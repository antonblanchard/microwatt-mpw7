module RAM32_1RW1R (CLK,
    EN0,
    EN1,
    VPWR,
    VGND,
    A0,
    A1,
    Di0,
    Do0,
    Do1,
    WE0);
 input CLK;
 input EN0;
 input EN1;
 input VPWR;
 input VGND;
 input [4:0] A0;
 input [4:0] A1;
 input [63:0] Di0;
 output [63:0] Do0;
 output [63:0] Do1;
 input [7:0] WE0;

 wire \A0BUF[0].X ;
 wire \A0BUF[1].X ;
 wire \A0BUF[2].X ;
 wire \A0BUF[3].X ;
 wire \A0BUF[4].X ;
 wire \A1BUF[0].X ;
 wire \A1BUF[1].X ;
 wire \A1BUF[2].X ;
 wire \A1BUF[3].X ;
 wire \A1BUF[4].X ;
 wire \BYTE[0].FLOATBUF0[0].A ;
 wire \BYTE[0].FLOATBUF0[0].TE_B ;
 wire \BYTE[0].FLOATBUF0[0].Z ;
 wire \BYTE[0].FLOATBUF0[1].Z ;
 wire \BYTE[0].FLOATBUF0[2].Z ;
 wire \BYTE[0].FLOATBUF0[3].Z ;
 wire \BYTE[0].FLOATBUF0[4].Z ;
 wire \BYTE[0].FLOATBUF0[5].Z ;
 wire \BYTE[0].FLOATBUF0[6].Z ;
 wire \BYTE[0].FLOATBUF0[7].Z ;
 wire \BYTE[0].FLOATBUF1[0].A ;
 wire \BYTE[0].FLOATBUF1[0].TE_B ;
 wire \BYTE[0].FLOATBUF1[0].Z ;
 wire \BYTE[0].FLOATBUF1[1].Z ;
 wire \BYTE[0].FLOATBUF1[2].Z ;
 wire \BYTE[0].FLOATBUF1[3].Z ;
 wire \BYTE[0].FLOATBUF1[4].Z ;
 wire \BYTE[0].FLOATBUF1[5].Z ;
 wire \BYTE[0].FLOATBUF1[6].Z ;
 wire \BYTE[0].FLOATBUF1[7].Z ;
 wire \BYTE[1].FLOATBUF0[10].A ;
 wire \BYTE[1].FLOATBUF0[10].TE_B ;
 wire \BYTE[1].FLOATBUF0[10].Z ;
 wire \BYTE[1].FLOATBUF0[11].Z ;
 wire \BYTE[1].FLOATBUF0[12].Z ;
 wire \BYTE[1].FLOATBUF0[13].Z ;
 wire \BYTE[1].FLOATBUF0[14].Z ;
 wire \BYTE[1].FLOATBUF0[15].Z ;
 wire \BYTE[1].FLOATBUF0[8].Z ;
 wire \BYTE[1].FLOATBUF0[9].Z ;
 wire \BYTE[1].FLOATBUF1[10].A ;
 wire \BYTE[1].FLOATBUF1[10].TE_B ;
 wire \BYTE[1].FLOATBUF1[10].Z ;
 wire \BYTE[1].FLOATBUF1[11].Z ;
 wire \BYTE[1].FLOATBUF1[12].Z ;
 wire \BYTE[1].FLOATBUF1[13].Z ;
 wire \BYTE[1].FLOATBUF1[14].Z ;
 wire \BYTE[1].FLOATBUF1[15].Z ;
 wire \BYTE[1].FLOATBUF1[8].Z ;
 wire \BYTE[1].FLOATBUF1[9].Z ;
 wire \BYTE[2].FLOATBUF0[16].A ;
 wire \BYTE[2].FLOATBUF0[16].TE_B ;
 wire \BYTE[2].FLOATBUF0[16].Z ;
 wire \BYTE[2].FLOATBUF0[17].Z ;
 wire \BYTE[2].FLOATBUF0[18].Z ;
 wire \BYTE[2].FLOATBUF0[19].Z ;
 wire \BYTE[2].FLOATBUF0[20].Z ;
 wire \BYTE[2].FLOATBUF0[21].Z ;
 wire \BYTE[2].FLOATBUF0[22].Z ;
 wire \BYTE[2].FLOATBUF0[23].Z ;
 wire \BYTE[2].FLOATBUF1[16].A ;
 wire \BYTE[2].FLOATBUF1[16].TE_B ;
 wire \BYTE[2].FLOATBUF1[16].Z ;
 wire \BYTE[2].FLOATBUF1[17].Z ;
 wire \BYTE[2].FLOATBUF1[18].Z ;
 wire \BYTE[2].FLOATBUF1[19].Z ;
 wire \BYTE[2].FLOATBUF1[20].Z ;
 wire \BYTE[2].FLOATBUF1[21].Z ;
 wire \BYTE[2].FLOATBUF1[22].Z ;
 wire \BYTE[2].FLOATBUF1[23].Z ;
 wire \BYTE[3].FLOATBUF0[24].A ;
 wire \BYTE[3].FLOATBUF0[24].TE_B ;
 wire \BYTE[3].FLOATBUF0[24].Z ;
 wire \BYTE[3].FLOATBUF0[25].Z ;
 wire \BYTE[3].FLOATBUF0[26].Z ;
 wire \BYTE[3].FLOATBUF0[27].Z ;
 wire \BYTE[3].FLOATBUF0[28].Z ;
 wire \BYTE[3].FLOATBUF0[29].Z ;
 wire \BYTE[3].FLOATBUF0[30].Z ;
 wire \BYTE[3].FLOATBUF0[31].Z ;
 wire \BYTE[3].FLOATBUF1[24].A ;
 wire \BYTE[3].FLOATBUF1[24].TE_B ;
 wire \BYTE[3].FLOATBUF1[24].Z ;
 wire \BYTE[3].FLOATBUF1[25].Z ;
 wire \BYTE[3].FLOATBUF1[26].Z ;
 wire \BYTE[3].FLOATBUF1[27].Z ;
 wire \BYTE[3].FLOATBUF1[28].Z ;
 wire \BYTE[3].FLOATBUF1[29].Z ;
 wire \BYTE[3].FLOATBUF1[30].Z ;
 wire \BYTE[3].FLOATBUF1[31].Z ;
 wire \BYTE[4].FLOATBUF0[32].A ;
 wire \BYTE[4].FLOATBUF0[32].TE_B ;
 wire \BYTE[4].FLOATBUF0[32].Z ;
 wire \BYTE[4].FLOATBUF0[33].Z ;
 wire \BYTE[4].FLOATBUF0[34].Z ;
 wire \BYTE[4].FLOATBUF0[35].Z ;
 wire \BYTE[4].FLOATBUF0[36].Z ;
 wire \BYTE[4].FLOATBUF0[37].Z ;
 wire \BYTE[4].FLOATBUF0[38].Z ;
 wire \BYTE[4].FLOATBUF0[39].Z ;
 wire \BYTE[4].FLOATBUF1[32].A ;
 wire \BYTE[4].FLOATBUF1[32].TE_B ;
 wire \BYTE[4].FLOATBUF1[32].Z ;
 wire \BYTE[4].FLOATBUF1[33].Z ;
 wire \BYTE[4].FLOATBUF1[34].Z ;
 wire \BYTE[4].FLOATBUF1[35].Z ;
 wire \BYTE[4].FLOATBUF1[36].Z ;
 wire \BYTE[4].FLOATBUF1[37].Z ;
 wire \BYTE[4].FLOATBUF1[38].Z ;
 wire \BYTE[4].FLOATBUF1[39].Z ;
 wire \BYTE[5].FLOATBUF0[40].A ;
 wire \BYTE[5].FLOATBUF0[40].TE_B ;
 wire \BYTE[5].FLOATBUF0[40].Z ;
 wire \BYTE[5].FLOATBUF0[41].Z ;
 wire \BYTE[5].FLOATBUF0[42].Z ;
 wire \BYTE[5].FLOATBUF0[43].Z ;
 wire \BYTE[5].FLOATBUF0[44].Z ;
 wire \BYTE[5].FLOATBUF0[45].Z ;
 wire \BYTE[5].FLOATBUF0[46].Z ;
 wire \BYTE[5].FLOATBUF0[47].Z ;
 wire \BYTE[5].FLOATBUF1[40].A ;
 wire \BYTE[5].FLOATBUF1[40].TE_B ;
 wire \BYTE[5].FLOATBUF1[40].Z ;
 wire \BYTE[5].FLOATBUF1[41].Z ;
 wire \BYTE[5].FLOATBUF1[42].Z ;
 wire \BYTE[5].FLOATBUF1[43].Z ;
 wire \BYTE[5].FLOATBUF1[44].Z ;
 wire \BYTE[5].FLOATBUF1[45].Z ;
 wire \BYTE[5].FLOATBUF1[46].Z ;
 wire \BYTE[5].FLOATBUF1[47].Z ;
 wire \BYTE[6].FLOATBUF0[48].A ;
 wire \BYTE[6].FLOATBUF0[48].TE_B ;
 wire \BYTE[6].FLOATBUF0[48].Z ;
 wire \BYTE[6].FLOATBUF0[49].Z ;
 wire \BYTE[6].FLOATBUF0[50].Z ;
 wire \BYTE[6].FLOATBUF0[51].Z ;
 wire \BYTE[6].FLOATBUF0[52].Z ;
 wire \BYTE[6].FLOATBUF0[53].Z ;
 wire \BYTE[6].FLOATBUF0[54].Z ;
 wire \BYTE[6].FLOATBUF0[55].Z ;
 wire \BYTE[6].FLOATBUF1[48].A ;
 wire \BYTE[6].FLOATBUF1[48].TE_B ;
 wire \BYTE[6].FLOATBUF1[48].Z ;
 wire \BYTE[6].FLOATBUF1[49].Z ;
 wire \BYTE[6].FLOATBUF1[50].Z ;
 wire \BYTE[6].FLOATBUF1[51].Z ;
 wire \BYTE[6].FLOATBUF1[52].Z ;
 wire \BYTE[6].FLOATBUF1[53].Z ;
 wire \BYTE[6].FLOATBUF1[54].Z ;
 wire \BYTE[6].FLOATBUF1[55].Z ;
 wire \BYTE[7].FLOATBUF0[56].A ;
 wire \BYTE[7].FLOATBUF0[56].TE_B ;
 wire \BYTE[7].FLOATBUF0[56].Z ;
 wire \BYTE[7].FLOATBUF0[57].Z ;
 wire \BYTE[7].FLOATBUF0[58].Z ;
 wire \BYTE[7].FLOATBUF0[59].Z ;
 wire \BYTE[7].FLOATBUF0[60].Z ;
 wire \BYTE[7].FLOATBUF0[61].Z ;
 wire \BYTE[7].FLOATBUF0[62].Z ;
 wire \BYTE[7].FLOATBUF0[63].Z ;
 wire \BYTE[7].FLOATBUF1[56].A ;
 wire \BYTE[7].FLOATBUF1[56].TE_B ;
 wire \BYTE[7].FLOATBUF1[56].Z ;
 wire \BYTE[7].FLOATBUF1[57].Z ;
 wire \BYTE[7].FLOATBUF1[58].Z ;
 wire \BYTE[7].FLOATBUF1[59].Z ;
 wire \BYTE[7].FLOATBUF1[60].Z ;
 wire \BYTE[7].FLOATBUF1[61].Z ;
 wire \BYTE[7].FLOATBUF1[62].Z ;
 wire \BYTE[7].FLOATBUF1[63].Z ;
 wire \CLKBUF.X ;
 wire \DEC0.EN ;
 wire \DEC1.EN ;
 wire \DIBUF[0].X ;
 wire \DIBUF[10].X ;
 wire \DIBUF[11].X ;
 wire \DIBUF[12].X ;
 wire \DIBUF[13].X ;
 wire \DIBUF[14].X ;
 wire \DIBUF[15].X ;
 wire \DIBUF[16].X ;
 wire \DIBUF[17].X ;
 wire \DIBUF[18].X ;
 wire \DIBUF[19].X ;
 wire \DIBUF[1].X ;
 wire \DIBUF[20].X ;
 wire \DIBUF[21].X ;
 wire \DIBUF[22].X ;
 wire \DIBUF[23].X ;
 wire \DIBUF[24].X ;
 wire \DIBUF[25].X ;
 wire \DIBUF[26].X ;
 wire \DIBUF[27].X ;
 wire \DIBUF[28].X ;
 wire \DIBUF[29].X ;
 wire \DIBUF[2].X ;
 wire \DIBUF[30].X ;
 wire \DIBUF[31].X ;
 wire \DIBUF[32].X ;
 wire \DIBUF[33].X ;
 wire \DIBUF[34].X ;
 wire \DIBUF[35].X ;
 wire \DIBUF[36].X ;
 wire \DIBUF[37].X ;
 wire \DIBUF[38].X ;
 wire \DIBUF[39].X ;
 wire \DIBUF[3].X ;
 wire \DIBUF[40].X ;
 wire \DIBUF[41].X ;
 wire \DIBUF[42].X ;
 wire \DIBUF[43].X ;
 wire \DIBUF[44].X ;
 wire \DIBUF[45].X ;
 wire \DIBUF[46].X ;
 wire \DIBUF[47].X ;
 wire \DIBUF[48].X ;
 wire \DIBUF[49].X ;
 wire \DIBUF[4].X ;
 wire \DIBUF[50].X ;
 wire \DIBUF[51].X ;
 wire \DIBUF[52].X ;
 wire \DIBUF[53].X ;
 wire \DIBUF[54].X ;
 wire \DIBUF[55].X ;
 wire \DIBUF[56].X ;
 wire \DIBUF[57].X ;
 wire \DIBUF[58].X ;
 wire \DIBUF[59].X ;
 wire \DIBUF[5].X ;
 wire \DIBUF[60].X ;
 wire \DIBUF[61].X ;
 wire \DIBUF[62].X ;
 wire \DIBUF[63].X ;
 wire \DIBUF[6].X ;
 wire \DIBUF[7].X ;
 wire \DIBUF[8].X ;
 wire \DIBUF[9].X ;
 wire \Do0_REG.CLKBUF[0] ;
 wire \Do0_REG.CLKBUF[1] ;
 wire \Do0_REG.CLKBUF[2] ;
 wire \Do0_REG.CLKBUF[3] ;
 wire \Do0_REG.CLKBUF[4] ;
 wire \Do0_REG.CLKBUF[5] ;
 wire \Do0_REG.CLKBUF[6] ;
 wire \Do0_REG.CLKBUF[7] ;
 wire \Do0_REG.CLK_buf ;
 wire \Do1_REG.CLKBUF[0] ;
 wire \Do1_REG.CLKBUF[1] ;
 wire \Do1_REG.CLKBUF[2] ;
 wire \Do1_REG.CLKBUF[3] ;
 wire \Do1_REG.CLKBUF[4] ;
 wire \Do1_REG.CLKBUF[5] ;
 wire \Do1_REG.CLKBUF[6] ;
 wire \Do1_REG.CLKBUF[7] ;
 wire \Do1_REG.CLK_buf ;
 wire \SLICE[0].RAM8.CLKBUF.X ;
 wire \SLICE[0].RAM8.DEC0.A_buf[0] ;
 wire \SLICE[0].RAM8.DEC0.A_buf[1] ;
 wire \SLICE[0].RAM8.DEC0.A_buf[2] ;
 wire \SLICE[0].RAM8.DEC0.EN ;
 wire \SLICE[0].RAM8.DEC0.EN_buf ;
 wire \SLICE[0].RAM8.DEC1.A_buf[0] ;
 wire \SLICE[0].RAM8.DEC1.A_buf[1] ;
 wire \SLICE[0].RAM8.DEC1.A_buf[2] ;
 wire \SLICE[0].RAM8.DEC1.EN ;
 wire \SLICE[0].RAM8.DEC1.EN_buf ;
 wire \SLICE[0].RAM8.WEBUF[0].A ;
 wire \SLICE[0].RAM8.WEBUF[0].X ;
 wire \SLICE[0].RAM8.WEBUF[1].A ;
 wire \SLICE[0].RAM8.WEBUF[1].X ;
 wire \SLICE[0].RAM8.WEBUF[2].A ;
 wire \SLICE[0].RAM8.WEBUF[2].X ;
 wire \SLICE[0].RAM8.WEBUF[3].A ;
 wire \SLICE[0].RAM8.WEBUF[3].X ;
 wire \SLICE[0].RAM8.WEBUF[4].A ;
 wire \SLICE[0].RAM8.WEBUF[4].X ;
 wire \SLICE[0].RAM8.WEBUF[5].A ;
 wire \SLICE[0].RAM8.WEBUF[5].X ;
 wire \SLICE[0].RAM8.WEBUF[6].A ;
 wire \SLICE[0].RAM8.WEBUF[6].X ;
 wire \SLICE[0].RAM8.WEBUF[7].A ;
 wire \SLICE[0].RAM8.WEBUF[7].X ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1 ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[0].W.SEL0 ;
 wire \SLICE[0].RAM8.WORD[0].W.SEL1 ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1 ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[1].W.SEL0 ;
 wire \SLICE[0].RAM8.WORD[1].W.SEL1 ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1 ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[2].W.SEL0 ;
 wire \SLICE[0].RAM8.WORD[2].W.SEL1 ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1 ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[3].W.SEL0 ;
 wire \SLICE[0].RAM8.WORD[3].W.SEL1 ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1 ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[4].W.SEL0 ;
 wire \SLICE[0].RAM8.WORD[4].W.SEL1 ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1 ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[5].W.SEL0 ;
 wire \SLICE[0].RAM8.WORD[5].W.SEL1 ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1 ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[6].W.SEL0 ;
 wire \SLICE[0].RAM8.WORD[6].W.SEL1 ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1 ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[7].W.SEL0 ;
 wire \SLICE[0].RAM8.WORD[7].W.SEL1 ;
 wire \SLICE[1].RAM8.CLKBUF.X ;
 wire \SLICE[1].RAM8.DEC0.A_buf[0] ;
 wire \SLICE[1].RAM8.DEC0.A_buf[1] ;
 wire \SLICE[1].RAM8.DEC0.A_buf[2] ;
 wire \SLICE[1].RAM8.DEC0.EN ;
 wire \SLICE[1].RAM8.DEC0.EN_buf ;
 wire \SLICE[1].RAM8.DEC1.A_buf[0] ;
 wire \SLICE[1].RAM8.DEC1.A_buf[1] ;
 wire \SLICE[1].RAM8.DEC1.A_buf[2] ;
 wire \SLICE[1].RAM8.DEC1.EN ;
 wire \SLICE[1].RAM8.DEC1.EN_buf ;
 wire \SLICE[1].RAM8.WEBUF[0].X ;
 wire \SLICE[1].RAM8.WEBUF[1].X ;
 wire \SLICE[1].RAM8.WEBUF[2].X ;
 wire \SLICE[1].RAM8.WEBUF[3].X ;
 wire \SLICE[1].RAM8.WEBUF[4].X ;
 wire \SLICE[1].RAM8.WEBUF[5].X ;
 wire \SLICE[1].RAM8.WEBUF[6].X ;
 wire \SLICE[1].RAM8.WEBUF[7].X ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1 ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[0].W.SEL0 ;
 wire \SLICE[1].RAM8.WORD[0].W.SEL1 ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1 ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[1].W.SEL0 ;
 wire \SLICE[1].RAM8.WORD[1].W.SEL1 ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1 ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[2].W.SEL0 ;
 wire \SLICE[1].RAM8.WORD[2].W.SEL1 ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1 ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[3].W.SEL0 ;
 wire \SLICE[1].RAM8.WORD[3].W.SEL1 ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1 ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[4].W.SEL0 ;
 wire \SLICE[1].RAM8.WORD[4].W.SEL1 ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1 ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[5].W.SEL0 ;
 wire \SLICE[1].RAM8.WORD[5].W.SEL1 ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1 ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[6].W.SEL0 ;
 wire \SLICE[1].RAM8.WORD[6].W.SEL1 ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1 ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[7].W.SEL0 ;
 wire \SLICE[1].RAM8.WORD[7].W.SEL1 ;
 wire \SLICE[2].RAM8.CLKBUF.X ;
 wire \SLICE[2].RAM8.DEC0.A_buf[0] ;
 wire \SLICE[2].RAM8.DEC0.A_buf[1] ;
 wire \SLICE[2].RAM8.DEC0.A_buf[2] ;
 wire \SLICE[2].RAM8.DEC0.EN ;
 wire \SLICE[2].RAM8.DEC0.EN_buf ;
 wire \SLICE[2].RAM8.DEC1.A_buf[0] ;
 wire \SLICE[2].RAM8.DEC1.A_buf[1] ;
 wire \SLICE[2].RAM8.DEC1.A_buf[2] ;
 wire \SLICE[2].RAM8.DEC1.EN ;
 wire \SLICE[2].RAM8.DEC1.EN_buf ;
 wire \SLICE[2].RAM8.WEBUF[0].X ;
 wire \SLICE[2].RAM8.WEBUF[1].X ;
 wire \SLICE[2].RAM8.WEBUF[2].X ;
 wire \SLICE[2].RAM8.WEBUF[3].X ;
 wire \SLICE[2].RAM8.WEBUF[4].X ;
 wire \SLICE[2].RAM8.WEBUF[5].X ;
 wire \SLICE[2].RAM8.WEBUF[6].X ;
 wire \SLICE[2].RAM8.WEBUF[7].X ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1 ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[0].W.SEL0 ;
 wire \SLICE[2].RAM8.WORD[0].W.SEL1 ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1 ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[1].W.SEL0 ;
 wire \SLICE[2].RAM8.WORD[1].W.SEL1 ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1 ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[2].W.SEL0 ;
 wire \SLICE[2].RAM8.WORD[2].W.SEL1 ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1 ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[3].W.SEL0 ;
 wire \SLICE[2].RAM8.WORD[3].W.SEL1 ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1 ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[4].W.SEL0 ;
 wire \SLICE[2].RAM8.WORD[4].W.SEL1 ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1 ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[5].W.SEL0 ;
 wire \SLICE[2].RAM8.WORD[5].W.SEL1 ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1 ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[6].W.SEL0 ;
 wire \SLICE[2].RAM8.WORD[6].W.SEL1 ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1 ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[7].W.SEL0 ;
 wire \SLICE[2].RAM8.WORD[7].W.SEL1 ;
 wire \SLICE[3].RAM8.CLKBUF.X ;
 wire \SLICE[3].RAM8.DEC0.A_buf[0] ;
 wire \SLICE[3].RAM8.DEC0.A_buf[1] ;
 wire \SLICE[3].RAM8.DEC0.A_buf[2] ;
 wire \SLICE[3].RAM8.DEC0.EN ;
 wire \SLICE[3].RAM8.DEC0.EN_buf ;
 wire \SLICE[3].RAM8.DEC1.A_buf[0] ;
 wire \SLICE[3].RAM8.DEC1.A_buf[1] ;
 wire \SLICE[3].RAM8.DEC1.A_buf[2] ;
 wire \SLICE[3].RAM8.DEC1.EN ;
 wire \SLICE[3].RAM8.DEC1.EN_buf ;
 wire \SLICE[3].RAM8.WEBUF[0].X ;
 wire \SLICE[3].RAM8.WEBUF[1].X ;
 wire \SLICE[3].RAM8.WEBUF[2].X ;
 wire \SLICE[3].RAM8.WEBUF[3].X ;
 wire \SLICE[3].RAM8.WEBUF[4].X ;
 wire \SLICE[3].RAM8.WEBUF[5].X ;
 wire \SLICE[3].RAM8.WEBUF[6].X ;
 wire \SLICE[3].RAM8.WEBUF[7].X ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1 ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[0].W.SEL0 ;
 wire \SLICE[3].RAM8.WORD[0].W.SEL1 ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1 ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[1].W.SEL0 ;
 wire \SLICE[3].RAM8.WORD[1].W.SEL1 ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1 ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[2].W.SEL0 ;
 wire \SLICE[3].RAM8.WORD[2].W.SEL1 ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1 ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[3].W.SEL0 ;
 wire \SLICE[3].RAM8.WORD[3].W.SEL1 ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1 ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[4].W.SEL0 ;
 wire \SLICE[3].RAM8.WORD[4].W.SEL1 ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1 ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[5].W.SEL0 ;
 wire \SLICE[3].RAM8.WORD[5].W.SEL1 ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1 ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[6].W.SEL0 ;
 wire \SLICE[3].RAM8.WORD[6].W.SEL1 ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1 ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[7].W.SEL0 ;
 wire \SLICE[3].RAM8.WORD[7].W.SEL1 ;

 sky130_fd_sc_hd__clkbuf_2 \A0BUF[0].__cell__  (.A(A0[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \A0BUF[1].__cell__  (.A(A0[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \A0BUF[2].__cell__  (.A(A0[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \A0BUF[3].__cell__  (.A(A0[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\A0BUF[3].X ));
 sky130_fd_sc_hd__clkbuf_2 \A0BUF[4].__cell__  (.A(A0[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\A0BUF[4].X ));
 sky130_fd_sc_hd__clkbuf_2 \A1BUF[0].__cell__  (.A(A1[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\A1BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \A1BUF[1].__cell__  (.A(A1[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\A1BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \A1BUF[2].__cell__  (.A(A1[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\A1BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \A1BUF[3].__cell__  (.A(A1[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\A1BUF[3].X ));
 sky130_fd_sc_hd__clkbuf_2 \A1BUF[4].__cell__  (.A(A1[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\A1BUF[4].X ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[0].FLOATBUF0[0].__cell__  (.A(\BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BYTE[0].FLOATBUF0[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[0].FLOATBUF0[1].__cell__  (.A(\BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BYTE[0].FLOATBUF0[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[0].FLOATBUF0[2].__cell__  (.A(\BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BYTE[0].FLOATBUF0[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[0].FLOATBUF0[3].__cell__  (.A(\BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BYTE[0].FLOATBUF0[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[0].FLOATBUF0[4].__cell__  (.A(\BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BYTE[0].FLOATBUF0[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[0].FLOATBUF0[5].__cell__  (.A(\BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BYTE[0].FLOATBUF0[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[0].FLOATBUF0[6].__cell__  (.A(\BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BYTE[0].FLOATBUF0[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[0].FLOATBUF0[7].__cell__  (.A(\BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BYTE[0].FLOATBUF0[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[0].FLOATBUF1[0].__cell__  (.A(\BYTE[0].FLOATBUF1[0].A ),
    .TE_B(\BYTE[0].FLOATBUF1[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[0].FLOATBUF1[1].__cell__  (.A(\BYTE[0].FLOATBUF1[0].A ),
    .TE_B(\BYTE[0].FLOATBUF1[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[0].FLOATBUF1[2].__cell__  (.A(\BYTE[0].FLOATBUF1[0].A ),
    .TE_B(\BYTE[0].FLOATBUF1[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[0].FLOATBUF1[3].__cell__  (.A(\BYTE[0].FLOATBUF1[0].A ),
    .TE_B(\BYTE[0].FLOATBUF1[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[0].FLOATBUF1[4].__cell__  (.A(\BYTE[0].FLOATBUF1[0].A ),
    .TE_B(\BYTE[0].FLOATBUF1[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[0].FLOATBUF1[5].__cell__  (.A(\BYTE[0].FLOATBUF1[0].A ),
    .TE_B(\BYTE[0].FLOATBUF1[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[0].FLOATBUF1[6].__cell__  (.A(\BYTE[0].FLOATBUF1[0].A ),
    .TE_B(\BYTE[0].FLOATBUF1[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[0].FLOATBUF1[7].__cell__  (.A(\BYTE[0].FLOATBUF1[0].A ),
    .TE_B(\BYTE[0].FLOATBUF1[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[1].FLOATBUF0[10].__cell__  (.A(\BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BYTE[1].FLOATBUF0[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[1].FLOATBUF0[11].__cell__  (.A(\BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BYTE[1].FLOATBUF0[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[1].FLOATBUF0[12].__cell__  (.A(\BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BYTE[1].FLOATBUF0[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[1].FLOATBUF0[13].__cell__  (.A(\BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BYTE[1].FLOATBUF0[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[1].FLOATBUF0[14].__cell__  (.A(\BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BYTE[1].FLOATBUF0[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[1].FLOATBUF0[15].__cell__  (.A(\BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BYTE[1].FLOATBUF0[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[1].FLOATBUF0[8].__cell__  (.A(\BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BYTE[1].FLOATBUF0[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[1].FLOATBUF0[9].__cell__  (.A(\BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BYTE[1].FLOATBUF0[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[1].FLOATBUF1[10].__cell__  (.A(\BYTE[1].FLOATBUF1[10].A ),
    .TE_B(\BYTE[1].FLOATBUF1[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[1].FLOATBUF1[11].__cell__  (.A(\BYTE[1].FLOATBUF1[10].A ),
    .TE_B(\BYTE[1].FLOATBUF1[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[1].FLOATBUF1[12].__cell__  (.A(\BYTE[1].FLOATBUF1[10].A ),
    .TE_B(\BYTE[1].FLOATBUF1[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[1].FLOATBUF1[13].__cell__  (.A(\BYTE[1].FLOATBUF1[10].A ),
    .TE_B(\BYTE[1].FLOATBUF1[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[1].FLOATBUF1[14].__cell__  (.A(\BYTE[1].FLOATBUF1[10].A ),
    .TE_B(\BYTE[1].FLOATBUF1[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[1].FLOATBUF1[15].__cell__  (.A(\BYTE[1].FLOATBUF1[10].A ),
    .TE_B(\BYTE[1].FLOATBUF1[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[1].FLOATBUF1[8].__cell__  (.A(\BYTE[1].FLOATBUF1[10].A ),
    .TE_B(\BYTE[1].FLOATBUF1[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[1].FLOATBUF1[9].__cell__  (.A(\BYTE[1].FLOATBUF1[10].A ),
    .TE_B(\BYTE[1].FLOATBUF1[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[2].FLOATBUF0[16].__cell__  (.A(\BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BYTE[2].FLOATBUF0[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[2].FLOATBUF0[17].__cell__  (.A(\BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BYTE[2].FLOATBUF0[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[2].FLOATBUF0[18].__cell__  (.A(\BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BYTE[2].FLOATBUF0[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[2].FLOATBUF0[19].__cell__  (.A(\BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BYTE[2].FLOATBUF0[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[2].FLOATBUF0[20].__cell__  (.A(\BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BYTE[2].FLOATBUF0[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[2].FLOATBUF0[21].__cell__  (.A(\BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BYTE[2].FLOATBUF0[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[2].FLOATBUF0[22].__cell__  (.A(\BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BYTE[2].FLOATBUF0[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[2].FLOATBUF0[23].__cell__  (.A(\BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BYTE[2].FLOATBUF0[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[2].FLOATBUF1[16].__cell__  (.A(\BYTE[2].FLOATBUF1[16].A ),
    .TE_B(\BYTE[2].FLOATBUF1[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[2].FLOATBUF1[17].__cell__  (.A(\BYTE[2].FLOATBUF1[16].A ),
    .TE_B(\BYTE[2].FLOATBUF1[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[2].FLOATBUF1[18].__cell__  (.A(\BYTE[2].FLOATBUF1[16].A ),
    .TE_B(\BYTE[2].FLOATBUF1[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[2].FLOATBUF1[19].__cell__  (.A(\BYTE[2].FLOATBUF1[16].A ),
    .TE_B(\BYTE[2].FLOATBUF1[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[2].FLOATBUF1[20].__cell__  (.A(\BYTE[2].FLOATBUF1[16].A ),
    .TE_B(\BYTE[2].FLOATBUF1[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[2].FLOATBUF1[21].__cell__  (.A(\BYTE[2].FLOATBUF1[16].A ),
    .TE_B(\BYTE[2].FLOATBUF1[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[2].FLOATBUF1[22].__cell__  (.A(\BYTE[2].FLOATBUF1[16].A ),
    .TE_B(\BYTE[2].FLOATBUF1[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[2].FLOATBUF1[23].__cell__  (.A(\BYTE[2].FLOATBUF1[16].A ),
    .TE_B(\BYTE[2].FLOATBUF1[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[3].FLOATBUF0[24].__cell__  (.A(\BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BYTE[3].FLOATBUF0[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[3].FLOATBUF0[25].__cell__  (.A(\BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BYTE[3].FLOATBUF0[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[3].FLOATBUF0[26].__cell__  (.A(\BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BYTE[3].FLOATBUF0[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[3].FLOATBUF0[27].__cell__  (.A(\BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BYTE[3].FLOATBUF0[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[3].FLOATBUF0[28].__cell__  (.A(\BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BYTE[3].FLOATBUF0[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[3].FLOATBUF0[29].__cell__  (.A(\BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BYTE[3].FLOATBUF0[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[3].FLOATBUF0[30].__cell__  (.A(\BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BYTE[3].FLOATBUF0[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[3].FLOATBUF0[31].__cell__  (.A(\BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BYTE[3].FLOATBUF0[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[3].FLOATBUF1[24].__cell__  (.A(\BYTE[3].FLOATBUF1[24].A ),
    .TE_B(\BYTE[3].FLOATBUF1[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[3].FLOATBUF1[25].__cell__  (.A(\BYTE[3].FLOATBUF1[24].A ),
    .TE_B(\BYTE[3].FLOATBUF1[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[3].FLOATBUF1[26].__cell__  (.A(\BYTE[3].FLOATBUF1[24].A ),
    .TE_B(\BYTE[3].FLOATBUF1[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[3].FLOATBUF1[27].__cell__  (.A(\BYTE[3].FLOATBUF1[24].A ),
    .TE_B(\BYTE[3].FLOATBUF1[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[3].FLOATBUF1[28].__cell__  (.A(\BYTE[3].FLOATBUF1[24].A ),
    .TE_B(\BYTE[3].FLOATBUF1[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[3].FLOATBUF1[29].__cell__  (.A(\BYTE[3].FLOATBUF1[24].A ),
    .TE_B(\BYTE[3].FLOATBUF1[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[3].FLOATBUF1[30].__cell__  (.A(\BYTE[3].FLOATBUF1[24].A ),
    .TE_B(\BYTE[3].FLOATBUF1[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[3].FLOATBUF1[31].__cell__  (.A(\BYTE[3].FLOATBUF1[24].A ),
    .TE_B(\BYTE[3].FLOATBUF1[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[4].FLOATBUF0[32].__cell__  (.A(\BYTE[4].FLOATBUF0[32].A ),
    .TE_B(\BYTE[4].FLOATBUF0[32].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[4].FLOATBUF0[33].__cell__  (.A(\BYTE[4].FLOATBUF0[32].A ),
    .TE_B(\BYTE[4].FLOATBUF0[32].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[4].FLOATBUF0[34].__cell__  (.A(\BYTE[4].FLOATBUF0[32].A ),
    .TE_B(\BYTE[4].FLOATBUF0[32].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[4].FLOATBUF0[35].__cell__  (.A(\BYTE[4].FLOATBUF0[32].A ),
    .TE_B(\BYTE[4].FLOATBUF0[32].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[4].FLOATBUF0[36].__cell__  (.A(\BYTE[4].FLOATBUF0[32].A ),
    .TE_B(\BYTE[4].FLOATBUF0[32].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[4].FLOATBUF0[37].__cell__  (.A(\BYTE[4].FLOATBUF0[32].A ),
    .TE_B(\BYTE[4].FLOATBUF0[32].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[4].FLOATBUF0[38].__cell__  (.A(\BYTE[4].FLOATBUF0[32].A ),
    .TE_B(\BYTE[4].FLOATBUF0[32].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[4].FLOATBUF0[39].__cell__  (.A(\BYTE[4].FLOATBUF0[32].A ),
    .TE_B(\BYTE[4].FLOATBUF0[32].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[4].FLOATBUF1[32].__cell__  (.A(\BYTE[4].FLOATBUF1[32].A ),
    .TE_B(\BYTE[4].FLOATBUF1[32].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[4].FLOATBUF1[33].__cell__  (.A(\BYTE[4].FLOATBUF1[32].A ),
    .TE_B(\BYTE[4].FLOATBUF1[32].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[4].FLOATBUF1[34].__cell__  (.A(\BYTE[4].FLOATBUF1[32].A ),
    .TE_B(\BYTE[4].FLOATBUF1[32].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[4].FLOATBUF1[35].__cell__  (.A(\BYTE[4].FLOATBUF1[32].A ),
    .TE_B(\BYTE[4].FLOATBUF1[32].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[4].FLOATBUF1[36].__cell__  (.A(\BYTE[4].FLOATBUF1[32].A ),
    .TE_B(\BYTE[4].FLOATBUF1[32].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[4].FLOATBUF1[37].__cell__  (.A(\BYTE[4].FLOATBUF1[32].A ),
    .TE_B(\BYTE[4].FLOATBUF1[32].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[4].FLOATBUF1[38].__cell__  (.A(\BYTE[4].FLOATBUF1[32].A ),
    .TE_B(\BYTE[4].FLOATBUF1[32].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[4].FLOATBUF1[39].__cell__  (.A(\BYTE[4].FLOATBUF1[32].A ),
    .TE_B(\BYTE[4].FLOATBUF1[32].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[5].FLOATBUF0[40].__cell__  (.A(\BYTE[5].FLOATBUF0[40].A ),
    .TE_B(\BYTE[5].FLOATBUF0[40].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[5].FLOATBUF0[41].__cell__  (.A(\BYTE[5].FLOATBUF0[40].A ),
    .TE_B(\BYTE[5].FLOATBUF0[40].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[5].FLOATBUF0[42].__cell__  (.A(\BYTE[5].FLOATBUF0[40].A ),
    .TE_B(\BYTE[5].FLOATBUF0[40].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[5].FLOATBUF0[43].__cell__  (.A(\BYTE[5].FLOATBUF0[40].A ),
    .TE_B(\BYTE[5].FLOATBUF0[40].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[5].FLOATBUF0[44].__cell__  (.A(\BYTE[5].FLOATBUF0[40].A ),
    .TE_B(\BYTE[5].FLOATBUF0[40].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[5].FLOATBUF0[45].__cell__  (.A(\BYTE[5].FLOATBUF0[40].A ),
    .TE_B(\BYTE[5].FLOATBUF0[40].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[5].FLOATBUF0[46].__cell__  (.A(\BYTE[5].FLOATBUF0[40].A ),
    .TE_B(\BYTE[5].FLOATBUF0[40].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[5].FLOATBUF0[47].__cell__  (.A(\BYTE[5].FLOATBUF0[40].A ),
    .TE_B(\BYTE[5].FLOATBUF0[40].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[5].FLOATBUF1[40].__cell__  (.A(\BYTE[5].FLOATBUF1[40].A ),
    .TE_B(\BYTE[5].FLOATBUF1[40].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[5].FLOATBUF1[41].__cell__  (.A(\BYTE[5].FLOATBUF1[40].A ),
    .TE_B(\BYTE[5].FLOATBUF1[40].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[5].FLOATBUF1[42].__cell__  (.A(\BYTE[5].FLOATBUF1[40].A ),
    .TE_B(\BYTE[5].FLOATBUF1[40].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[5].FLOATBUF1[43].__cell__  (.A(\BYTE[5].FLOATBUF1[40].A ),
    .TE_B(\BYTE[5].FLOATBUF1[40].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[5].FLOATBUF1[44].__cell__  (.A(\BYTE[5].FLOATBUF1[40].A ),
    .TE_B(\BYTE[5].FLOATBUF1[40].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[5].FLOATBUF1[45].__cell__  (.A(\BYTE[5].FLOATBUF1[40].A ),
    .TE_B(\BYTE[5].FLOATBUF1[40].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[5].FLOATBUF1[46].__cell__  (.A(\BYTE[5].FLOATBUF1[40].A ),
    .TE_B(\BYTE[5].FLOATBUF1[40].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[5].FLOATBUF1[47].__cell__  (.A(\BYTE[5].FLOATBUF1[40].A ),
    .TE_B(\BYTE[5].FLOATBUF1[40].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[6].FLOATBUF0[48].__cell__  (.A(\BYTE[6].FLOATBUF0[48].A ),
    .TE_B(\BYTE[6].FLOATBUF0[48].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[6].FLOATBUF0[49].__cell__  (.A(\BYTE[6].FLOATBUF0[48].A ),
    .TE_B(\BYTE[6].FLOATBUF0[48].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[6].FLOATBUF0[50].__cell__  (.A(\BYTE[6].FLOATBUF0[48].A ),
    .TE_B(\BYTE[6].FLOATBUF0[48].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[6].FLOATBUF0[51].__cell__  (.A(\BYTE[6].FLOATBUF0[48].A ),
    .TE_B(\BYTE[6].FLOATBUF0[48].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[6].FLOATBUF0[52].__cell__  (.A(\BYTE[6].FLOATBUF0[48].A ),
    .TE_B(\BYTE[6].FLOATBUF0[48].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[6].FLOATBUF0[53].__cell__  (.A(\BYTE[6].FLOATBUF0[48].A ),
    .TE_B(\BYTE[6].FLOATBUF0[48].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[6].FLOATBUF0[54].__cell__  (.A(\BYTE[6].FLOATBUF0[48].A ),
    .TE_B(\BYTE[6].FLOATBUF0[48].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[6].FLOATBUF0[55].__cell__  (.A(\BYTE[6].FLOATBUF0[48].A ),
    .TE_B(\BYTE[6].FLOATBUF0[48].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[6].FLOATBUF1[48].__cell__  (.A(\BYTE[6].FLOATBUF1[48].A ),
    .TE_B(\BYTE[6].FLOATBUF1[48].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[6].FLOATBUF1[49].__cell__  (.A(\BYTE[6].FLOATBUF1[48].A ),
    .TE_B(\BYTE[6].FLOATBUF1[48].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[6].FLOATBUF1[50].__cell__  (.A(\BYTE[6].FLOATBUF1[48].A ),
    .TE_B(\BYTE[6].FLOATBUF1[48].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[6].FLOATBUF1[51].__cell__  (.A(\BYTE[6].FLOATBUF1[48].A ),
    .TE_B(\BYTE[6].FLOATBUF1[48].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[6].FLOATBUF1[52].__cell__  (.A(\BYTE[6].FLOATBUF1[48].A ),
    .TE_B(\BYTE[6].FLOATBUF1[48].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[6].FLOATBUF1[53].__cell__  (.A(\BYTE[6].FLOATBUF1[48].A ),
    .TE_B(\BYTE[6].FLOATBUF1[48].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[6].FLOATBUF1[54].__cell__  (.A(\BYTE[6].FLOATBUF1[48].A ),
    .TE_B(\BYTE[6].FLOATBUF1[48].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[6].FLOATBUF1[55].__cell__  (.A(\BYTE[6].FLOATBUF1[48].A ),
    .TE_B(\BYTE[6].FLOATBUF1[48].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[7].FLOATBUF0[56].__cell__  (.A(\BYTE[7].FLOATBUF0[56].A ),
    .TE_B(\BYTE[7].FLOATBUF0[56].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[7].FLOATBUF0[57].__cell__  (.A(\BYTE[7].FLOATBUF0[56].A ),
    .TE_B(\BYTE[7].FLOATBUF0[56].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[7].FLOATBUF0[58].__cell__  (.A(\BYTE[7].FLOATBUF0[56].A ),
    .TE_B(\BYTE[7].FLOATBUF0[56].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[7].FLOATBUF0[59].__cell__  (.A(\BYTE[7].FLOATBUF0[56].A ),
    .TE_B(\BYTE[7].FLOATBUF0[56].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[7].FLOATBUF0[60].__cell__  (.A(\BYTE[7].FLOATBUF0[56].A ),
    .TE_B(\BYTE[7].FLOATBUF0[56].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[7].FLOATBUF0[61].__cell__  (.A(\BYTE[7].FLOATBUF0[56].A ),
    .TE_B(\BYTE[7].FLOATBUF0[56].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[7].FLOATBUF0[62].__cell__  (.A(\BYTE[7].FLOATBUF0[56].A ),
    .TE_B(\BYTE[7].FLOATBUF0[56].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[7].FLOATBUF0[63].__cell__  (.A(\BYTE[7].FLOATBUF0[56].A ),
    .TE_B(\BYTE[7].FLOATBUF0[56].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[7].FLOATBUF1[56].__cell__  (.A(\BYTE[7].FLOATBUF1[56].A ),
    .TE_B(\BYTE[7].FLOATBUF1[56].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[7].FLOATBUF1[57].__cell__  (.A(\BYTE[7].FLOATBUF1[56].A ),
    .TE_B(\BYTE[7].FLOATBUF1[56].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[7].FLOATBUF1[58].__cell__  (.A(\BYTE[7].FLOATBUF1[56].A ),
    .TE_B(\BYTE[7].FLOATBUF1[56].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[7].FLOATBUF1[59].__cell__  (.A(\BYTE[7].FLOATBUF1[56].A ),
    .TE_B(\BYTE[7].FLOATBUF1[56].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[7].FLOATBUF1[60].__cell__  (.A(\BYTE[7].FLOATBUF1[56].A ),
    .TE_B(\BYTE[7].FLOATBUF1[56].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[7].FLOATBUF1[61].__cell__  (.A(\BYTE[7].FLOATBUF1[56].A ),
    .TE_B(\BYTE[7].FLOATBUF1[56].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[7].FLOATBUF1[62].__cell__  (.A(\BYTE[7].FLOATBUF1[56].A ),
    .TE_B(\BYTE[7].FLOATBUF1[56].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \BYTE[7].FLOATBUF1[63].__cell__  (.A(\BYTE[7].FLOATBUF1[56].A ),
    .TE_B(\BYTE[7].FLOATBUF1[56].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__clkbuf_4 \CLKBUF.__cell__  (.A(CLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\CLKBUF.X ));
 sky130_fd_sc_hd__nor3b_2 \DEC0.AND0  (.A(\A0BUF[3].X ),
    .B(\A0BUF[4].X ),
    .C_N(\DEC0.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and3b_2 \DEC0.AND1  (.A_N(\A0BUF[4].X ),
    .B(\A0BUF[3].X ),
    .C(\DEC0.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and3b_2 \DEC0.AND2  (.A_N(\A0BUF[3].X ),
    .B(\A0BUF[4].X ),
    .C(\DEC0.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and3_2 \DEC0.AND3  (.A(\A0BUF[4].X ),
    .B(\A0BUF[3].X ),
    .C(\DEC0.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__nor3b_2 \DEC1.AND0  (.A(\A1BUF[3].X ),
    .B(\A1BUF[4].X ),
    .C_N(\DEC1.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.DEC1.EN ));
 sky130_fd_sc_hd__and3b_2 \DEC1.AND1  (.A_N(\A1BUF[4].X ),
    .B(\A1BUF[3].X ),
    .C(\DEC1.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.DEC1.EN ));
 sky130_fd_sc_hd__and3b_2 \DEC1.AND2  (.A_N(\A1BUF[3].X ),
    .B(\A1BUF[4].X ),
    .C(\DEC1.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.DEC1.EN ));
 sky130_fd_sc_hd__and3_2 \DEC1.AND3  (.A(\A1BUF[4].X ),
    .B(\A1BUF[3].X ),
    .C(\DEC1.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.DEC1.EN ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[0].__cell__  (.A(Di0[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[10].__cell__  (.A(Di0[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[10].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[11].__cell__  (.A(Di0[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[11].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[12].__cell__  (.A(Di0[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[12].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[13].__cell__  (.A(Di0[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[13].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[14].__cell__  (.A(Di0[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[14].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[15].__cell__  (.A(Di0[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[15].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[16].__cell__  (.A(Di0[16]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[16].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[17].__cell__  (.A(Di0[17]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[17].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[18].__cell__  (.A(Di0[18]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[18].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[19].__cell__  (.A(Di0[19]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[19].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[1].__cell__  (.A(Di0[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[20].__cell__  (.A(Di0[20]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[20].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[21].__cell__  (.A(Di0[21]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[21].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[22].__cell__  (.A(Di0[22]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[22].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[23].__cell__  (.A(Di0[23]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[23].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[24].__cell__  (.A(Di0[24]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[24].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[25].__cell__  (.A(Di0[25]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[25].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[26].__cell__  (.A(Di0[26]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[26].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[27].__cell__  (.A(Di0[27]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[27].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[28].__cell__  (.A(Di0[28]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[28].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[29].__cell__  (.A(Di0[29]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[29].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[2].__cell__  (.A(Di0[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[30].__cell__  (.A(Di0[30]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[30].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[31].__cell__  (.A(Di0[31]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[31].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[32].__cell__  (.A(Di0[32]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[32].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[33].__cell__  (.A(Di0[33]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[33].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[34].__cell__  (.A(Di0[34]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[34].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[35].__cell__  (.A(Di0[35]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[35].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[36].__cell__  (.A(Di0[36]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[36].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[37].__cell__  (.A(Di0[37]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[37].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[38].__cell__  (.A(Di0[38]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[38].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[39].__cell__  (.A(Di0[39]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[39].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[3].__cell__  (.A(Di0[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[3].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[40].__cell__  (.A(Di0[40]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[40].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[41].__cell__  (.A(Di0[41]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[41].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[42].__cell__  (.A(Di0[42]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[42].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[43].__cell__  (.A(Di0[43]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[43].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[44].__cell__  (.A(Di0[44]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[44].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[45].__cell__  (.A(Di0[45]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[45].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[46].__cell__  (.A(Di0[46]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[46].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[47].__cell__  (.A(Di0[47]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[47].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[48].__cell__  (.A(Di0[48]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[48].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[49].__cell__  (.A(Di0[49]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[49].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[4].__cell__  (.A(Di0[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[4].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[50].__cell__  (.A(Di0[50]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[50].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[51].__cell__  (.A(Di0[51]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[51].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[52].__cell__  (.A(Di0[52]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[52].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[53].__cell__  (.A(Di0[53]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[53].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[54].__cell__  (.A(Di0[54]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[54].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[55].__cell__  (.A(Di0[55]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[55].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[56].__cell__  (.A(Di0[56]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[56].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[57].__cell__  (.A(Di0[57]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[57].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[58].__cell__  (.A(Di0[58]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[58].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[59].__cell__  (.A(Di0[59]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[59].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[5].__cell__  (.A(Di0[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[5].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[60].__cell__  (.A(Di0[60]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[60].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[61].__cell__  (.A(Di0[61]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[61].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[62].__cell__  (.A(Di0[62]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[62].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[63].__cell__  (.A(Di0[63]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[63].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[6].__cell__  (.A(Di0[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[6].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[7].__cell__  (.A(Di0[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[7].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[8].__cell__  (.A(Di0[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[8].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[9].__cell__  (.A(Di0[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[9].X ));
 sky130_fd_sc_hd__clkbuf_4 \Do0_REG.Do_CLKBUF[0]  (.A(\Do0_REG.CLK_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Do0_REG.CLKBUF[0] ));
 sky130_fd_sc_hd__clkbuf_4 \Do0_REG.Do_CLKBUF[1]  (.A(\Do0_REG.CLK_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Do0_REG.CLKBUF[1] ));
 sky130_fd_sc_hd__clkbuf_4 \Do0_REG.Do_CLKBUF[2]  (.A(\Do0_REG.CLK_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Do0_REG.CLKBUF[2] ));
 sky130_fd_sc_hd__clkbuf_4 \Do0_REG.Do_CLKBUF[3]  (.A(\Do0_REG.CLK_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Do0_REG.CLKBUF[3] ));
 sky130_fd_sc_hd__clkbuf_4 \Do0_REG.Do_CLKBUF[4]  (.A(\Do0_REG.CLK_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Do0_REG.CLKBUF[4] ));
 sky130_fd_sc_hd__clkbuf_4 \Do0_REG.Do_CLKBUF[5]  (.A(\Do0_REG.CLK_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Do0_REG.CLKBUF[5] ));
 sky130_fd_sc_hd__clkbuf_4 \Do0_REG.Do_CLKBUF[6]  (.A(\Do0_REG.CLK_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Do0_REG.CLKBUF[6] ));
 sky130_fd_sc_hd__clkbuf_4 \Do0_REG.Do_CLKBUF[7]  (.A(\Do0_REG.CLK_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Do0_REG.CLKBUF[7] ));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[0].DIODE[0]  (.DIODE(\BYTE[0].FLOATBUF0[0].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[0].DIODE[1]  (.DIODE(\BYTE[0].FLOATBUF0[1].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[0].DIODE[2]  (.DIODE(\BYTE[0].FLOATBUF0[2].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[0].DIODE[3]  (.DIODE(\BYTE[0].FLOATBUF0[3].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[0].DIODE[4]  (.DIODE(\BYTE[0].FLOATBUF0[4].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[0].DIODE[5]  (.DIODE(\BYTE[0].FLOATBUF0[5].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[0].DIODE[6]  (.DIODE(\BYTE[0].FLOATBUF0[6].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[0].DIODE[7]  (.DIODE(\BYTE[0].FLOATBUF0[7].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[0].Do_FF[0]  (.CLK(\Do0_REG.CLKBUF[0] ),
    .D(\BYTE[0].FLOATBUF0[0].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[0]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[0].Do_FF[1]  (.CLK(\Do0_REG.CLKBUF[0] ),
    .D(\BYTE[0].FLOATBUF0[1].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[1]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[0].Do_FF[2]  (.CLK(\Do0_REG.CLKBUF[0] ),
    .D(\BYTE[0].FLOATBUF0[2].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[2]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[0].Do_FF[3]  (.CLK(\Do0_REG.CLKBUF[0] ),
    .D(\BYTE[0].FLOATBUF0[3].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[3]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[0].Do_FF[4]  (.CLK(\Do0_REG.CLKBUF[0] ),
    .D(\BYTE[0].FLOATBUF0[4].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[4]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[0].Do_FF[5]  (.CLK(\Do0_REG.CLKBUF[0] ),
    .D(\BYTE[0].FLOATBUF0[5].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[5]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[0].Do_FF[6]  (.CLK(\Do0_REG.CLKBUF[0] ),
    .D(\BYTE[0].FLOATBUF0[6].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[6]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[0].Do_FF[7]  (.CLK(\Do0_REG.CLKBUF[0] ),
    .D(\BYTE[0].FLOATBUF0[7].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[7]));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[1].DIODE[0]  (.DIODE(\BYTE[1].FLOATBUF0[8].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[1].DIODE[1]  (.DIODE(\BYTE[1].FLOATBUF0[9].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[1].DIODE[2]  (.DIODE(\BYTE[1].FLOATBUF0[10].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[1].DIODE[3]  (.DIODE(\BYTE[1].FLOATBUF0[11].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[1].DIODE[4]  (.DIODE(\BYTE[1].FLOATBUF0[12].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[1].DIODE[5]  (.DIODE(\BYTE[1].FLOATBUF0[13].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[1].DIODE[6]  (.DIODE(\BYTE[1].FLOATBUF0[14].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[1].DIODE[7]  (.DIODE(\BYTE[1].FLOATBUF0[15].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[1].Do_FF[0]  (.CLK(\Do0_REG.CLKBUF[1] ),
    .D(\BYTE[1].FLOATBUF0[8].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[8]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[1].Do_FF[1]  (.CLK(\Do0_REG.CLKBUF[1] ),
    .D(\BYTE[1].FLOATBUF0[9].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[9]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[1].Do_FF[2]  (.CLK(\Do0_REG.CLKBUF[1] ),
    .D(\BYTE[1].FLOATBUF0[10].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[10]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[1].Do_FF[3]  (.CLK(\Do0_REG.CLKBUF[1] ),
    .D(\BYTE[1].FLOATBUF0[11].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[11]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[1].Do_FF[4]  (.CLK(\Do0_REG.CLKBUF[1] ),
    .D(\BYTE[1].FLOATBUF0[12].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[12]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[1].Do_FF[5]  (.CLK(\Do0_REG.CLKBUF[1] ),
    .D(\BYTE[1].FLOATBUF0[13].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[13]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[1].Do_FF[6]  (.CLK(\Do0_REG.CLKBUF[1] ),
    .D(\BYTE[1].FLOATBUF0[14].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[14]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[1].Do_FF[7]  (.CLK(\Do0_REG.CLKBUF[1] ),
    .D(\BYTE[1].FLOATBUF0[15].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[15]));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[2].DIODE[0]  (.DIODE(\BYTE[2].FLOATBUF0[16].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[2].DIODE[1]  (.DIODE(\BYTE[2].FLOATBUF0[17].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[2].DIODE[2]  (.DIODE(\BYTE[2].FLOATBUF0[18].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[2].DIODE[3]  (.DIODE(\BYTE[2].FLOATBUF0[19].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[2].DIODE[4]  (.DIODE(\BYTE[2].FLOATBUF0[20].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[2].DIODE[5]  (.DIODE(\BYTE[2].FLOATBUF0[21].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[2].DIODE[6]  (.DIODE(\BYTE[2].FLOATBUF0[22].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[2].DIODE[7]  (.DIODE(\BYTE[2].FLOATBUF0[23].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[2].Do_FF[0]  (.CLK(\Do0_REG.CLKBUF[2] ),
    .D(\BYTE[2].FLOATBUF0[16].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[16]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[2].Do_FF[1]  (.CLK(\Do0_REG.CLKBUF[2] ),
    .D(\BYTE[2].FLOATBUF0[17].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[17]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[2].Do_FF[2]  (.CLK(\Do0_REG.CLKBUF[2] ),
    .D(\BYTE[2].FLOATBUF0[18].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[18]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[2].Do_FF[3]  (.CLK(\Do0_REG.CLKBUF[2] ),
    .D(\BYTE[2].FLOATBUF0[19].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[19]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[2].Do_FF[4]  (.CLK(\Do0_REG.CLKBUF[2] ),
    .D(\BYTE[2].FLOATBUF0[20].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[20]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[2].Do_FF[5]  (.CLK(\Do0_REG.CLKBUF[2] ),
    .D(\BYTE[2].FLOATBUF0[21].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[21]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[2].Do_FF[6]  (.CLK(\Do0_REG.CLKBUF[2] ),
    .D(\BYTE[2].FLOATBUF0[22].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[22]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[2].Do_FF[7]  (.CLK(\Do0_REG.CLKBUF[2] ),
    .D(\BYTE[2].FLOATBUF0[23].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[23]));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[3].DIODE[0]  (.DIODE(\BYTE[3].FLOATBUF0[24].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[3].DIODE[1]  (.DIODE(\BYTE[3].FLOATBUF0[25].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[3].DIODE[2]  (.DIODE(\BYTE[3].FLOATBUF0[26].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[3].DIODE[3]  (.DIODE(\BYTE[3].FLOATBUF0[27].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[3].DIODE[4]  (.DIODE(\BYTE[3].FLOATBUF0[28].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[3].DIODE[5]  (.DIODE(\BYTE[3].FLOATBUF0[29].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[3].DIODE[6]  (.DIODE(\BYTE[3].FLOATBUF0[30].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[3].DIODE[7]  (.DIODE(\BYTE[3].FLOATBUF0[31].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[3].Do_FF[0]  (.CLK(\Do0_REG.CLKBUF[3] ),
    .D(\BYTE[3].FLOATBUF0[24].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[24]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[3].Do_FF[1]  (.CLK(\Do0_REG.CLKBUF[3] ),
    .D(\BYTE[3].FLOATBUF0[25].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[25]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[3].Do_FF[2]  (.CLK(\Do0_REG.CLKBUF[3] ),
    .D(\BYTE[3].FLOATBUF0[26].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[26]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[3].Do_FF[3]  (.CLK(\Do0_REG.CLKBUF[3] ),
    .D(\BYTE[3].FLOATBUF0[27].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[27]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[3].Do_FF[4]  (.CLK(\Do0_REG.CLKBUF[3] ),
    .D(\BYTE[3].FLOATBUF0[28].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[28]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[3].Do_FF[5]  (.CLK(\Do0_REG.CLKBUF[3] ),
    .D(\BYTE[3].FLOATBUF0[29].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[29]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[3].Do_FF[6]  (.CLK(\Do0_REG.CLKBUF[3] ),
    .D(\BYTE[3].FLOATBUF0[30].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[30]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[3].Do_FF[7]  (.CLK(\Do0_REG.CLKBUF[3] ),
    .D(\BYTE[3].FLOATBUF0[31].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[31]));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[4].DIODE[0]  (.DIODE(\BYTE[4].FLOATBUF0[32].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[4].DIODE[1]  (.DIODE(\BYTE[4].FLOATBUF0[33].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[4].DIODE[2]  (.DIODE(\BYTE[4].FLOATBUF0[34].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[4].DIODE[3]  (.DIODE(\BYTE[4].FLOATBUF0[35].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[4].DIODE[4]  (.DIODE(\BYTE[4].FLOATBUF0[36].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[4].DIODE[5]  (.DIODE(\BYTE[4].FLOATBUF0[37].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[4].DIODE[6]  (.DIODE(\BYTE[4].FLOATBUF0[38].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[4].DIODE[7]  (.DIODE(\BYTE[4].FLOATBUF0[39].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[4].Do_FF[0]  (.CLK(\Do0_REG.CLKBUF[4] ),
    .D(\BYTE[4].FLOATBUF0[32].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[32]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[4].Do_FF[1]  (.CLK(\Do0_REG.CLKBUF[4] ),
    .D(\BYTE[4].FLOATBUF0[33].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[33]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[4].Do_FF[2]  (.CLK(\Do0_REG.CLKBUF[4] ),
    .D(\BYTE[4].FLOATBUF0[34].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[34]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[4].Do_FF[3]  (.CLK(\Do0_REG.CLKBUF[4] ),
    .D(\BYTE[4].FLOATBUF0[35].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[35]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[4].Do_FF[4]  (.CLK(\Do0_REG.CLKBUF[4] ),
    .D(\BYTE[4].FLOATBUF0[36].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[36]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[4].Do_FF[5]  (.CLK(\Do0_REG.CLKBUF[4] ),
    .D(\BYTE[4].FLOATBUF0[37].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[37]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[4].Do_FF[6]  (.CLK(\Do0_REG.CLKBUF[4] ),
    .D(\BYTE[4].FLOATBUF0[38].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[38]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[4].Do_FF[7]  (.CLK(\Do0_REG.CLKBUF[4] ),
    .D(\BYTE[4].FLOATBUF0[39].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[39]));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[5].DIODE[0]  (.DIODE(\BYTE[5].FLOATBUF0[40].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[5].DIODE[1]  (.DIODE(\BYTE[5].FLOATBUF0[41].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[5].DIODE[2]  (.DIODE(\BYTE[5].FLOATBUF0[42].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[5].DIODE[3]  (.DIODE(\BYTE[5].FLOATBUF0[43].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[5].DIODE[4]  (.DIODE(\BYTE[5].FLOATBUF0[44].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[5].DIODE[5]  (.DIODE(\BYTE[5].FLOATBUF0[45].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[5].DIODE[6]  (.DIODE(\BYTE[5].FLOATBUF0[46].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[5].DIODE[7]  (.DIODE(\BYTE[5].FLOATBUF0[47].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[5].Do_FF[0]  (.CLK(\Do0_REG.CLKBUF[5] ),
    .D(\BYTE[5].FLOATBUF0[40].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[40]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[5].Do_FF[1]  (.CLK(\Do0_REG.CLKBUF[5] ),
    .D(\BYTE[5].FLOATBUF0[41].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[41]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[5].Do_FF[2]  (.CLK(\Do0_REG.CLKBUF[5] ),
    .D(\BYTE[5].FLOATBUF0[42].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[42]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[5].Do_FF[3]  (.CLK(\Do0_REG.CLKBUF[5] ),
    .D(\BYTE[5].FLOATBUF0[43].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[43]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[5].Do_FF[4]  (.CLK(\Do0_REG.CLKBUF[5] ),
    .D(\BYTE[5].FLOATBUF0[44].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[44]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[5].Do_FF[5]  (.CLK(\Do0_REG.CLKBUF[5] ),
    .D(\BYTE[5].FLOATBUF0[45].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[45]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[5].Do_FF[6]  (.CLK(\Do0_REG.CLKBUF[5] ),
    .D(\BYTE[5].FLOATBUF0[46].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[46]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[5].Do_FF[7]  (.CLK(\Do0_REG.CLKBUF[5] ),
    .D(\BYTE[5].FLOATBUF0[47].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[47]));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[6].DIODE[0]  (.DIODE(\BYTE[6].FLOATBUF0[48].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[6].DIODE[1]  (.DIODE(\BYTE[6].FLOATBUF0[49].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[6].DIODE[2]  (.DIODE(\BYTE[6].FLOATBUF0[50].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[6].DIODE[3]  (.DIODE(\BYTE[6].FLOATBUF0[51].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[6].DIODE[4]  (.DIODE(\BYTE[6].FLOATBUF0[52].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[6].DIODE[5]  (.DIODE(\BYTE[6].FLOATBUF0[53].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[6].DIODE[6]  (.DIODE(\BYTE[6].FLOATBUF0[54].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[6].DIODE[7]  (.DIODE(\BYTE[6].FLOATBUF0[55].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[6].Do_FF[0]  (.CLK(\Do0_REG.CLKBUF[6] ),
    .D(\BYTE[6].FLOATBUF0[48].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[48]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[6].Do_FF[1]  (.CLK(\Do0_REG.CLKBUF[6] ),
    .D(\BYTE[6].FLOATBUF0[49].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[49]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[6].Do_FF[2]  (.CLK(\Do0_REG.CLKBUF[6] ),
    .D(\BYTE[6].FLOATBUF0[50].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[50]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[6].Do_FF[3]  (.CLK(\Do0_REG.CLKBUF[6] ),
    .D(\BYTE[6].FLOATBUF0[51].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[51]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[6].Do_FF[4]  (.CLK(\Do0_REG.CLKBUF[6] ),
    .D(\BYTE[6].FLOATBUF0[52].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[52]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[6].Do_FF[5]  (.CLK(\Do0_REG.CLKBUF[6] ),
    .D(\BYTE[6].FLOATBUF0[53].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[53]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[6].Do_FF[6]  (.CLK(\Do0_REG.CLKBUF[6] ),
    .D(\BYTE[6].FLOATBUF0[54].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[54]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[6].Do_FF[7]  (.CLK(\Do0_REG.CLKBUF[6] ),
    .D(\BYTE[6].FLOATBUF0[55].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[55]));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[7].DIODE[0]  (.DIODE(\BYTE[7].FLOATBUF0[56].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[7].DIODE[1]  (.DIODE(\BYTE[7].FLOATBUF0[57].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[7].DIODE[2]  (.DIODE(\BYTE[7].FLOATBUF0[58].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[7].DIODE[3]  (.DIODE(\BYTE[7].FLOATBUF0[59].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[7].DIODE[4]  (.DIODE(\BYTE[7].FLOATBUF0[60].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[7].DIODE[5]  (.DIODE(\BYTE[7].FLOATBUF0[61].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[7].DIODE[6]  (.DIODE(\BYTE[7].FLOATBUF0[62].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0_REG.OUTREG_BYTE[7].DIODE[7]  (.DIODE(\BYTE[7].FLOATBUF0[63].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[7].Do_FF[0]  (.CLK(\Do0_REG.CLKBUF[7] ),
    .D(\BYTE[7].FLOATBUF0[56].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[56]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[7].Do_FF[1]  (.CLK(\Do0_REG.CLKBUF[7] ),
    .D(\BYTE[7].FLOATBUF0[57].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[57]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[7].Do_FF[2]  (.CLK(\Do0_REG.CLKBUF[7] ),
    .D(\BYTE[7].FLOATBUF0[58].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[58]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[7].Do_FF[3]  (.CLK(\Do0_REG.CLKBUF[7] ),
    .D(\BYTE[7].FLOATBUF0[59].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[59]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[7].Do_FF[4]  (.CLK(\Do0_REG.CLKBUF[7] ),
    .D(\BYTE[7].FLOATBUF0[60].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[60]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[7].Do_FF[5]  (.CLK(\Do0_REG.CLKBUF[7] ),
    .D(\BYTE[7].FLOATBUF0[61].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[61]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[7].Do_FF[6]  (.CLK(\Do0_REG.CLKBUF[7] ),
    .D(\BYTE[7].FLOATBUF0[62].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[62]));
 sky130_fd_sc_hd__dfxtp_1 \Do0_REG.OUTREG_BYTE[7].Do_FF[7]  (.CLK(\Do0_REG.CLKBUF[7] ),
    .D(\BYTE[7].FLOATBUF0[63].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do0[63]));
 sky130_fd_sc_hd__clkbuf_4 \Do0_REG.Root_CLKBUF  (.A(\CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Do0_REG.CLK_buf ));
 sky130_fd_sc_hd__clkbuf_4 \Do1_REG.Do_CLKBUF[0]  (.A(\Do1_REG.CLK_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Do1_REG.CLKBUF[0] ));
 sky130_fd_sc_hd__clkbuf_4 \Do1_REG.Do_CLKBUF[1]  (.A(\Do1_REG.CLK_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Do1_REG.CLKBUF[1] ));
 sky130_fd_sc_hd__clkbuf_4 \Do1_REG.Do_CLKBUF[2]  (.A(\Do1_REG.CLK_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Do1_REG.CLKBUF[2] ));
 sky130_fd_sc_hd__clkbuf_4 \Do1_REG.Do_CLKBUF[3]  (.A(\Do1_REG.CLK_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Do1_REG.CLKBUF[3] ));
 sky130_fd_sc_hd__clkbuf_4 \Do1_REG.Do_CLKBUF[4]  (.A(\Do1_REG.CLK_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Do1_REG.CLKBUF[4] ));
 sky130_fd_sc_hd__clkbuf_4 \Do1_REG.Do_CLKBUF[5]  (.A(\Do1_REG.CLK_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Do1_REG.CLKBUF[5] ));
 sky130_fd_sc_hd__clkbuf_4 \Do1_REG.Do_CLKBUF[6]  (.A(\Do1_REG.CLK_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Do1_REG.CLKBUF[6] ));
 sky130_fd_sc_hd__clkbuf_4 \Do1_REG.Do_CLKBUF[7]  (.A(\Do1_REG.CLK_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Do1_REG.CLKBUF[7] ));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[0].DIODE[0]  (.DIODE(\BYTE[0].FLOATBUF1[0].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[0].DIODE[1]  (.DIODE(\BYTE[0].FLOATBUF1[1].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[0].DIODE[2]  (.DIODE(\BYTE[0].FLOATBUF1[2].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[0].DIODE[3]  (.DIODE(\BYTE[0].FLOATBUF1[3].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[0].DIODE[4]  (.DIODE(\BYTE[0].FLOATBUF1[4].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[0].DIODE[5]  (.DIODE(\BYTE[0].FLOATBUF1[5].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[0].DIODE[6]  (.DIODE(\BYTE[0].FLOATBUF1[6].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[0].DIODE[7]  (.DIODE(\BYTE[0].FLOATBUF1[7].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[0].Do_FF[0]  (.CLK(\Do1_REG.CLKBUF[0] ),
    .D(\BYTE[0].FLOATBUF1[0].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[0]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[0].Do_FF[1]  (.CLK(\Do1_REG.CLKBUF[0] ),
    .D(\BYTE[0].FLOATBUF1[1].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[1]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[0].Do_FF[2]  (.CLK(\Do1_REG.CLKBUF[0] ),
    .D(\BYTE[0].FLOATBUF1[2].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[2]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[0].Do_FF[3]  (.CLK(\Do1_REG.CLKBUF[0] ),
    .D(\BYTE[0].FLOATBUF1[3].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[3]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[0].Do_FF[4]  (.CLK(\Do1_REG.CLKBUF[0] ),
    .D(\BYTE[0].FLOATBUF1[4].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[4]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[0].Do_FF[5]  (.CLK(\Do1_REG.CLKBUF[0] ),
    .D(\BYTE[0].FLOATBUF1[5].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[5]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[0].Do_FF[6]  (.CLK(\Do1_REG.CLKBUF[0] ),
    .D(\BYTE[0].FLOATBUF1[6].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[6]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[0].Do_FF[7]  (.CLK(\Do1_REG.CLKBUF[0] ),
    .D(\BYTE[0].FLOATBUF1[7].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[7]));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[1].DIODE[0]  (.DIODE(\BYTE[1].FLOATBUF1[8].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[1].DIODE[1]  (.DIODE(\BYTE[1].FLOATBUF1[9].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[1].DIODE[2]  (.DIODE(\BYTE[1].FLOATBUF1[10].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[1].DIODE[3]  (.DIODE(\BYTE[1].FLOATBUF1[11].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[1].DIODE[4]  (.DIODE(\BYTE[1].FLOATBUF1[12].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[1].DIODE[5]  (.DIODE(\BYTE[1].FLOATBUF1[13].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[1].DIODE[6]  (.DIODE(\BYTE[1].FLOATBUF1[14].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[1].DIODE[7]  (.DIODE(\BYTE[1].FLOATBUF1[15].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[1].Do_FF[0]  (.CLK(\Do1_REG.CLKBUF[1] ),
    .D(\BYTE[1].FLOATBUF1[8].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[8]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[1].Do_FF[1]  (.CLK(\Do1_REG.CLKBUF[1] ),
    .D(\BYTE[1].FLOATBUF1[9].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[9]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[1].Do_FF[2]  (.CLK(\Do1_REG.CLKBUF[1] ),
    .D(\BYTE[1].FLOATBUF1[10].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[10]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[1].Do_FF[3]  (.CLK(\Do1_REG.CLKBUF[1] ),
    .D(\BYTE[1].FLOATBUF1[11].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[11]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[1].Do_FF[4]  (.CLK(\Do1_REG.CLKBUF[1] ),
    .D(\BYTE[1].FLOATBUF1[12].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[12]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[1].Do_FF[5]  (.CLK(\Do1_REG.CLKBUF[1] ),
    .D(\BYTE[1].FLOATBUF1[13].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[13]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[1].Do_FF[6]  (.CLK(\Do1_REG.CLKBUF[1] ),
    .D(\BYTE[1].FLOATBUF1[14].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[14]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[1].Do_FF[7]  (.CLK(\Do1_REG.CLKBUF[1] ),
    .D(\BYTE[1].FLOATBUF1[15].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[15]));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[2].DIODE[0]  (.DIODE(\BYTE[2].FLOATBUF1[16].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[2].DIODE[1]  (.DIODE(\BYTE[2].FLOATBUF1[17].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[2].DIODE[2]  (.DIODE(\BYTE[2].FLOATBUF1[18].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[2].DIODE[3]  (.DIODE(\BYTE[2].FLOATBUF1[19].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[2].DIODE[4]  (.DIODE(\BYTE[2].FLOATBUF1[20].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[2].DIODE[5]  (.DIODE(\BYTE[2].FLOATBUF1[21].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[2].DIODE[6]  (.DIODE(\BYTE[2].FLOATBUF1[22].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[2].DIODE[7]  (.DIODE(\BYTE[2].FLOATBUF1[23].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[2].Do_FF[0]  (.CLK(\Do1_REG.CLKBUF[2] ),
    .D(\BYTE[2].FLOATBUF1[16].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[16]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[2].Do_FF[1]  (.CLK(\Do1_REG.CLKBUF[2] ),
    .D(\BYTE[2].FLOATBUF1[17].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[17]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[2].Do_FF[2]  (.CLK(\Do1_REG.CLKBUF[2] ),
    .D(\BYTE[2].FLOATBUF1[18].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[18]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[2].Do_FF[3]  (.CLK(\Do1_REG.CLKBUF[2] ),
    .D(\BYTE[2].FLOATBUF1[19].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[19]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[2].Do_FF[4]  (.CLK(\Do1_REG.CLKBUF[2] ),
    .D(\BYTE[2].FLOATBUF1[20].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[20]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[2].Do_FF[5]  (.CLK(\Do1_REG.CLKBUF[2] ),
    .D(\BYTE[2].FLOATBUF1[21].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[21]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[2].Do_FF[6]  (.CLK(\Do1_REG.CLKBUF[2] ),
    .D(\BYTE[2].FLOATBUF1[22].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[22]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[2].Do_FF[7]  (.CLK(\Do1_REG.CLKBUF[2] ),
    .D(\BYTE[2].FLOATBUF1[23].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[23]));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[3].DIODE[0]  (.DIODE(\BYTE[3].FLOATBUF1[24].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[3].DIODE[1]  (.DIODE(\BYTE[3].FLOATBUF1[25].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[3].DIODE[2]  (.DIODE(\BYTE[3].FLOATBUF1[26].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[3].DIODE[3]  (.DIODE(\BYTE[3].FLOATBUF1[27].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[3].DIODE[4]  (.DIODE(\BYTE[3].FLOATBUF1[28].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[3].DIODE[5]  (.DIODE(\BYTE[3].FLOATBUF1[29].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[3].DIODE[6]  (.DIODE(\BYTE[3].FLOATBUF1[30].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[3].DIODE[7]  (.DIODE(\BYTE[3].FLOATBUF1[31].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[3].Do_FF[0]  (.CLK(\Do1_REG.CLKBUF[3] ),
    .D(\BYTE[3].FLOATBUF1[24].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[24]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[3].Do_FF[1]  (.CLK(\Do1_REG.CLKBUF[3] ),
    .D(\BYTE[3].FLOATBUF1[25].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[25]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[3].Do_FF[2]  (.CLK(\Do1_REG.CLKBUF[3] ),
    .D(\BYTE[3].FLOATBUF1[26].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[26]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[3].Do_FF[3]  (.CLK(\Do1_REG.CLKBUF[3] ),
    .D(\BYTE[3].FLOATBUF1[27].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[27]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[3].Do_FF[4]  (.CLK(\Do1_REG.CLKBUF[3] ),
    .D(\BYTE[3].FLOATBUF1[28].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[28]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[3].Do_FF[5]  (.CLK(\Do1_REG.CLKBUF[3] ),
    .D(\BYTE[3].FLOATBUF1[29].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[29]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[3].Do_FF[6]  (.CLK(\Do1_REG.CLKBUF[3] ),
    .D(\BYTE[3].FLOATBUF1[30].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[30]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[3].Do_FF[7]  (.CLK(\Do1_REG.CLKBUF[3] ),
    .D(\BYTE[3].FLOATBUF1[31].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[31]));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[4].DIODE[0]  (.DIODE(\BYTE[4].FLOATBUF1[32].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[4].DIODE[1]  (.DIODE(\BYTE[4].FLOATBUF1[33].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[4].DIODE[2]  (.DIODE(\BYTE[4].FLOATBUF1[34].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[4].DIODE[3]  (.DIODE(\BYTE[4].FLOATBUF1[35].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[4].DIODE[4]  (.DIODE(\BYTE[4].FLOATBUF1[36].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[4].DIODE[5]  (.DIODE(\BYTE[4].FLOATBUF1[37].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[4].DIODE[6]  (.DIODE(\BYTE[4].FLOATBUF1[38].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[4].DIODE[7]  (.DIODE(\BYTE[4].FLOATBUF1[39].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[4].Do_FF[0]  (.CLK(\Do1_REG.CLKBUF[4] ),
    .D(\BYTE[4].FLOATBUF1[32].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[32]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[4].Do_FF[1]  (.CLK(\Do1_REG.CLKBUF[4] ),
    .D(\BYTE[4].FLOATBUF1[33].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[33]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[4].Do_FF[2]  (.CLK(\Do1_REG.CLKBUF[4] ),
    .D(\BYTE[4].FLOATBUF1[34].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[34]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[4].Do_FF[3]  (.CLK(\Do1_REG.CLKBUF[4] ),
    .D(\BYTE[4].FLOATBUF1[35].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[35]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[4].Do_FF[4]  (.CLK(\Do1_REG.CLKBUF[4] ),
    .D(\BYTE[4].FLOATBUF1[36].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[36]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[4].Do_FF[5]  (.CLK(\Do1_REG.CLKBUF[4] ),
    .D(\BYTE[4].FLOATBUF1[37].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[37]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[4].Do_FF[6]  (.CLK(\Do1_REG.CLKBUF[4] ),
    .D(\BYTE[4].FLOATBUF1[38].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[38]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[4].Do_FF[7]  (.CLK(\Do1_REG.CLKBUF[4] ),
    .D(\BYTE[4].FLOATBUF1[39].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[39]));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[5].DIODE[0]  (.DIODE(\BYTE[5].FLOATBUF1[40].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[5].DIODE[1]  (.DIODE(\BYTE[5].FLOATBUF1[41].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[5].DIODE[2]  (.DIODE(\BYTE[5].FLOATBUF1[42].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[5].DIODE[3]  (.DIODE(\BYTE[5].FLOATBUF1[43].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[5].DIODE[4]  (.DIODE(\BYTE[5].FLOATBUF1[44].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[5].DIODE[5]  (.DIODE(\BYTE[5].FLOATBUF1[45].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[5].DIODE[6]  (.DIODE(\BYTE[5].FLOATBUF1[46].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[5].DIODE[7]  (.DIODE(\BYTE[5].FLOATBUF1[47].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[5].Do_FF[0]  (.CLK(\Do1_REG.CLKBUF[5] ),
    .D(\BYTE[5].FLOATBUF1[40].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[40]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[5].Do_FF[1]  (.CLK(\Do1_REG.CLKBUF[5] ),
    .D(\BYTE[5].FLOATBUF1[41].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[41]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[5].Do_FF[2]  (.CLK(\Do1_REG.CLKBUF[5] ),
    .D(\BYTE[5].FLOATBUF1[42].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[42]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[5].Do_FF[3]  (.CLK(\Do1_REG.CLKBUF[5] ),
    .D(\BYTE[5].FLOATBUF1[43].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[43]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[5].Do_FF[4]  (.CLK(\Do1_REG.CLKBUF[5] ),
    .D(\BYTE[5].FLOATBUF1[44].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[44]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[5].Do_FF[5]  (.CLK(\Do1_REG.CLKBUF[5] ),
    .D(\BYTE[5].FLOATBUF1[45].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[45]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[5].Do_FF[6]  (.CLK(\Do1_REG.CLKBUF[5] ),
    .D(\BYTE[5].FLOATBUF1[46].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[46]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[5].Do_FF[7]  (.CLK(\Do1_REG.CLKBUF[5] ),
    .D(\BYTE[5].FLOATBUF1[47].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[47]));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[6].DIODE[0]  (.DIODE(\BYTE[6].FLOATBUF1[48].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[6].DIODE[1]  (.DIODE(\BYTE[6].FLOATBUF1[49].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[6].DIODE[2]  (.DIODE(\BYTE[6].FLOATBUF1[50].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[6].DIODE[3]  (.DIODE(\BYTE[6].FLOATBUF1[51].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[6].DIODE[4]  (.DIODE(\BYTE[6].FLOATBUF1[52].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[6].DIODE[5]  (.DIODE(\BYTE[6].FLOATBUF1[53].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[6].DIODE[6]  (.DIODE(\BYTE[6].FLOATBUF1[54].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[6].DIODE[7]  (.DIODE(\BYTE[6].FLOATBUF1[55].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[6].Do_FF[0]  (.CLK(\Do1_REG.CLKBUF[6] ),
    .D(\BYTE[6].FLOATBUF1[48].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[48]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[6].Do_FF[1]  (.CLK(\Do1_REG.CLKBUF[6] ),
    .D(\BYTE[6].FLOATBUF1[49].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[49]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[6].Do_FF[2]  (.CLK(\Do1_REG.CLKBUF[6] ),
    .D(\BYTE[6].FLOATBUF1[50].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[50]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[6].Do_FF[3]  (.CLK(\Do1_REG.CLKBUF[6] ),
    .D(\BYTE[6].FLOATBUF1[51].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[51]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[6].Do_FF[4]  (.CLK(\Do1_REG.CLKBUF[6] ),
    .D(\BYTE[6].FLOATBUF1[52].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[52]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[6].Do_FF[5]  (.CLK(\Do1_REG.CLKBUF[6] ),
    .D(\BYTE[6].FLOATBUF1[53].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[53]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[6].Do_FF[6]  (.CLK(\Do1_REG.CLKBUF[6] ),
    .D(\BYTE[6].FLOATBUF1[54].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[54]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[6].Do_FF[7]  (.CLK(\Do1_REG.CLKBUF[6] ),
    .D(\BYTE[6].FLOATBUF1[55].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[55]));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[7].DIODE[0]  (.DIODE(\BYTE[7].FLOATBUF1[56].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[7].DIODE[1]  (.DIODE(\BYTE[7].FLOATBUF1[57].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[7].DIODE[2]  (.DIODE(\BYTE[7].FLOATBUF1[58].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[7].DIODE[3]  (.DIODE(\BYTE[7].FLOATBUF1[59].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[7].DIODE[4]  (.DIODE(\BYTE[7].FLOATBUF1[60].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[7].DIODE[5]  (.DIODE(\BYTE[7].FLOATBUF1[61].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[7].DIODE[6]  (.DIODE(\BYTE[7].FLOATBUF1[62].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do1_REG.OUTREG_BYTE[7].DIODE[7]  (.DIODE(\BYTE[7].FLOATBUF1[63].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[7].Do_FF[0]  (.CLK(\Do1_REG.CLKBUF[7] ),
    .D(\BYTE[7].FLOATBUF1[56].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[56]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[7].Do_FF[1]  (.CLK(\Do1_REG.CLKBUF[7] ),
    .D(\BYTE[7].FLOATBUF1[57].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[57]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[7].Do_FF[2]  (.CLK(\Do1_REG.CLKBUF[7] ),
    .D(\BYTE[7].FLOATBUF1[58].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[58]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[7].Do_FF[3]  (.CLK(\Do1_REG.CLKBUF[7] ),
    .D(\BYTE[7].FLOATBUF1[59].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[59]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[7].Do_FF[4]  (.CLK(\Do1_REG.CLKBUF[7] ),
    .D(\BYTE[7].FLOATBUF1[60].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[60]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[7].Do_FF[5]  (.CLK(\Do1_REG.CLKBUF[7] ),
    .D(\BYTE[7].FLOATBUF1[61].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[61]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[7].Do_FF[6]  (.CLK(\Do1_REG.CLKBUF[7] ),
    .D(\BYTE[7].FLOATBUF1[62].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[62]));
 sky130_fd_sc_hd__dfxtp_1 \Do1_REG.OUTREG_BYTE[7].Do_FF[7]  (.CLK(\Do1_REG.CLKBUF[7] ),
    .D(\BYTE[7].FLOATBUF1[63].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Do1[63]));
 sky130_fd_sc_hd__clkbuf_4 \Do1_REG.Root_CLKBUF  (.A(\CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Do1_REG.CLK_buf ));
 sky130_fd_sc_hd__clkbuf_2 \EN0BUF.__cell__  (.A(EN0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \EN1BUF.__cell__  (.A(EN1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DEC1.EN ));
 sky130_fd_sc_hd__clkbuf_2 \FBUFENBUF0[0].__cell__  (.A(EN0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\BYTE[0].FLOATBUF0[0].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \FBUFENBUF0[1].__cell__  (.A(EN0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\BYTE[1].FLOATBUF0[10].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \FBUFENBUF0[2].__cell__  (.A(EN0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\BYTE[2].FLOATBUF0[16].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \FBUFENBUF0[3].__cell__  (.A(EN0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\BYTE[3].FLOATBUF0[24].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \FBUFENBUF0[4].__cell__  (.A(EN0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\BYTE[4].FLOATBUF0[32].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \FBUFENBUF0[5].__cell__  (.A(EN0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\BYTE[5].FLOATBUF0[40].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \FBUFENBUF0[6].__cell__  (.A(EN0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\BYTE[6].FLOATBUF0[48].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \FBUFENBUF0[7].__cell__  (.A(EN0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\BYTE[7].FLOATBUF0[56].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \FBUFENBUF1[0].__cell__  (.A(EN1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\BYTE[0].FLOATBUF1[0].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \FBUFENBUF1[1].__cell__  (.A(EN1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\BYTE[1].FLOATBUF1[10].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \FBUFENBUF1[2].__cell__  (.A(EN1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\BYTE[2].FLOATBUF1[16].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \FBUFENBUF1[3].__cell__  (.A(EN1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\BYTE[3].FLOATBUF1[24].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \FBUFENBUF1[4].__cell__  (.A(EN1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\BYTE[4].FLOATBUF1[32].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \FBUFENBUF1[5].__cell__  (.A(EN1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\BYTE[5].FLOATBUF1[40].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \FBUFENBUF1[6].__cell__  (.A(EN1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\BYTE[6].FLOATBUF1[48].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \FBUFENBUF1[7].__cell__  (.A(EN1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\BYTE[7].FLOATBUF1[56].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.CLKBUF.__cell__  (.A(\CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.DEC0.ABUF[0]  (.A(\A0BUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.DEC0.ABUF[1]  (.A(\A0BUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.DEC0.ABUF[2]  (.A(\A0BUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \SLICE[0].RAM8.DEC0.AND0  (.A(\SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D_N(\SLICE[0].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE[0].RAM8.DEC0.AND1  (.A_N(\SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\SLICE[0].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE[0].RAM8.DEC0.AND2  (.A_N(\SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\SLICE[0].RAM8.DEC0.A_buf[1] ),
    .D(\SLICE[0].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \SLICE[0].RAM8.DEC0.AND3  (.A_N(\SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B(\SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\SLICE[0].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE[0].RAM8.DEC0.AND4  (.A_N(\SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B_N(\SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE[0].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \SLICE[0].RAM8.DEC0.AND5  (.A_N(\SLICE[0].RAM8.DEC0.A_buf[1] ),
    .B(\SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE[0].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \SLICE[0].RAM8.DEC0.AND6  (.A_N(\SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE[0].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \SLICE[0].RAM8.DEC0.AND7  (.A(\SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE[0].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.DEC0.ENBUF  (.A(\SLICE[0].RAM8.DEC0.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.DEC1.ABUF[0]  (.A(\A1BUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.DEC1.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.DEC1.ABUF[1]  (.A(\A1BUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.DEC1.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.DEC1.ABUF[2]  (.A(\A1BUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.DEC1.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \SLICE[0].RAM8.DEC1.AND0  (.A(\SLICE[0].RAM8.DEC1.A_buf[0] ),
    .B(\SLICE[0].RAM8.DEC1.A_buf[1] ),
    .C(\SLICE[0].RAM8.DEC1.A_buf[2] ),
    .D_N(\SLICE[0].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[0].W.SEL1 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE[0].RAM8.DEC1.AND1  (.A_N(\SLICE[0].RAM8.DEC1.A_buf[2] ),
    .B_N(\SLICE[0].RAM8.DEC1.A_buf[1] ),
    .C(\SLICE[0].RAM8.DEC1.A_buf[0] ),
    .D(\SLICE[0].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[1].W.SEL1 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE[0].RAM8.DEC1.AND2  (.A_N(\SLICE[0].RAM8.DEC1.A_buf[2] ),
    .B_N(\SLICE[0].RAM8.DEC1.A_buf[0] ),
    .C(\SLICE[0].RAM8.DEC1.A_buf[1] ),
    .D(\SLICE[0].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[2].W.SEL1 ));
 sky130_fd_sc_hd__and4b_2 \SLICE[0].RAM8.DEC1.AND3  (.A_N(\SLICE[0].RAM8.DEC1.A_buf[2] ),
    .B(\SLICE[0].RAM8.DEC1.A_buf[1] ),
    .C(\SLICE[0].RAM8.DEC1.A_buf[0] ),
    .D(\SLICE[0].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[3].W.SEL1 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE[0].RAM8.DEC1.AND4  (.A_N(\SLICE[0].RAM8.DEC1.A_buf[0] ),
    .B_N(\SLICE[0].RAM8.DEC1.A_buf[1] ),
    .C(\SLICE[0].RAM8.DEC1.A_buf[2] ),
    .D(\SLICE[0].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[4].W.SEL1 ));
 sky130_fd_sc_hd__and4b_2 \SLICE[0].RAM8.DEC1.AND5  (.A_N(\SLICE[0].RAM8.DEC1.A_buf[1] ),
    .B(\SLICE[0].RAM8.DEC1.A_buf[0] ),
    .C(\SLICE[0].RAM8.DEC1.A_buf[2] ),
    .D(\SLICE[0].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[5].W.SEL1 ));
 sky130_fd_sc_hd__and4b_2 \SLICE[0].RAM8.DEC1.AND6  (.A_N(\SLICE[0].RAM8.DEC1.A_buf[0] ),
    .B(\SLICE[0].RAM8.DEC1.A_buf[1] ),
    .C(\SLICE[0].RAM8.DEC1.A_buf[2] ),
    .D(\SLICE[0].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[6].W.SEL1 ));
 sky130_fd_sc_hd__and4_2 \SLICE[0].RAM8.DEC1.AND7  (.A(\SLICE[0].RAM8.DEC1.A_buf[0] ),
    .B(\SLICE[0].RAM8.DEC1.A_buf[1] ),
    .C(\SLICE[0].RAM8.DEC1.A_buf[2] ),
    .D(\SLICE[0].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[7].W.SEL1 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.DEC1.ENBUF  (.A(\SLICE[0].RAM8.DEC1.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.DEC1.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.WEBUF[0].__cell__  (.A(\SLICE[0].RAM8.WEBUF[0].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WEBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.WEBUF[1].__cell__  (.A(\SLICE[0].RAM8.WEBUF[1].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WEBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.WEBUF[2].__cell__  (.A(\SLICE[0].RAM8.WEBUF[2].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WEBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.WEBUF[3].__cell__  (.A(\SLICE[0].RAM8.WEBUF[3].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WEBUF[3].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.WEBUF[4].__cell__  (.A(\SLICE[0].RAM8.WEBUF[4].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WEBUF[4].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.WEBUF[5].__cell__  (.A(\SLICE[0].RAM8.WEBUF[5].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WEBUF[5].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.WEBUF[6].__cell__  (.A(\SLICE[0].RAM8.WEBUF[6].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WEBUF[6].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.WEBUF[7].__cell__  (.A(\SLICE[0].RAM8.WEBUF[7].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WEBUF[7].X ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.CGAND  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[0].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[0].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.CGAND  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[0].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[0].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.CGAND  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[0].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[0].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.CGAND  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[0].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[0].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[0].RAM8.WORD[0].W.CLKBUF  (.A(\SLICE[0].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.WORD[0].W.SEL0BUF  (.A(\SLICE[0].RAM8.WORD[0].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.WORD[0].W.SEL1BUF  (.A(\SLICE[0].RAM8.WORD[0].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.CGAND  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[1].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[1].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.CGAND  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[1].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[1].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.CGAND  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[1].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[1].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.CGAND  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[1].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[1].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[0].RAM8.WORD[1].W.CLKBUF  (.A(\SLICE[0].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.WORD[1].W.SEL0BUF  (.A(\SLICE[0].RAM8.WORD[1].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.WORD[1].W.SEL1BUF  (.A(\SLICE[0].RAM8.WORD[1].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.CGAND  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[2].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[2].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.CGAND  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[2].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[2].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.CGAND  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[2].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[2].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.CGAND  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[2].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[2].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[0].RAM8.WORD[2].W.CLKBUF  (.A(\SLICE[0].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.WORD[2].W.SEL0BUF  (.A(\SLICE[0].RAM8.WORD[2].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.WORD[2].W.SEL1BUF  (.A(\SLICE[0].RAM8.WORD[2].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.CGAND  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[3].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[3].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.CGAND  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[3].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[3].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.CGAND  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[3].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[3].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.CGAND  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[3].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[3].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[0].RAM8.WORD[3].W.CLKBUF  (.A(\SLICE[0].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.WORD[3].W.SEL0BUF  (.A(\SLICE[0].RAM8.WORD[3].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.WORD[3].W.SEL1BUF  (.A(\SLICE[0].RAM8.WORD[3].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.CGAND  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[4].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[4].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.CGAND  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[4].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[4].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.CGAND  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[4].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[4].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.CGAND  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[4].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[4].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[0].RAM8.WORD[4].W.CLKBUF  (.A(\SLICE[0].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.WORD[4].W.SEL0BUF  (.A(\SLICE[0].RAM8.WORD[4].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.WORD[4].W.SEL1BUF  (.A(\SLICE[0].RAM8.WORD[4].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.CGAND  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[5].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[5].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.CGAND  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[5].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[5].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.CGAND  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[5].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[5].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.CGAND  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[5].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[5].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[0].RAM8.WORD[5].W.CLKBUF  (.A(\SLICE[0].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.WORD[5].W.SEL0BUF  (.A(\SLICE[0].RAM8.WORD[5].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.WORD[5].W.SEL1BUF  (.A(\SLICE[0].RAM8.WORD[5].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.CGAND  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[6].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[6].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.CGAND  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[6].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[6].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.CGAND  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[6].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[6].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.CGAND  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[6].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[6].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[0].RAM8.WORD[6].W.CLKBUF  (.A(\SLICE[0].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.WORD[6].W.SEL0BUF  (.A(\SLICE[0].RAM8.WORD[6].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.WORD[6].W.SEL1BUF  (.A(\SLICE[0].RAM8.WORD[6].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.CGAND  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[7].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[7].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.CGAND  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[7].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[7].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.CGAND  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[7].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[7].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.CGAND  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[0].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.SEL0INV  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.SEL1INV  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[0].RAM8.WORD[7].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[0].RAM8.WORD[7].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[0].RAM8.WORD[7].W.CLKBUF  (.A(\SLICE[0].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.WORD[7].W.SEL0BUF  (.A(\SLICE[0].RAM8.WORD[7].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[0].RAM8.WORD[7].W.SEL1BUF  (.A(\SLICE[0].RAM8.WORD[7].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.CLKBUF.__cell__  (.A(\CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.DEC0.ABUF[0]  (.A(\A0BUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.DEC0.ABUF[1]  (.A(\A0BUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.DEC0.ABUF[2]  (.A(\A0BUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \SLICE[1].RAM8.DEC0.AND0  (.A(\SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D_N(\SLICE[1].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE[1].RAM8.DEC0.AND1  (.A_N(\SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\SLICE[1].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE[1].RAM8.DEC0.AND2  (.A_N(\SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\SLICE[1].RAM8.DEC0.A_buf[1] ),
    .D(\SLICE[1].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \SLICE[1].RAM8.DEC0.AND3  (.A_N(\SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B(\SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\SLICE[1].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE[1].RAM8.DEC0.AND4  (.A_N(\SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B_N(\SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE[1].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \SLICE[1].RAM8.DEC0.AND5  (.A_N(\SLICE[1].RAM8.DEC0.A_buf[1] ),
    .B(\SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE[1].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \SLICE[1].RAM8.DEC0.AND6  (.A_N(\SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE[1].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \SLICE[1].RAM8.DEC0.AND7  (.A(\SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE[1].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.DEC0.ENBUF  (.A(\SLICE[1].RAM8.DEC0.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.DEC1.ABUF[0]  (.A(\A1BUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.DEC1.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.DEC1.ABUF[1]  (.A(\A1BUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.DEC1.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.DEC1.ABUF[2]  (.A(\A1BUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.DEC1.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \SLICE[1].RAM8.DEC1.AND0  (.A(\SLICE[1].RAM8.DEC1.A_buf[0] ),
    .B(\SLICE[1].RAM8.DEC1.A_buf[1] ),
    .C(\SLICE[1].RAM8.DEC1.A_buf[2] ),
    .D_N(\SLICE[1].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[0].W.SEL1 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE[1].RAM8.DEC1.AND1  (.A_N(\SLICE[1].RAM8.DEC1.A_buf[2] ),
    .B_N(\SLICE[1].RAM8.DEC1.A_buf[1] ),
    .C(\SLICE[1].RAM8.DEC1.A_buf[0] ),
    .D(\SLICE[1].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[1].W.SEL1 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE[1].RAM8.DEC1.AND2  (.A_N(\SLICE[1].RAM8.DEC1.A_buf[2] ),
    .B_N(\SLICE[1].RAM8.DEC1.A_buf[0] ),
    .C(\SLICE[1].RAM8.DEC1.A_buf[1] ),
    .D(\SLICE[1].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[2].W.SEL1 ));
 sky130_fd_sc_hd__and4b_2 \SLICE[1].RAM8.DEC1.AND3  (.A_N(\SLICE[1].RAM8.DEC1.A_buf[2] ),
    .B(\SLICE[1].RAM8.DEC1.A_buf[1] ),
    .C(\SLICE[1].RAM8.DEC1.A_buf[0] ),
    .D(\SLICE[1].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[3].W.SEL1 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE[1].RAM8.DEC1.AND4  (.A_N(\SLICE[1].RAM8.DEC1.A_buf[0] ),
    .B_N(\SLICE[1].RAM8.DEC1.A_buf[1] ),
    .C(\SLICE[1].RAM8.DEC1.A_buf[2] ),
    .D(\SLICE[1].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[4].W.SEL1 ));
 sky130_fd_sc_hd__and4b_2 \SLICE[1].RAM8.DEC1.AND5  (.A_N(\SLICE[1].RAM8.DEC1.A_buf[1] ),
    .B(\SLICE[1].RAM8.DEC1.A_buf[0] ),
    .C(\SLICE[1].RAM8.DEC1.A_buf[2] ),
    .D(\SLICE[1].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[5].W.SEL1 ));
 sky130_fd_sc_hd__and4b_2 \SLICE[1].RAM8.DEC1.AND6  (.A_N(\SLICE[1].RAM8.DEC1.A_buf[0] ),
    .B(\SLICE[1].RAM8.DEC1.A_buf[1] ),
    .C(\SLICE[1].RAM8.DEC1.A_buf[2] ),
    .D(\SLICE[1].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[6].W.SEL1 ));
 sky130_fd_sc_hd__and4_2 \SLICE[1].RAM8.DEC1.AND7  (.A(\SLICE[1].RAM8.DEC1.A_buf[0] ),
    .B(\SLICE[1].RAM8.DEC1.A_buf[1] ),
    .C(\SLICE[1].RAM8.DEC1.A_buf[2] ),
    .D(\SLICE[1].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[7].W.SEL1 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.DEC1.ENBUF  (.A(\SLICE[1].RAM8.DEC1.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.DEC1.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.WEBUF[0].__cell__  (.A(\SLICE[0].RAM8.WEBUF[0].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WEBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.WEBUF[1].__cell__  (.A(\SLICE[0].RAM8.WEBUF[1].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WEBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.WEBUF[2].__cell__  (.A(\SLICE[0].RAM8.WEBUF[2].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WEBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.WEBUF[3].__cell__  (.A(\SLICE[0].RAM8.WEBUF[3].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WEBUF[3].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.WEBUF[4].__cell__  (.A(\SLICE[0].RAM8.WEBUF[4].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WEBUF[4].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.WEBUF[5].__cell__  (.A(\SLICE[0].RAM8.WEBUF[5].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WEBUF[5].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.WEBUF[6].__cell__  (.A(\SLICE[0].RAM8.WEBUF[6].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WEBUF[6].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.WEBUF[7].__cell__  (.A(\SLICE[0].RAM8.WEBUF[7].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WEBUF[7].X ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.CGAND  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[0].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[0].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.CGAND  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[0].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[0].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.CGAND  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[0].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[0].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.CGAND  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[0].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[0].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[1].RAM8.WORD[0].W.CLKBUF  (.A(\SLICE[1].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.WORD[0].W.SEL0BUF  (.A(\SLICE[1].RAM8.WORD[0].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.WORD[0].W.SEL1BUF  (.A(\SLICE[1].RAM8.WORD[0].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.CGAND  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[1].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[1].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.CGAND  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[1].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[1].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.CGAND  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[1].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[1].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.CGAND  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[1].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[1].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[1].RAM8.WORD[1].W.CLKBUF  (.A(\SLICE[1].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.WORD[1].W.SEL0BUF  (.A(\SLICE[1].RAM8.WORD[1].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.WORD[1].W.SEL1BUF  (.A(\SLICE[1].RAM8.WORD[1].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.CGAND  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[2].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[2].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.CGAND  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[2].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[2].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.CGAND  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[2].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[2].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.CGAND  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[2].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[2].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[1].RAM8.WORD[2].W.CLKBUF  (.A(\SLICE[1].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.WORD[2].W.SEL0BUF  (.A(\SLICE[1].RAM8.WORD[2].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.WORD[2].W.SEL1BUF  (.A(\SLICE[1].RAM8.WORD[2].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.CGAND  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[3].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[3].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.CGAND  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[3].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[3].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.CGAND  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[3].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[3].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.CGAND  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[3].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[3].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[1].RAM8.WORD[3].W.CLKBUF  (.A(\SLICE[1].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.WORD[3].W.SEL0BUF  (.A(\SLICE[1].RAM8.WORD[3].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.WORD[3].W.SEL1BUF  (.A(\SLICE[1].RAM8.WORD[3].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.CGAND  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[4].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[4].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.CGAND  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[4].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[4].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.CGAND  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[4].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[4].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.CGAND  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[4].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[4].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[1].RAM8.WORD[4].W.CLKBUF  (.A(\SLICE[1].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.WORD[4].W.SEL0BUF  (.A(\SLICE[1].RAM8.WORD[4].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.WORD[4].W.SEL1BUF  (.A(\SLICE[1].RAM8.WORD[4].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.CGAND  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[5].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[5].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.CGAND  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[5].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[5].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.CGAND  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[5].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[5].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.CGAND  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[5].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[5].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[1].RAM8.WORD[5].W.CLKBUF  (.A(\SLICE[1].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.WORD[5].W.SEL0BUF  (.A(\SLICE[1].RAM8.WORD[5].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.WORD[5].W.SEL1BUF  (.A(\SLICE[1].RAM8.WORD[5].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.CGAND  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[6].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[6].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.CGAND  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[6].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[6].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.CGAND  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[6].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[6].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.CGAND  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[6].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[6].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[1].RAM8.WORD[6].W.CLKBUF  (.A(\SLICE[1].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.WORD[6].W.SEL0BUF  (.A(\SLICE[1].RAM8.WORD[6].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.WORD[6].W.SEL1BUF  (.A(\SLICE[1].RAM8.WORD[6].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.CGAND  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[7].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[7].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.CGAND  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[7].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[7].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.CGAND  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[7].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[7].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.CGAND  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[1].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.SEL0INV  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.SEL1INV  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[1].RAM8.WORD[7].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[1].RAM8.WORD[7].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[1].RAM8.WORD[7].W.CLKBUF  (.A(\SLICE[1].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.WORD[7].W.SEL0BUF  (.A(\SLICE[1].RAM8.WORD[7].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[1].RAM8.WORD[7].W.SEL1BUF  (.A(\SLICE[1].RAM8.WORD[7].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.CLKBUF.__cell__  (.A(\CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.DEC0.ABUF[0]  (.A(\A0BUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.DEC0.ABUF[1]  (.A(\A0BUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.DEC0.ABUF[2]  (.A(\A0BUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \SLICE[2].RAM8.DEC0.AND0  (.A(\SLICE[2].RAM8.DEC0.A_buf[0] ),
    .B(\SLICE[2].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE[2].RAM8.DEC0.A_buf[2] ),
    .D_N(\SLICE[2].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE[2].RAM8.DEC0.AND1  (.A_N(\SLICE[2].RAM8.DEC0.A_buf[2] ),
    .B_N(\SLICE[2].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE[2].RAM8.DEC0.A_buf[0] ),
    .D(\SLICE[2].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE[2].RAM8.DEC0.AND2  (.A_N(\SLICE[2].RAM8.DEC0.A_buf[2] ),
    .B_N(\SLICE[2].RAM8.DEC0.A_buf[0] ),
    .C(\SLICE[2].RAM8.DEC0.A_buf[1] ),
    .D(\SLICE[2].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \SLICE[2].RAM8.DEC0.AND3  (.A_N(\SLICE[2].RAM8.DEC0.A_buf[2] ),
    .B(\SLICE[2].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE[2].RAM8.DEC0.A_buf[0] ),
    .D(\SLICE[2].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE[2].RAM8.DEC0.AND4  (.A_N(\SLICE[2].RAM8.DEC0.A_buf[0] ),
    .B_N(\SLICE[2].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE[2].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE[2].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \SLICE[2].RAM8.DEC0.AND5  (.A_N(\SLICE[2].RAM8.DEC0.A_buf[1] ),
    .B(\SLICE[2].RAM8.DEC0.A_buf[0] ),
    .C(\SLICE[2].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE[2].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \SLICE[2].RAM8.DEC0.AND6  (.A_N(\SLICE[2].RAM8.DEC0.A_buf[0] ),
    .B(\SLICE[2].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE[2].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE[2].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \SLICE[2].RAM8.DEC0.AND7  (.A(\SLICE[2].RAM8.DEC0.A_buf[0] ),
    .B(\SLICE[2].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE[2].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE[2].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.DEC0.ENBUF  (.A(\SLICE[2].RAM8.DEC0.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.DEC1.ABUF[0]  (.A(\A1BUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.DEC1.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.DEC1.ABUF[1]  (.A(\A1BUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.DEC1.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.DEC1.ABUF[2]  (.A(\A1BUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.DEC1.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \SLICE[2].RAM8.DEC1.AND0  (.A(\SLICE[2].RAM8.DEC1.A_buf[0] ),
    .B(\SLICE[2].RAM8.DEC1.A_buf[1] ),
    .C(\SLICE[2].RAM8.DEC1.A_buf[2] ),
    .D_N(\SLICE[2].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[0].W.SEL1 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE[2].RAM8.DEC1.AND1  (.A_N(\SLICE[2].RAM8.DEC1.A_buf[2] ),
    .B_N(\SLICE[2].RAM8.DEC1.A_buf[1] ),
    .C(\SLICE[2].RAM8.DEC1.A_buf[0] ),
    .D(\SLICE[2].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[1].W.SEL1 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE[2].RAM8.DEC1.AND2  (.A_N(\SLICE[2].RAM8.DEC1.A_buf[2] ),
    .B_N(\SLICE[2].RAM8.DEC1.A_buf[0] ),
    .C(\SLICE[2].RAM8.DEC1.A_buf[1] ),
    .D(\SLICE[2].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[2].W.SEL1 ));
 sky130_fd_sc_hd__and4b_2 \SLICE[2].RAM8.DEC1.AND3  (.A_N(\SLICE[2].RAM8.DEC1.A_buf[2] ),
    .B(\SLICE[2].RAM8.DEC1.A_buf[1] ),
    .C(\SLICE[2].RAM8.DEC1.A_buf[0] ),
    .D(\SLICE[2].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[3].W.SEL1 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE[2].RAM8.DEC1.AND4  (.A_N(\SLICE[2].RAM8.DEC1.A_buf[0] ),
    .B_N(\SLICE[2].RAM8.DEC1.A_buf[1] ),
    .C(\SLICE[2].RAM8.DEC1.A_buf[2] ),
    .D(\SLICE[2].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[4].W.SEL1 ));
 sky130_fd_sc_hd__and4b_2 \SLICE[2].RAM8.DEC1.AND5  (.A_N(\SLICE[2].RAM8.DEC1.A_buf[1] ),
    .B(\SLICE[2].RAM8.DEC1.A_buf[0] ),
    .C(\SLICE[2].RAM8.DEC1.A_buf[2] ),
    .D(\SLICE[2].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[5].W.SEL1 ));
 sky130_fd_sc_hd__and4b_2 \SLICE[2].RAM8.DEC1.AND6  (.A_N(\SLICE[2].RAM8.DEC1.A_buf[0] ),
    .B(\SLICE[2].RAM8.DEC1.A_buf[1] ),
    .C(\SLICE[2].RAM8.DEC1.A_buf[2] ),
    .D(\SLICE[2].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[6].W.SEL1 ));
 sky130_fd_sc_hd__and4_2 \SLICE[2].RAM8.DEC1.AND7  (.A(\SLICE[2].RAM8.DEC1.A_buf[0] ),
    .B(\SLICE[2].RAM8.DEC1.A_buf[1] ),
    .C(\SLICE[2].RAM8.DEC1.A_buf[2] ),
    .D(\SLICE[2].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[7].W.SEL1 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.DEC1.ENBUF  (.A(\SLICE[2].RAM8.DEC1.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.DEC1.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.WEBUF[0].__cell__  (.A(\SLICE[0].RAM8.WEBUF[0].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WEBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.WEBUF[1].__cell__  (.A(\SLICE[0].RAM8.WEBUF[1].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WEBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.WEBUF[2].__cell__  (.A(\SLICE[0].RAM8.WEBUF[2].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WEBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.WEBUF[3].__cell__  (.A(\SLICE[0].RAM8.WEBUF[3].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WEBUF[3].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.WEBUF[4].__cell__  (.A(\SLICE[0].RAM8.WEBUF[4].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WEBUF[4].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.WEBUF[5].__cell__  (.A(\SLICE[0].RAM8.WEBUF[5].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WEBUF[5].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.WEBUF[6].__cell__  (.A(\SLICE[0].RAM8.WEBUF[6].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WEBUF[6].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.WEBUF[7].__cell__  (.A(\SLICE[0].RAM8.WEBUF[7].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WEBUF[7].X ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.CGAND  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[0].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[0].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.CGAND  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[0].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[0].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.CGAND  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[0].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[0].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.CGAND  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[0].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[0].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[2].RAM8.WORD[0].W.CLKBUF  (.A(\SLICE[2].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.WORD[0].W.SEL0BUF  (.A(\SLICE[2].RAM8.WORD[0].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.WORD[0].W.SEL1BUF  (.A(\SLICE[2].RAM8.WORD[0].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.CGAND  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[1].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[1].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.CGAND  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[1].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[1].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.CGAND  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[1].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[1].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.CGAND  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[1].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[1].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[2].RAM8.WORD[1].W.CLKBUF  (.A(\SLICE[2].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.WORD[1].W.SEL0BUF  (.A(\SLICE[2].RAM8.WORD[1].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.WORD[1].W.SEL1BUF  (.A(\SLICE[2].RAM8.WORD[1].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.CGAND  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[2].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[2].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.CGAND  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[2].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[2].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.CGAND  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[2].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[2].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.CGAND  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[2].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[2].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[2].RAM8.WORD[2].W.CLKBUF  (.A(\SLICE[2].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.WORD[2].W.SEL0BUF  (.A(\SLICE[2].RAM8.WORD[2].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.WORD[2].W.SEL1BUF  (.A(\SLICE[2].RAM8.WORD[2].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.CGAND  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[3].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[3].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.CGAND  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[3].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[3].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.CGAND  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[3].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[3].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.CGAND  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[3].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[3].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[2].RAM8.WORD[3].W.CLKBUF  (.A(\SLICE[2].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.WORD[3].W.SEL0BUF  (.A(\SLICE[2].RAM8.WORD[3].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.WORD[3].W.SEL1BUF  (.A(\SLICE[2].RAM8.WORD[3].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.CGAND  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[4].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[4].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.CGAND  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[4].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[4].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.CGAND  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[4].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[4].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.CGAND  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[4].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[4].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[2].RAM8.WORD[4].W.CLKBUF  (.A(\SLICE[2].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.WORD[4].W.SEL0BUF  (.A(\SLICE[2].RAM8.WORD[4].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.WORD[4].W.SEL1BUF  (.A(\SLICE[2].RAM8.WORD[4].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.CGAND  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[5].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[5].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.CGAND  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[5].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[5].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.CGAND  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[5].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[5].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.CGAND  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[5].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[5].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[2].RAM8.WORD[5].W.CLKBUF  (.A(\SLICE[2].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.WORD[5].W.SEL0BUF  (.A(\SLICE[2].RAM8.WORD[5].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.WORD[5].W.SEL1BUF  (.A(\SLICE[2].RAM8.WORD[5].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.CGAND  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[6].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[6].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.CGAND  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[6].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[6].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.CGAND  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[6].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[6].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.CGAND  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[6].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[6].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[2].RAM8.WORD[6].W.CLKBUF  (.A(\SLICE[2].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.WORD[6].W.SEL0BUF  (.A(\SLICE[2].RAM8.WORD[6].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.WORD[6].W.SEL1BUF  (.A(\SLICE[2].RAM8.WORD[6].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.CGAND  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[7].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[7].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.CGAND  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[7].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[7].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.CGAND  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[7].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[7].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.CGAND  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[2].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.SEL0INV  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.SEL1INV  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[2].RAM8.WORD[7].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[2].RAM8.WORD[7].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[2].RAM8.WORD[7].W.CLKBUF  (.A(\SLICE[2].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.WORD[7].W.SEL0BUF  (.A(\SLICE[2].RAM8.WORD[7].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[2].RAM8.WORD[7].W.SEL1BUF  (.A(\SLICE[2].RAM8.WORD[7].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.CLKBUF.__cell__  (.A(\CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.DEC0.ABUF[0]  (.A(\A0BUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.DEC0.ABUF[1]  (.A(\A0BUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.DEC0.ABUF[2]  (.A(\A0BUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \SLICE[3].RAM8.DEC0.AND0  (.A(\SLICE[3].RAM8.DEC0.A_buf[0] ),
    .B(\SLICE[3].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE[3].RAM8.DEC0.A_buf[2] ),
    .D_N(\SLICE[3].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE[3].RAM8.DEC0.AND1  (.A_N(\SLICE[3].RAM8.DEC0.A_buf[2] ),
    .B_N(\SLICE[3].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE[3].RAM8.DEC0.A_buf[0] ),
    .D(\SLICE[3].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE[3].RAM8.DEC0.AND2  (.A_N(\SLICE[3].RAM8.DEC0.A_buf[2] ),
    .B_N(\SLICE[3].RAM8.DEC0.A_buf[0] ),
    .C(\SLICE[3].RAM8.DEC0.A_buf[1] ),
    .D(\SLICE[3].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \SLICE[3].RAM8.DEC0.AND3  (.A_N(\SLICE[3].RAM8.DEC0.A_buf[2] ),
    .B(\SLICE[3].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE[3].RAM8.DEC0.A_buf[0] ),
    .D(\SLICE[3].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE[3].RAM8.DEC0.AND4  (.A_N(\SLICE[3].RAM8.DEC0.A_buf[0] ),
    .B_N(\SLICE[3].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE[3].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE[3].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \SLICE[3].RAM8.DEC0.AND5  (.A_N(\SLICE[3].RAM8.DEC0.A_buf[1] ),
    .B(\SLICE[3].RAM8.DEC0.A_buf[0] ),
    .C(\SLICE[3].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE[3].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \SLICE[3].RAM8.DEC0.AND6  (.A_N(\SLICE[3].RAM8.DEC0.A_buf[0] ),
    .B(\SLICE[3].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE[3].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE[3].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \SLICE[3].RAM8.DEC0.AND7  (.A(\SLICE[3].RAM8.DEC0.A_buf[0] ),
    .B(\SLICE[3].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE[3].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE[3].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.DEC0.ENBUF  (.A(\SLICE[3].RAM8.DEC0.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.DEC1.ABUF[0]  (.A(\A1BUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.DEC1.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.DEC1.ABUF[1]  (.A(\A1BUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.DEC1.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.DEC1.ABUF[2]  (.A(\A1BUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.DEC1.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \SLICE[3].RAM8.DEC1.AND0  (.A(\SLICE[3].RAM8.DEC1.A_buf[0] ),
    .B(\SLICE[3].RAM8.DEC1.A_buf[1] ),
    .C(\SLICE[3].RAM8.DEC1.A_buf[2] ),
    .D_N(\SLICE[3].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[0].W.SEL1 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE[3].RAM8.DEC1.AND1  (.A_N(\SLICE[3].RAM8.DEC1.A_buf[2] ),
    .B_N(\SLICE[3].RAM8.DEC1.A_buf[1] ),
    .C(\SLICE[3].RAM8.DEC1.A_buf[0] ),
    .D(\SLICE[3].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[1].W.SEL1 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE[3].RAM8.DEC1.AND2  (.A_N(\SLICE[3].RAM8.DEC1.A_buf[2] ),
    .B_N(\SLICE[3].RAM8.DEC1.A_buf[0] ),
    .C(\SLICE[3].RAM8.DEC1.A_buf[1] ),
    .D(\SLICE[3].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[2].W.SEL1 ));
 sky130_fd_sc_hd__and4b_2 \SLICE[3].RAM8.DEC1.AND3  (.A_N(\SLICE[3].RAM8.DEC1.A_buf[2] ),
    .B(\SLICE[3].RAM8.DEC1.A_buf[1] ),
    .C(\SLICE[3].RAM8.DEC1.A_buf[0] ),
    .D(\SLICE[3].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[3].W.SEL1 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE[3].RAM8.DEC1.AND4  (.A_N(\SLICE[3].RAM8.DEC1.A_buf[0] ),
    .B_N(\SLICE[3].RAM8.DEC1.A_buf[1] ),
    .C(\SLICE[3].RAM8.DEC1.A_buf[2] ),
    .D(\SLICE[3].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[4].W.SEL1 ));
 sky130_fd_sc_hd__and4b_2 \SLICE[3].RAM8.DEC1.AND5  (.A_N(\SLICE[3].RAM8.DEC1.A_buf[1] ),
    .B(\SLICE[3].RAM8.DEC1.A_buf[0] ),
    .C(\SLICE[3].RAM8.DEC1.A_buf[2] ),
    .D(\SLICE[3].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[5].W.SEL1 ));
 sky130_fd_sc_hd__and4b_2 \SLICE[3].RAM8.DEC1.AND6  (.A_N(\SLICE[3].RAM8.DEC1.A_buf[0] ),
    .B(\SLICE[3].RAM8.DEC1.A_buf[1] ),
    .C(\SLICE[3].RAM8.DEC1.A_buf[2] ),
    .D(\SLICE[3].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[6].W.SEL1 ));
 sky130_fd_sc_hd__and4_2 \SLICE[3].RAM8.DEC1.AND7  (.A(\SLICE[3].RAM8.DEC1.A_buf[0] ),
    .B(\SLICE[3].RAM8.DEC1.A_buf[1] ),
    .C(\SLICE[3].RAM8.DEC1.A_buf[2] ),
    .D(\SLICE[3].RAM8.DEC1.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[7].W.SEL1 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.DEC1.ENBUF  (.A(\SLICE[3].RAM8.DEC1.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.DEC1.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.WEBUF[0].__cell__  (.A(\SLICE[0].RAM8.WEBUF[0].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WEBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.WEBUF[1].__cell__  (.A(\SLICE[0].RAM8.WEBUF[1].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WEBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.WEBUF[2].__cell__  (.A(\SLICE[0].RAM8.WEBUF[2].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WEBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.WEBUF[3].__cell__  (.A(\SLICE[0].RAM8.WEBUF[3].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WEBUF[3].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.WEBUF[4].__cell__  (.A(\SLICE[0].RAM8.WEBUF[4].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WEBUF[4].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.WEBUF[5].__cell__  (.A(\SLICE[0].RAM8.WEBUF[5].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WEBUF[5].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.WEBUF[6].__cell__  (.A(\SLICE[0].RAM8.WEBUF[6].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WEBUF[6].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.WEBUF[7].__cell__  (.A(\SLICE[0].RAM8.WEBUF[7].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WEBUF[7].X ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.CGAND  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[0].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[0].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.CGAND  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[0].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[0].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.CGAND  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[0].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[0].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.CGAND  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[0].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[0].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[3].RAM8.WORD[0].W.CLKBUF  (.A(\SLICE[3].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.WORD[0].W.SEL0BUF  (.A(\SLICE[3].RAM8.WORD[0].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.WORD[0].W.SEL1BUF  (.A(\SLICE[3].RAM8.WORD[0].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.CGAND  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[1].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[1].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.CGAND  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[1].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[1].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.CGAND  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[1].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[1].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.CGAND  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[1].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[1].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[3].RAM8.WORD[1].W.CLKBUF  (.A(\SLICE[3].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.WORD[1].W.SEL0BUF  (.A(\SLICE[3].RAM8.WORD[1].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.WORD[1].W.SEL1BUF  (.A(\SLICE[3].RAM8.WORD[1].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.CGAND  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[2].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[2].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.CGAND  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[2].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[2].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.CGAND  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[2].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[2].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.CGAND  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[2].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[2].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[3].RAM8.WORD[2].W.CLKBUF  (.A(\SLICE[3].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.WORD[2].W.SEL0BUF  (.A(\SLICE[3].RAM8.WORD[2].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.WORD[2].W.SEL1BUF  (.A(\SLICE[3].RAM8.WORD[2].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.CGAND  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[3].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[3].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.CGAND  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[3].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[3].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.CGAND  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[3].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[3].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.CGAND  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[3].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[3].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[3].RAM8.WORD[3].W.CLKBUF  (.A(\SLICE[3].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.WORD[3].W.SEL0BUF  (.A(\SLICE[3].RAM8.WORD[3].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.WORD[3].W.SEL1BUF  (.A(\SLICE[3].RAM8.WORD[3].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.CGAND  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[4].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[4].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.CGAND  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[4].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[4].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.CGAND  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[4].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[4].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.CGAND  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[4].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[4].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[3].RAM8.WORD[4].W.CLKBUF  (.A(\SLICE[3].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.WORD[4].W.SEL0BUF  (.A(\SLICE[3].RAM8.WORD[4].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.WORD[4].W.SEL1BUF  (.A(\SLICE[3].RAM8.WORD[4].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.CGAND  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[5].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[5].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.CGAND  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[5].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[5].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.CGAND  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[5].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[5].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.CGAND  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[5].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[5].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[3].RAM8.WORD[5].W.CLKBUF  (.A(\SLICE[3].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.WORD[5].W.SEL0BUF  (.A(\SLICE[3].RAM8.WORD[5].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.WORD[5].W.SEL1BUF  (.A(\SLICE[3].RAM8.WORD[5].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.CGAND  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[6].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[6].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.CGAND  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[6].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[6].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.CGAND  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[6].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[6].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.CGAND  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[6].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[6].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[3].RAM8.WORD[6].W.CLKBUF  (.A(\SLICE[3].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.WORD[6].W.SEL0BUF  (.A(\SLICE[3].RAM8.WORD[6].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.WORD[6].W.SEL1BUF  (.A(\SLICE[3].RAM8.WORD[6].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[32].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[32].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[32].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[33].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[33].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[33].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[34].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[34].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[34].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[35].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[35].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[35].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[36].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[36].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[36].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[37].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[37].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[37].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[38].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[38].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[38].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF0[39].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[4].FLOATBUF1[39].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[39].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.CGAND  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[7].W.BYTE[4].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[7].W.BYTE[4].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[40].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[40].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[40].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[41].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[41].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[41].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[42].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[42].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[42].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[43].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[43].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[43].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[44].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[44].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[44].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[45].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[45].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[45].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[46].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[46].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[46].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF0[47].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[5].FLOATBUF1[47].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[47].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.CGAND  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[5].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[7].W.BYTE[5].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[7].W.BYTE[5].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[48].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[48].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[48].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[49].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[49].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[49].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[50].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[50].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[50].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[51].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[51].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[51].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[52].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[52].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[52].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[53].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[53].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[53].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[54].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[54].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[54].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF0[55].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[6].FLOATBUF1[55].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[55].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.CGAND  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[6].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[7].W.BYTE[6].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[7].W.BYTE[6].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.BIT[0].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[56].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.BIT[0].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[0] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[56].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[56].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.BIT[1].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[57].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.BIT[1].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[1] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[57].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[57].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.BIT[2].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[58].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.BIT[2].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[2] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[58].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[58].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.BIT[3].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[59].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.BIT[3].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[3] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[59].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[59].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.BIT[4].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[60].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.BIT[4].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[4] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[60].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[60].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.BIT[5].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[61].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.BIT[5].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[5] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[61].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[61].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.BIT[6].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[62].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.BIT[6].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[6] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[62].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[62].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.BIT[7].OBUF0  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF0[63].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.BIT[7].OBUF1  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[7] ),
    .TE_B(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\BYTE[7].FLOATBUF1[63].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[63].X ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.CGAND  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE[3].RAM8.WEBUF[7].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.DIODE_CLK  (.DIODE(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.SEL0INV  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.SEL0_B ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.SEL1INV  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.SEL1_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.CLK_B ),
    .GATE(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE[3].RAM8.WORD[7].W.BYTE[7].B.genblk1.CLKINV  (.A(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE[3].RAM8.WORD[7].W.BYTE[7].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE[3].RAM8.WORD[7].W.CLKBUF  (.A(\SLICE[3].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.WORD[7].W.SEL0BUF  (.A(\SLICE[3].RAM8.WORD[7].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE[3].RAM8.WORD[7].W.SEL1BUF  (.A(\SLICE[3].RAM8.WORD[7].W.SEL1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1 ));
 sky130_fd_sc_hd__conb_1 \TIE0[0].__cell__  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(\BYTE[0].FLOATBUF0[0].A ));
 sky130_fd_sc_hd__conb_1 \TIE0[1].__cell__  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(\BYTE[1].FLOATBUF0[10].A ));
 sky130_fd_sc_hd__conb_1 \TIE0[2].__cell__  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(\BYTE[2].FLOATBUF0[16].A ));
 sky130_fd_sc_hd__conb_1 \TIE0[3].__cell__  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(\BYTE[3].FLOATBUF0[24].A ));
 sky130_fd_sc_hd__conb_1 \TIE0[4].__cell__  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(\BYTE[4].FLOATBUF0[32].A ));
 sky130_fd_sc_hd__conb_1 \TIE0[5].__cell__  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(\BYTE[5].FLOATBUF0[40].A ));
 sky130_fd_sc_hd__conb_1 \TIE0[6].__cell__  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(\BYTE[6].FLOATBUF0[48].A ));
 sky130_fd_sc_hd__conb_1 \TIE0[7].__cell__  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(\BYTE[7].FLOATBUF0[56].A ));
 sky130_fd_sc_hd__conb_1 \TIE1[0].__cell__  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(\BYTE[0].FLOATBUF1[0].A ));
 sky130_fd_sc_hd__conb_1 \TIE1[1].__cell__  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(\BYTE[1].FLOATBUF1[10].A ));
 sky130_fd_sc_hd__conb_1 \TIE1[2].__cell__  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(\BYTE[2].FLOATBUF1[16].A ));
 sky130_fd_sc_hd__conb_1 \TIE1[3].__cell__  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(\BYTE[3].FLOATBUF1[24].A ));
 sky130_fd_sc_hd__conb_1 \TIE1[4].__cell__  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(\BYTE[4].FLOATBUF1[32].A ));
 sky130_fd_sc_hd__conb_1 \TIE1[5].__cell__  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(\BYTE[5].FLOATBUF1[40].A ));
 sky130_fd_sc_hd__conb_1 \TIE1[6].__cell__  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(\BYTE[6].FLOATBUF1[48].A ));
 sky130_fd_sc_hd__conb_1 \TIE1[7].__cell__  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(\BYTE[7].FLOATBUF1[56].A ));
 sky130_fd_sc_hd__clkbuf_2 \WEBUF[0].__cell__  (.A(WE0[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WEBUF[0].A ));
 sky130_fd_sc_hd__clkbuf_2 \WEBUF[1].__cell__  (.A(WE0[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WEBUF[1].A ));
 sky130_fd_sc_hd__clkbuf_2 \WEBUF[2].__cell__  (.A(WE0[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WEBUF[2].A ));
 sky130_fd_sc_hd__clkbuf_2 \WEBUF[3].__cell__  (.A(WE0[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WEBUF[3].A ));
 sky130_fd_sc_hd__clkbuf_2 \WEBUF[4].__cell__  (.A(WE0[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WEBUF[4].A ));
 sky130_fd_sc_hd__clkbuf_2 \WEBUF[5].__cell__  (.A(WE0[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WEBUF[5].A ));
 sky130_fd_sc_hd__clkbuf_2 \WEBUF[6].__cell__  (.A(WE0[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WEBUF[6].A ));
 sky130_fd_sc_hd__clkbuf_2 \WEBUF[7].__cell__  (.A(WE0[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE[0].RAM8.WEBUF[7].A ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_0_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_1_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_1_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_2_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_2_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_2_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_3_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_3_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_4_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_4_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_4_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_5_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_5_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_7_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_8_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_8_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_9_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_9_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_10_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_10_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_10_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_11_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_11_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_12_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_12_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_12_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_13_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_13_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_14_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_14_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_14_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_15_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_15_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_16_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_16_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_16_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_17_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_72 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_72 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_72 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_72 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_2_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_2_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_3_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_3_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_4_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_4_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_5_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_5_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_5_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_6_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_6_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_7_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_7_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_8_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_8_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_8_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_73 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_2_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_2_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_3_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_3_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_4_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_4_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_5_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_5_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_6_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_6_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_7_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_7_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_8_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_8_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_72 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_72 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_72 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_72 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_10_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_10_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_11_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_11_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_12_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_12_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_13_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_13_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_13_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_14_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_14_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_15_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_15_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_16_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_16_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_16_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_73 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_10_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_10_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_11_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_11_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_12_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_12_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_13_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_13_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_14_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_14_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_15_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_15_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_16_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_16_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_72 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_72 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_72 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_72 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_18_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 fill_18_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 fill_18_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_19_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 fill_19_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_19_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_20_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_20_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_21_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_21_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_21_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_22_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_22_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_22_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_23_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_23_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 fill_23_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_24_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_24_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_24_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_24_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_73 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_18_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_18_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_19_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_19_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_20_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_20_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_21_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_21_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_22_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_22_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_23_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_23_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_24_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_24_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_72 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_72 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_72 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_72 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_26_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_26_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_27_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_27_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_28_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 fill_28_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_29_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_29_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_29_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_30_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_30_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_30_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_31_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_31_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_32_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 fill_32_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_73 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_26_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_26_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_27_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_27_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_28_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_28_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_29_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_29_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_30_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_30_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_31_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_31_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_32_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_32_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_72 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_73 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_74 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_75 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_76 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_77 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_78 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_79 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_80 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_81 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_82 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_83 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_84 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_85 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_86 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_87 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_88 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_89 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_90 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_91 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_92 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_93 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_94 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_95 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_96 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_97 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_98 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_99 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_100 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_101 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_103 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_104 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_106 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_107 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_109 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_110 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_112 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_113 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_115 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_116 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_118 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_119 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_121 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_122 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_124 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_125 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_72 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_75 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_78 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_81 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_84 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_87 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_90 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_93 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_96 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_99 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_129 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_132 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_135 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_138 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_141 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_0_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_145 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_1_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_1_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_1_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_1_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_1_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_1_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_1_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_1_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_1_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_1_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_1_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_1_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_1_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_1_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_1_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_1_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_1_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_1_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_1_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_1_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_1_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_1_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_1_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_1_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_1_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_1_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_1_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_1_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_1_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_2_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_2_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_2_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_2_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_2_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_2_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_2_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_2_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_2_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_2_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_2_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_2_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_2_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_2_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_2_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_2_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_2_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_2_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_2_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_2_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_2_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_2_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_2_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_2_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_2_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_2_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_2_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_2_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_2_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_2_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_3_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_3_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_3_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_3_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_3_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_3_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_3_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_3_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_3_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_3_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_3_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_3_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_3_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_3_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_3_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_3_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_3_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_3_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_3_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_3_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_3_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_3_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_3_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_3_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_3_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_3_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_3_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_3_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_3_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_3_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_4_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_4_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_4_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_4_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_4_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_4_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_4_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_4_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_4_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_4_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_4_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_4_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_4_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_4_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_4_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_4_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_4_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_4_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_4_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_4_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_4_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_4_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_4_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_4_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_4_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_4_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_4_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_4_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_4_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 fill_4_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_5_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_5_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_5_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_5_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_5_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_5_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_5_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_5_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_5_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_5_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_5_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_5_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_5_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_5_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_5_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_5_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_5_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_5_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_5_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_5_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_5_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_5_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_5_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_5_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_5_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_5_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_5_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_5_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_5_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_5_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_6_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_6_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_6_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_6_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_6_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_6_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_6_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_6_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_6_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_6_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_6_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_6_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_6_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_6_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_6_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_6_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_6_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_6_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_6_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_6_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_6_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_6_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_6_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_6_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_6_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_6_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_6_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_6_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_6_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_6_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_7_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_7_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_7_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_7_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_7_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_7_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_7_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_7_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_7_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_7_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_7_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_7_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_7_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_7_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_7_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_7_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_7_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_7_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_7_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_7_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_7_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_7_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_7_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_7_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_7_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_7_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_7_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_7_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_7_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 fill_7_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_8_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_8_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_8_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_8_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_8_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_8_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_8_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_8_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_8_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_8_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_8_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_8_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_8_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_8_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_8_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_8_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_8_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_8_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_8_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_8_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_8_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_8_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_8_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_8_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_8_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_8_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_8_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_8_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_8_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_8_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_9_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_9_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_9_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_9_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_9_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_9_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_9_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_9_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_9_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_9_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_9_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_9_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_9_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_9_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_9_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_9_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_9_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_9_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_9_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_9_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_9_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_9_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_9_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_9_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_9_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_9_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_9_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 fill_9_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_9_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_9_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_10_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_10_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_10_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_10_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_10_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_10_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_10_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_10_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_10_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_10_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_10_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_10_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_10_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_10_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_10_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_10_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_10_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_10_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_10_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_10_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_10_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_10_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_10_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_10_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_10_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_10_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_10_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_10_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_10_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_10_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_11_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_11_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_11_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_11_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_11_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_11_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_11_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_11_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_11_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_11_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_11_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_11_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_11_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_11_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_11_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_11_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_11_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_11_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_11_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_11_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_11_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_11_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_11_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_11_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_11_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_11_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_11_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_11_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_11_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_11_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_12_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_12_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_12_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_12_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_12_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_12_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_12_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_12_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_12_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_12_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_12_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_12_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_12_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_12_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_12_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_12_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_12_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_12_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_12_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_12_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_12_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_12_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_12_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_12_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_12_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_12_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_12_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_12_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_12_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 fill_12_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_13_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_13_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_13_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_13_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_13_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_13_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_13_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_13_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_13_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_13_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_13_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_13_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_13_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_13_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_13_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_13_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_13_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_13_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_13_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_13_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_13_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_13_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_13_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_13_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_13_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_13_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_13_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_13_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_13_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_13_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_14_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_14_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_14_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_14_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_14_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_14_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_14_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_14_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_14_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_14_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_14_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_14_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_14_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_14_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_14_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_14_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_14_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_14_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_14_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_14_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_14_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_14_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_14_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_14_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_14_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_14_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_14_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_14_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_14_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_14_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_14_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_15_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_15_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_15_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_15_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_15_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_15_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_15_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_15_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_15_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_15_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_15_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_15_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_15_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_15_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_15_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_15_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_15_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_15_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_15_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_15_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_15_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_15_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_15_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_15_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_15_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_15_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_15_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_15_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_15_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_15_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_15_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_16_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_16_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_16_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_16_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_16_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_16_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_16_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_16_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_16_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_16_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_16_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_16_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_16_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_16_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_16_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_16_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_16_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_16_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_16_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_16_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_16_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_16_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_16_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_16_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_16_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_16_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_16_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_16_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_16_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 fill_16_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_18_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_18_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_18_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_18_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_18_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_18_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_18_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_18_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_18_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_18_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_19_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_19_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_19_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_19_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_19_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_19_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_19_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_19_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_19_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_19_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_19_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_19_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_19_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_19_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_19_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_19_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_19_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_19_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_19_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_19_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_19_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_19_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_19_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_19_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_19_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_19_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_19_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_19_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_19_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_19_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_20_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_20_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_20_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_20_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_20_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_20_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_20_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_20_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_20_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_20_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_20_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_20_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_20_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_20_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_20_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_20_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_20_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_20_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_20_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_20_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_20_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_20_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_20_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_20_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_20_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_20_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_20_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_20_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_20_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 fill_20_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_21_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_21_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_21_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_21_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_21_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_21_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_21_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_21_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_21_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_21_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_21_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_21_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_21_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_21_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_21_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_21_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_21_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_21_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_21_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_21_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_21_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_21_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_21_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_21_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_21_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_21_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_21_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_21_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_21_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_21_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_22_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_22_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_22_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_22_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_22_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_22_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_22_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_22_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_22_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_22_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_22_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_22_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_22_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_22_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_22_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_22_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_22_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_22_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_22_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_22_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_22_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_22_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_22_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_22_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_22_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_22_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_22_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_22_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_22_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_22_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_22_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_23_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_23_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_23_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_23_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_23_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_23_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_23_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_23_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_23_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_23_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_23_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_23_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_23_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_23_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_23_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_23_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_23_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_23_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_23_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_23_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_23_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_23_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_23_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_23_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_23_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_23_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_23_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_23_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_23_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_23_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_23_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_24_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_24_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_24_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_24_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_24_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_24_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_24_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_24_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_24_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_24_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_24_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_24_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_24_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_24_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_24_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_24_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_24_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_24_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_24_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_24_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_24_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_24_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_24_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_24_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_24_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_24_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_24_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_24_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_24_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 fill_24_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_25_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_25_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_25_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_25_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_25_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_25_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_25_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_25_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_25_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_25_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_25_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_25_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_25_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_25_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_25_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_25_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_25_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_25_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_25_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_25_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_25_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_25_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_25_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_25_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_25_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_25_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_25_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_25_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_25_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 fill_25_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_25_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_26_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_26_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_26_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_26_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_26_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_26_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_26_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_26_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_26_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_26_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_26_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_26_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_26_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_26_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_26_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_26_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_26_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_26_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_26_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_26_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_26_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_26_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_26_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_26_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_26_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_26_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_26_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_26_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_26_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 fill_26_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 fill_26_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_27_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_27_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_27_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_27_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_27_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_27_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_27_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_27_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_27_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_27_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_27_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_27_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_27_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_27_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_27_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_27_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_27_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_27_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_27_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_27_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_27_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_27_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_27_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_27_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_27_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_27_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_27_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_27_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_27_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_27_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 fill_27_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_28_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_28_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_28_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_28_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_28_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_28_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_28_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_28_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_28_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_28_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_28_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_28_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_28_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_28_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_28_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_28_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_28_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_28_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_28_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_28_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_28_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_28_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_28_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_28_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_28_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_28_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_28_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_28_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_28_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_28_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_28_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_29_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_29_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_29_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_29_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_29_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_29_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_29_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_29_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_29_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_29_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_29_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_29_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_29_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_29_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_29_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_29_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_29_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_29_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_29_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_29_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_29_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_29_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_29_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_29_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_29_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_29_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_29_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_29_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_29_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_29_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_29_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_29_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_30_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_30_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_30_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_30_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_30_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_30_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_30_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_30_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_30_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_30_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_30_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_30_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_30_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_30_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_30_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_30_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_30_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_30_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_30_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_30_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_30_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_30_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_30_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_30_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_30_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_30_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_30_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_30_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_30_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_30_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 fill_30_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_31_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_31_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_31_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_31_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_31_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_31_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_31_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_31_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_31_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_31_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_31_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_31_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_31_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_31_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_31_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_31_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_31_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_31_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_31_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_31_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_31_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_31_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_31_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_31_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_31_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_31_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_31_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_31_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_31_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_31_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 fill_31_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_32_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_32_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_32_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_32_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_32_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_32_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_32_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_32_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_32_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_32_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_32_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_32_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_32_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_32_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_32_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_32_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_32_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_32_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_32_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_32_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_32_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_32_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_32_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_32_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_32_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_32_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_32_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_32_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_32_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_32_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 fill_32_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_32_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_72 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_75 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_78 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_81 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_84 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_87 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_90 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_93 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_96 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_99 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_129 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_132 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_135 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_138 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_141 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_144 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_147 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_150 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_153 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_33_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 fill_33_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
endmodule
