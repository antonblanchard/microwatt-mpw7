* NGSPICE file created from multiply_add_64x64.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fa_1 abstract view
.subckt sky130_fd_sc_hd__fa_1 A B CIN VGND VNB VPB VPWR COUT SUM
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ha_1 abstract view
.subckt sky130_fd_sc_hd__ha_1 A B VGND VNB VPB VPWR COUT SUM
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fa_2 abstract view
.subckt sky130_fd_sc_hd__fa_2 A B CIN VGND VNB VPB VPWR COUT SUM
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ha_2 abstract view
.subckt sky130_fd_sc_hd__ha_2 A B VGND VNB VPB VPWR COUT SUM
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

.subckt multiply_add_64x64 VGND VPWR a[0] a[10] a[11] a[12] a[13] a[14] a[15] a[16]
+ a[17] a[18] a[19] a[1] a[20] a[21] a[22] a[23] a[24] a[25] a[26] a[27] a[28] a[29]
+ a[2] a[30] a[31] a[32] a[33] a[34] a[35] a[36] a[37] a[38] a[39] a[3] a[40] a[41]
+ a[42] a[43] a[44] a[45] a[46] a[47] a[48] a[49] a[4] a[50] a[51] a[52] a[53] a[54]
+ a[55] a[56] a[57] a[58] a[59] a[5] a[60] a[61] a[62] a[63] a[6] a[7] a[8] a[9] b[0]
+ b[10] b[11] b[12] b[13] b[14] b[15] b[16] b[17] b[18] b[19] b[1] b[20] b[21] b[22]
+ b[23] b[24] b[25] b[26] b[27] b[28] b[29] b[2] b[30] b[31] b[32] b[33] b[34] b[35]
+ b[36] b[37] b[38] b[39] b[3] b[40] b[41] b[42] b[43] b[44] b[45] b[46] b[47] b[48]
+ b[49] b[4] b[50] b[51] b[52] b[53] b[54] b[55] b[56] b[57] b[58] b[59] b[5] b[60]
+ b[61] b[62] b[63] b[6] b[7] b[8] b[9] c[0] c[100] c[101] c[102] c[103] c[104] c[105]
+ c[106] c[107] c[108] c[109] c[10] c[110] c[111] c[112] c[113] c[114] c[115] c[116]
+ c[117] c[118] c[119] c[11] c[120] c[121] c[122] c[123] c[124] c[125] c[126] c[127]
+ c[12] c[13] c[14] c[15] c[16] c[17] c[18] c[19] c[1] c[20] c[21] c[22] c[23] c[24]
+ c[25] c[26] c[27] c[28] c[29] c[2] c[30] c[31] c[32] c[33] c[34] c[35] c[36] c[37]
+ c[38] c[39] c[3] c[40] c[41] c[42] c[43] c[44] c[45] c[46] c[47] c[48] c[49] c[4]
+ c[50] c[51] c[52] c[53] c[54] c[55] c[56] c[57] c[58] c[59] c[5] c[60] c[61] c[62]
+ c[63] c[64] c[65] c[66] c[67] c[68] c[69] c[6] c[70] c[71] c[72] c[73] c[74] c[75]
+ c[76] c[77] c[78] c[79] c[7] c[80] c[81] c[82] c[83] c[84] c[85] c[86] c[87] c[88]
+ c[89] c[8] c[90] c[91] c[92] c[93] c[94] c[95] c[96] c[97] c[98] c[99] c[9] clk
+ o[0] o[100] o[101] o[102] o[103] o[104] o[105] o[106] o[107] o[108] o[109] o[10]
+ o[110] o[111] o[112] o[113] o[114] o[115] o[116] o[117] o[118] o[119] o[11] o[120]
+ o[121] o[122] o[123] o[124] o[125] o[126] o[127] o[12] o[13] o[14] o[15] o[16] o[17]
+ o[18] o[19] o[1] o[20] o[21] o[22] o[23] o[24] o[25] o[26] o[27] o[28] o[29] o[2]
+ o[30] o[31] o[32] o[33] o[34] o[35] o[36] o[37] o[38] o[39] o[3] o[40] o[41] o[42]
+ o[43] o[44] o[45] o[46] o[47] o[48] o[49] o[4] o[50] o[51] o[52] o[53] o[54] o[55]
+ o[56] o[57] o[58] o[59] o[5] o[60] o[61] o[62] o[63] o[64] o[65] o[66] o[67] o[68]
+ o[69] o[6] o[70] o[71] o[72] o[73] o[74] o[75] o[76] o[77] o[78] o[79] o[7] o[80]
+ o[81] o[82] o[83] o[84] o[85] o[86] o[87] o[88] o[89] o[8] o[90] o[91] o[92] o[93]
+ o[94] o[95] o[96] o[97] o[98] o[99] o[9] rst
XFILLER_39_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0367_ clknet_leaf_190_clk booth_b44_m31 VGND VGND VPWR VPWR pp_row75_17 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_57_8 c$16 s$19 s$21 VGND VGND VPWR VPWR c$490 s$491 sky130_fd_sc_hd__fa_1
XFILLER_95_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2106_ clknet_leaf_33_clk booth_b46_m12 VGND VGND VPWR VPWR pp_row58_23 sky130_fd_sc_hd__dfxtp_1
X_0298_ clknet_leaf_201_clk booth_b36_m37 VGND VGND VPWR VPWR pp_row73_14 sky130_fd_sc_hd__dfxtp_1
X_2037_ clknet_leaf_83_clk booth_b46_m10 VGND VGND VPWR VPWR pp_row56_23 sky130_fd_sc_hd__dfxtp_1
XFILLER_82_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_104_0 net1906 pp_row104_1 pp_row104_2 VGND VGND VPWR VPWR c$1956 s$1957
+ sky130_fd_sc_hd__fa_1
XFILLER_35_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_606 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1290 t$5064 net1663 VGND VGND VPWR VPWR booth_b18_m25 sky130_fd_sc_hd__xor2_1
XFILLER_167_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_90_2 pp_row90_6 pp_row90_7 pp_row90_8 VGND VGND VPWR VPWR c$1022 s$1023
+ sky130_fd_sc_hd__fa_1
XFILLER_191_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_83_1 pp_row83_3 pp_row83_4 pp_row83_5 VGND VGND VPWR VPWR c$940 s$941
+ sky130_fd_sc_hd__fa_1
XFILLER_104_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_60_0 s$1457 c$2310 c$2312 VGND VGND VPWR VPWR c$3050 s$3051 sky130_fd_sc_hd__fa_1
XFILLER_131_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout820 net821 VGND VGND VPWR VPWR net820 sky130_fd_sc_hd__buf_4
XFILLER_89_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_76_0 pp_row76_5 pp_row76_6 pp_row76_7 VGND VGND VPWR VPWR c$816 s$817
+ sky130_fd_sc_hd__fa_1
XFILLER_104_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout831 net832 VGND VGND VPWR VPWR net831 sky130_fd_sc_hd__buf_4
XFILLER_120_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout842 net843 VGND VGND VPWR VPWR net842 sky130_fd_sc_hd__buf_6
Xfanout853 net854 VGND VGND VPWR VPWR net853 sky130_fd_sc_hd__clkbuf_4
Xfanout864 net865 VGND VGND VPWR VPWR net864 sky130_fd_sc_hd__buf_4
XFILLER_131_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout875 net877 VGND VGND VPWR VPWR net875 sky130_fd_sc_hd__buf_4
XFILLER_58_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout886 net888 VGND VGND VPWR VPWR net886 sky130_fd_sc_hd__buf_4
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout897 net898 VGND VGND VPWR VPWR net897 sky130_fd_sc_hd__clkbuf_4
XU$$3609 t$6249 net1319 VGND VGND VPWR VPWR booth_b52_m20 sky130_fd_sc_hd__xor2_1
XTAP_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2908 t$5891 net1372 VGND VGND VPWR VPWR booth_b42_m12 sky130_fd_sc_hd__xor2_1
XFILLER_172_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_202 net1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2919 net1151 net519 net1140 net792 VGND VGND VPWR VPWR t$5897 sky130_fd_sc_hd__a22o_1
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_213 net1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_224 net1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_ha_5_124_1 pp_row124_3 pp_row124_4 VGND VGND VPWR VPWR c$3894 s$3895 sky130_fd_sc_hd__ha_1
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_235 net1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_246 net1559 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_257 net1640 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_268 net1728 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_279 c$4242 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_98_1 c$1894 c$1896 c$1898 VGND VGND VPWR VPWR c$2624 s$2625 sky130_fd_sc_hd__fa_1
Xdadda_fa_6_75_0 c$3692 c$3694 s$3697 VGND VGND VPWR VPWR c$4046 s$4047 sky130_fd_sc_hd__fa_1
XFILLER_142_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1270_ clknet_leaf_10_clk booth_b16_m10 VGND VGND VPWR VPWR pp_row26_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_1_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0221_ clknet_leaf_200_clk booth_b18_m53 VGND VGND VPWR VPWR pp_row71_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_76_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$370 net1724 net533 net1715 net806 VGND VGND VPWR VPWR t$4594 sky130_fd_sc_hd__a22o_1
XU$$381 t$4599 net1280 VGND VGND VPWR VPWR booth_b4_m50 sky130_fd_sc_hd__xor2_1
XU$$392 net1614 net530 net1606 net803 VGND VGND VPWR VPWR t$4605 sky130_fd_sc_hd__a22o_1
XFILLER_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0985_ clknet_leaf_117_clk booth_b46_m54 VGND VGND VPWR VPWR pp_row100_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_93_0 pp_row93_6 pp_row93_7 pp_row93_8 VGND VGND VPWR VPWR c$1842 s$1843
+ sky130_fd_sc_hd__fa_1
XFILLER_156_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1606_ clknet_leaf_240_clk booth_b10_m32 VGND VGND VPWR VPWR pp_row42_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_160_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1537_ clknet_leaf_7_clk booth_b18_m21 VGND VGND VPWR VPWR pp_row39_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_59_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1468_ clknet_leaf_40_clk booth_b20_m16 VGND VGND VPWR VPWR pp_row36_10 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_62_6 c$52 c$54 c$56 VGND VGND VPWR VPWR c$576 s$577 sky130_fd_sc_hd__fa_1
XFILLER_74_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0419_ clknet_leaf_145_clk booth_b26_m51 VGND VGND VPWR VPWR pp_row77_7 sky130_fd_sc_hd__dfxtp_1
X_1399_ clknet_leaf_54_clk booth_b8_m25 VGND VGND VPWR VPWR pp_row33_4 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_55_5 pp_row55_20 pp_row55_21 pp_row55_22 VGND VGND VPWR VPWR c$448 s$449
+ sky130_fd_sc_hd__fa_1
XFILLER_55_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_48_4 pp_row48_12 pp_row48_13 pp_row48_14 VGND VGND VPWR VPWR c$324 s$325
+ sky130_fd_sc_hd__fa_1
XFILLER_27_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_18_2 s$1987 s$1989 s$1991 VGND VGND VPWR VPWR c$2802 s$2803 sky130_fd_sc_hd__fa_1
XFILLER_179_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_92_0 s$3767 c$4078 s$4081 VGND VGND VPWR VPWR c$4336 s$4337 sky130_fd_sc_hd__fa_1
XFILLER_163_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1604 net1606 VGND VGND VPWR VPWR net1604 sky130_fd_sc_hd__buf_4
XFILLER_77_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1615 net1619 VGND VGND VPWR VPWR net1615 sky130_fd_sc_hd__buf_4
Xfanout1626 net1627 VGND VGND VPWR VPWR net1626 sky130_fd_sc_hd__buf_4
Xfanout1637 net113 VGND VGND VPWR VPWR net1637 sky130_fd_sc_hd__buf_4
Xfanout650 sel_0$4967 VGND VGND VPWR VPWR net650 sky130_fd_sc_hd__buf_6
Xfanout1648 net111 VGND VGND VPWR VPWR net1648 sky130_fd_sc_hd__buf_6
XFILLER_77_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout661 net666 VGND VGND VPWR VPWR net661 sky130_fd_sc_hd__buf_4
XU$$4107 net1529 net453 net1804 net726 VGND VGND VPWR VPWR t$6503 sky130_fd_sc_hd__a22o_1
Xfanout1659 net1661 VGND VGND VPWR VPWR net1659 sky130_fd_sc_hd__clkbuf_8
XU$$4118 net1229 net434 net1125 net716 VGND VGND VPWR VPWR t$6510 sky130_fd_sc_hd__a22o_1
Xfanout672 net673 VGND VGND VPWR VPWR net672 sky130_fd_sc_hd__buf_4
XU$$4129 t$6515 net1269 VGND VGND VPWR VPWR booth_b60_m6 sky130_fd_sc_hd__xor2_1
Xfanout683 sel_1$4688 VGND VGND VPWR VPWR net683 sky130_fd_sc_hd__buf_6
XFILLER_120_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout694 net695 VGND VGND VPWR VPWR net694 sky130_fd_sc_hd__buf_4
XFILLER_19_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3406 net1618 net498 net1609 net771 VGND VGND VPWR VPWR t$6145 sky130_fd_sc_hd__a22o_1
XFILLER_58_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3417 t$6150 net1345 VGND VGND VPWR VPWR booth_b48_m61 sky130_fd_sc_hd__xor2_1
XFILLER_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3428 net1330 notblock$6155\[1\] VGND VGND VPWR VPWR t$6156 sky130_fd_sc_hd__and2_1
XTAP_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3439 net938 net488 net1677 net761 VGND VGND VPWR VPWR t$6163 sky130_fd_sc_hd__a22o_1
XFILLER_46_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_854 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2705 net1696 net545 net1688 net818 VGND VGND VPWR VPWR t$5787 sky130_fd_sc_hd__a22o_1
XTAP_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2716 t$5792 net1401 VGND VGND VPWR VPWR booth_b38_m53 sky130_fd_sc_hd__xor2_1
XU$$2727 net1592 net548 net1584 net821 VGND VGND VPWR VPWR t$5798 sky130_fd_sc_hd__a22o_1
XFILLER_160_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2738 t$5803 net1401 VGND VGND VPWR VPWR booth_b38_m64 sky130_fd_sc_hd__xor2_1
XFILLER_46_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2749 t$5810 net1376 VGND VGND VPWR VPWR booth_b40_m1 sky130_fd_sc_hd__xor2_1
XFILLER_61_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_20_2 pp_row20_6 pp_row20_7 pp_row20_8 VGND VGND VPWR VPWR c$2002 s$2003
+ sky130_fd_sc_hd__fa_1
XTAP_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_987 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_773 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_929 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0770_ clknet_leaf_138_clk booth_b28_m62 VGND VGND VPWR VPWR pp_row90_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_183_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2440_ clknet_leaf_75_clk booth_b58_m9 VGND VGND VPWR VPWR pp_row67_29 sky130_fd_sc_hd__dfxtp_1
XFILLER_170_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2371_ clknet_leaf_85_clk booth_b2_m64 VGND VGND VPWR VPWR pp_row66_1 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_72_5 s$755 s$757 s$759 VGND VGND VPWR VPWR c$1600 s$1601 sky130_fd_sc_hd__fa_2
XFILLER_97_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1322_ clknet_leaf_0_clk booth_b12_m17 VGND VGND VPWR VPWR pp_row29_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_69_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_65_4 s$623 s$625 s$627 VGND VGND VPWR VPWR c$1514 s$1515 sky130_fd_sc_hd__fa_2
XFILLER_111_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1253_ clknet_leaf_10_clk booth_b12_m13 VGND VGND VPWR VPWR pp_row25_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_58_3 c$490 s$493 s$495 VGND VGND VPWR VPWR c$1428 s$1429 sky130_fd_sc_hd__fa_1
XFILLER_110_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0204_ clknet_leaf_152_clk booth_b48_m22 VGND VGND VPWR VPWR pp_row70_22 sky130_fd_sc_hd__dfxtp_1
X_1184_ clknet_leaf_53_clk booth_b20_m0 VGND VGND VPWR VPWR pp_row20_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_37_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3940 net1693 net466 net1684 net739 VGND VGND VPWR VPWR t$6418 sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_28_1 s$2859 s$2861 s$2863 VGND VGND VPWR VPWR c$3510 s$3511 sky130_fd_sc_hd__fa_1
XU$$3951 t$6423 net1297 VGND VGND VPWR VPWR booth_b56_m54 sky130_fd_sc_hd__xor2_1
XU$$3962 net1584 net465 net1557 net738 VGND VGND VPWR VPWR t$6429 sky130_fd_sc_hd__a22o_1
XU$$3973 net1292 VGND VGND VPWR VPWR notblock$6435\[0\] sky130_fd_sc_hd__inv_1
XU$$3984 t$6441 net1282 VGND VGND VPWR VPWR booth_b58_m2 sky130_fd_sc_hd__xor2_1
XU$$3995 net1517 net455 net1510 net728 VGND VGND VPWR VPWR t$6447 sky130_fd_sc_hd__a22o_1
XFILLER_91_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0968_ clknet_leaf_116_clk booth_b46_m53 VGND VGND VPWR VPWR pp_row99_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_118_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_102_1 s$3303 s$3305 s$3307 VGND VGND VPWR VPWR c$3806 s$3807 sky130_fd_sc_hd__fa_1
XFILLER_118_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0899_ clknet_leaf_130_clk booth_b62_m58 VGND VGND VPWR VPWR pp_row120_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_160_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput264 net264 VGND VGND VPWR VPWR o[106] sky130_fd_sc_hd__buf_2
XFILLER_161_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput275 net275 VGND VGND VPWR VPWR o[116] sky130_fd_sc_hd__buf_2
XFILLER_0_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput286 net286 VGND VGND VPWR VPWR o[126] sky130_fd_sc_hd__buf_2
Xoutput297 net297 VGND VGND VPWR VPWR o[20] sky130_fd_sc_hd__buf_2
XFILLER_59_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_60_3 pp_row60_23 pp_row60_24 pp_row60_25 VGND VGND VPWR VPWR c$534 s$535
+ sky130_fd_sc_hd__fa_1
XFILLER_28_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_53_2 pp_row53_8 pp_row53_9 pp_row53_10 VGND VGND VPWR VPWR c$406 s$407
+ sky130_fd_sc_hd__fa_1
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_30_1 c$2074 c$2076 s$2079 VGND VGND VPWR VPWR c$2872 s$2873 sky130_fd_sc_hd__fa_1
Xdadda_fa_1_46_1 pp_row46_3 pp_row46_4 pp_row46_5 VGND VGND VPWR VPWR c$290 s$291
+ sky130_fd_sc_hd__fa_2
XFILLER_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_23_0 s$1053 c$2014 c$2016 VGND VGND VPWR VPWR c$2828 s$2829 sky130_fd_sc_hd__fa_1
Xdadda_fa_1_39_0 pp_row39_0 pp_row39_1 pp_row39_2 VGND VGND VPWR VPWR c$222 s$223
+ sky130_fd_sc_hd__fa_1
XFILLER_70_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_973 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_75_3 s$1631 s$1633 s$1635 VGND VGND VPWR VPWR c$2444 s$2445 sky130_fd_sc_hd__fa_1
XFILLER_140_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1401 net1402 VGND VGND VPWR VPWR net1401 sky130_fd_sc_hd__buf_4
Xfanout1412 net3 VGND VGND VPWR VPWR net1412 sky130_fd_sc_hd__buf_6
Xdadda_fa_3_68_2 c$1540 s$1543 s$1545 VGND VGND VPWR VPWR c$2386 s$2387 sky130_fd_sc_hd__fa_1
Xfanout1423 net1424 VGND VGND VPWR VPWR net1423 sky130_fd_sc_hd__buf_6
XFILLER_120_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1434 net1436 VGND VGND VPWR VPWR net1434 sky130_fd_sc_hd__buf_6
Xfanout1445 net1446 VGND VGND VPWR VPWR net1445 sky130_fd_sc_hd__buf_8
XFILLER_78_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1456 net22 VGND VGND VPWR VPWR net1456 sky130_fd_sc_hd__buf_6
Xfanout1467 net1468 VGND VGND VPWR VPWR net1467 sky130_fd_sc_hd__buf_4
XFILLER_171_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout480 net481 VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__buf_4
Xfanout1478 net1480 VGND VGND VPWR VPWR net1478 sky130_fd_sc_hd__buf_6
Xfanout1489 net1490 VGND VGND VPWR VPWR net1489 sky130_fd_sc_hd__buf_6
Xfanout491 net492 VGND VGND VPWR VPWR net491 sky130_fd_sc_hd__buf_2
Xdadda_fa_6_38_0 c$3544 c$3546 s$3549 VGND VGND VPWR VPWR c$3972 s$3973 sky130_fd_sc_hd__fa_1
XU$$3203 net1104 net506 net1096 net779 VGND VGND VPWR VPWR t$6042 sky130_fd_sc_hd__a22o_1
XU$$3214 t$6047 net1348 VGND VGND VPWR VPWR booth_b46_m28 sky130_fd_sc_hd__xor2_1
XU$$3225 net994 net504 net985 net777 VGND VGND VPWR VPWR t$6053 sky130_fd_sc_hd__a22o_1
XFILLER_185_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3236 t$6058 net1351 VGND VGND VPWR VPWR booth_b46_m39 sky130_fd_sc_hd__xor2_1
XFILLER_46_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2502 net1180 net554 net1171 net827 VGND VGND VPWR VPWR t$5684 sky130_fd_sc_hd__a22o_1
XU$$3247 net1726 net507 net1717 net780 VGND VGND VPWR VPWR t$6064 sky130_fd_sc_hd__a22o_1
XFILLER_47_876 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$18 c$4186 s$4189 VGND VGND VPWR VPWR final_adder.$signal$38 final_adder.$signal$1108
+ sky130_fd_sc_hd__ha_1
XU$$3258 t$6069 net1355 VGND VGND VPWR VPWR booth_b46_m50 sky130_fd_sc_hd__xor2_1
XU$$2513 t$5689 net1406 VGND VGND VPWR VPWR booth_b36_m20 sky130_fd_sc_hd__xor2_1
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$29 c$4208 s$4211 VGND VGND VPWR VPWR final_adder.$signal$60 final_adder.$signal$1119
+ sky130_fd_sc_hd__ha_1
XU$$2524 net1078 net555 net1070 net828 VGND VGND VPWR VPWR t$5695 sky130_fd_sc_hd__a22o_1
XU$$3269 net1618 net507 net1609 net780 VGND VGND VPWR VPWR t$6075 sky130_fd_sc_hd__a22o_1
XFILLER_185_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2535 t$5700 net1407 VGND VGND VPWR VPWR booth_b36_m31 sky130_fd_sc_hd__xor2_1
XU$$1801 net1524 net597 net1516 net870 VGND VGND VPWR VPWR t$5326 sky130_fd_sc_hd__a22o_1
XFILLER_146_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2546 net965 net553 net957 net826 VGND VGND VPWR VPWR t$5706 sky130_fd_sc_hd__a22o_1
XFILLER_146_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2557 t$5711 net1408 VGND VGND VPWR VPWR booth_b36_m42 sky130_fd_sc_hd__xor2_1
XFILLER_73_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1812 t$5331 net1460 VGND VGND VPWR VPWR booth_b26_m12 sky130_fd_sc_hd__xor2_1
XFILLER_181_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2568 net1696 net556 net1688 net829 VGND VGND VPWR VPWR t$5717 sky130_fd_sc_hd__a22o_1
XU$$1823 net1147 net594 net1139 net867 VGND VGND VPWR VPWR t$5337 sky130_fd_sc_hd__a22o_1
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2579 t$5722 net1409 VGND VGND VPWR VPWR booth_b36_m53 sky130_fd_sc_hd__xor2_1
XU$$1834 t$5342 net1458 VGND VGND VPWR VPWR booth_b26_m23 sky130_fd_sc_hd__xor2_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1845 net1049 net597 net1042 net870 VGND VGND VPWR VPWR t$5348 sky130_fd_sc_hd__a22o_1
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1856 t$5353 net1462 VGND VGND VPWR VPWR booth_b26_m34 sky130_fd_sc_hd__xor2_1
X_1940_ clknet_leaf_70_clk booth_b44_m9 VGND VGND VPWR VPWR pp_row53_22 sky130_fd_sc_hd__dfxtp_1
XFILLER_61_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1867 net944 net597 net928 net870 VGND VGND VPWR VPWR t$5359 sky130_fd_sc_hd__a22o_1
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1878 t$5364 net1464 VGND VGND VPWR VPWR booth_b26_m45 sky130_fd_sc_hd__xor2_1
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1889 net1659 net600 net1647 net873 VGND VGND VPWR VPWR t$5370 sky130_fd_sc_hd__a22o_1
XFILLER_187_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1871_ clknet_leaf_72_clk booth_b32_m19 VGND VGND VPWR VPWR pp_row51_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_187_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0822_ clknet_leaf_106_clk booth_b40_m52 VGND VGND VPWR VPWR pp_row92_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_80_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0753_ clknet_leaf_160_clk booth_b40_m49 VGND VGND VPWR VPWR pp_row89_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_192_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0684_ clknet_leaf_174_clk booth_b50_m36 VGND VGND VPWR VPWR pp_row86_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_192_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2423_ clknet_leaf_142_clk booth_b28_m39 VGND VGND VPWR VPWR pp_row67_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_130_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_70_2 c$700 c$702 c$704 VGND VGND VPWR VPWR c$1570 s$1571 sky130_fd_sc_hd__fa_2
X_2354_ clknet_leaf_75_clk booth_b38_m27 VGND VGND VPWR VPWR pp_row65_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_69_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_63_1 c$568 c$570 c$572 VGND VGND VPWR VPWR c$1484 s$1485 sky130_fd_sc_hd__fa_1
XFILLER_57_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1305_ clknet_leaf_122_clk booth_b62_m41 VGND VGND VPWR VPWR pp_row103_12 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$508 final_adder.p_new$520 final_adder.p_new$512 VGND VGND VPWR VPWR
+ final_adder.p_new$636 sky130_fd_sc_hd__and2_1
XFILLER_84_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_40_0 c$2924 c$2926 c$2928 VGND VGND VPWR VPWR c$3556 s$3557 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$519 final_adder.p_new$522 final_adder.g_new$531 final_adder.g_new$523
+ VGND VGND VPWR VPWR final_adder.g_new$647 sky130_fd_sc_hd__a21o_1
X_2285_ clknet_leaf_152_clk booth_b44_m19 VGND VGND VPWR VPWR pp_row63_22 sky130_fd_sc_hd__dfxtp_1
XFILLER_85_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_56_0 s$17 c$438 c$440 VGND VGND VPWR VPWR c$1398 s$1399 sky130_fd_sc_hd__fa_2
X_1236_ clknet_leaf_13_clk booth_b12_m12 VGND VGND VPWR VPWR pp_row24_6 sky130_fd_sc_hd__dfxtp_1
XU$$4460 net989 sel_0$6647 net980 net697 VGND VGND VPWR VPWR t$6684 sky130_fd_sc_hd__a22o_1
XU$$4471 t$6689 net1856 VGND VGND VPWR VPWR booth_b64_m40 sky130_fd_sc_hd__xor2_1
XFILLER_65_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4482 net1719 sel_0$6647 net1710 net699 VGND VGND VPWR VPWR t$6695 sky130_fd_sc_hd__a22o_1
XU$$4493 t$6700 net1867 VGND VGND VPWR VPWR booth_b64_m51 sky130_fd_sc_hd__xor2_1
XFILLER_64_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1167_ clknet_leaf_45_clk booth_b14_m5 VGND VGND VPWR VPWR pp_row19_7 sky130_fd_sc_hd__dfxtp_1
XU$$4427_1834 VGND VGND VPWR VPWR U$$4427_1834/HI net1834 sky130_fd_sc_hd__conb_1
XU$$3770 t$6331 net1303 VGND VGND VPWR VPWR booth_b54_m32 sky130_fd_sc_hd__xor2_1
XU$$3781 net962 net474 net953 net747 VGND VGND VPWR VPWR t$6337 sky130_fd_sc_hd__a22o_1
XU$$3792 t$6342 net1307 VGND VGND VPWR VPWR booth_b54_m43 sky130_fd_sc_hd__xor2_1
XFILLER_53_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1098_ clknet_leaf_59_clk booth_b8_m5 VGND VGND VPWR VPWR pp_row13_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_80_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_85_2 s$2521 s$2523 s$2525 VGND VGND VPWR VPWR c$3204 s$3205 sky130_fd_sc_hd__fa_1
XFILLER_118_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_78_1 c$2458 c$2460 s$2463 VGND VGND VPWR VPWR c$3160 s$3161 sky130_fd_sc_hd__fa_1
XFILLER_0_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_55_0 s$3619 c$4004 s$4007 VGND VGND VPWR VPWR c$4262 s$4263 sky130_fd_sc_hd__fa_1
XFILLER_173_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1096 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$903 t$4866 net1317 VGND VGND VPWR VPWR booth_b12_m37 sky130_fd_sc_hd__xor2_1
XFILLER_44_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$914 net1741 net398 net1733 net664 VGND VGND VPWR VPWR t$4872 sky130_fd_sc_hd__a22o_1
XFILLER_16_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$925 t$4877 net1317 VGND VGND VPWR VPWR booth_b12_m48 sky130_fd_sc_hd__xor2_1
XFILLER_71_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$936 net1633 net399 net1623 net665 VGND VGND VPWR VPWR t$4883 sky130_fd_sc_hd__a22o_1
XFILLER_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$947 t$4888 net1316 VGND VGND VPWR VPWR booth_b12_m59 sky130_fd_sc_hd__xor2_1
XFILLER_56_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$958 net1316 VGND VGND VPWR VPWR notsign$4894 sky130_fd_sc_hd__inv_1
XU$$969 net1123 net385 net1032 net651 VGND VGND VPWR VPWR t$4901 sky130_fd_sc_hd__a22o_1
XU$$1108 net1032 net646 net933 net919 VGND VGND VPWR VPWR t$4972 sky130_fd_sc_hd__a22o_1
XFILLER_71_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1119 t$4977 net1006 VGND VGND VPWR VPWR booth_b16_m8 sky130_fd_sc_hd__xor2_1
XFILLER_19_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_80_1 c$1678 c$1680 c$1682 VGND VGND VPWR VPWR c$2480 s$2481 sky130_fd_sc_hd__fa_1
XFILLER_98_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_73_0 s$779 c$1590 c$1592 VGND VGND VPWR VPWR c$2422 s$2423 sky130_fd_sc_hd__fa_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1220 net1223 VGND VGND VPWR VPWR net1220 sky130_fd_sc_hd__buf_4
XFILLER_152_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1231 net1232 VGND VGND VPWR VPWR net1231 sky130_fd_sc_hd__clkbuf_4
XFILLER_182_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1242 net1243 VGND VGND VPWR VPWR net1242 sky130_fd_sc_hd__buf_6
Xfanout1253 net62 VGND VGND VPWR VPWR net1253 sky130_fd_sc_hd__buf_6
XFILLER_39_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1264 net58 VGND VGND VPWR VPWR net1264 sky130_fd_sc_hd__clkbuf_4
XFILLER_121_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1275 net1276 VGND VGND VPWR VPWR net1275 sky130_fd_sc_hd__buf_4
XFILLER_93_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1286 net55 VGND VGND VPWR VPWR net1286 sky130_fd_sc_hd__buf_6
XFILLER_94_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3000 t$5937 net1373 VGND VGND VPWR VPWR booth_b42_m58 sky130_fd_sc_hd__xor2_1
X_2070_ clknet_leaf_36_clk booth_b42_m15 VGND VGND VPWR VPWR pp_row57_21 sky130_fd_sc_hd__dfxtp_1
Xfanout1297 net1299 VGND VGND VPWR VPWR net1297 sky130_fd_sc_hd__buf_6
XU$$3011 net1532 net525 net1786 net798 VGND VGND VPWR VPWR t$5943 sky130_fd_sc_hd__a22o_1
XU$$3022 net1228 net511 net1124 net784 VGND VGND VPWR VPWR t$5950 sky130_fd_sc_hd__a22o_1
XU$$3033 t$5955 net1362 VGND VGND VPWR VPWR booth_b44_m6 sky130_fd_sc_hd__xor2_1
X_1021_ clknet_leaf_249_clk net168 VGND VGND VPWR VPWR pp_row1_1 sky130_fd_sc_hd__dfxtp_2
XFILLER_47_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3044 net1217 net514 net1208 net787 VGND VGND VPWR VPWR t$5961 sky130_fd_sc_hd__a22o_1
XU$$3055 t$5966 net1358 VGND VGND VPWR VPWR booth_b44_m17 sky130_fd_sc_hd__xor2_1
XU$$2310 net1613 net574 net1606 net847 VGND VGND VPWR VPWR t$5585 sky130_fd_sc_hd__a22o_1
XU$$2321 t$5590 net1437 VGND VGND VPWR VPWR booth_b32_m61 sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_102_0 s$1949 c$2646 c$2648 VGND VGND VPWR VPWR c$3302 s$3303 sky130_fd_sc_hd__fa_1
XU$$3066 net1104 net517 net1096 net790 VGND VGND VPWR VPWR t$5972 sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_35_5 pp_row35_17 pp_row35_18 c$204 VGND VGND VPWR VPWR c$1156 s$1157 sky130_fd_sc_hd__fa_1
XFILLER_19_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2332 net1426 notblock$5595\[1\] VGND VGND VPWR VPWR t$5596 sky130_fd_sc_hd__and2_1
XU$$3077 t$5977 net1357 VGND VGND VPWR VPWR booth_b44_m28 sky130_fd_sc_hd__xor2_1
XU$$2343 net932 net560 net1671 net833 VGND VGND VPWR VPWR t$5603 sky130_fd_sc_hd__a22o_1
XU$$3088 net994 net512 net985 net785 VGND VGND VPWR VPWR t$5983 sky130_fd_sc_hd__a22o_1
XFILLER_62_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3099 t$5988 net1359 VGND VGND VPWR VPWR booth_b44_m39 sky130_fd_sc_hd__xor2_1
XU$$2354 t$5608 net1420 VGND VGND VPWR VPWR booth_b34_m9 sky130_fd_sc_hd__xor2_1
XU$$1620 t$5232 net1483 VGND VGND VPWR VPWR booth_b22_m53 sky130_fd_sc_hd__xor2_1
XU$$2365 net1176 net561 net1167 net834 VGND VGND VPWR VPWR t$5614 sky130_fd_sc_hd__a22o_1
XU$$2376 t$5619 net1423 VGND VGND VPWR VPWR booth_b34_m20 sky130_fd_sc_hd__xor2_1
XU$$1631 net1588 net617 net1579 net890 VGND VGND VPWR VPWR t$5238 sky130_fd_sc_hd__a22o_1
XU$$1642 t$5243 net1481 VGND VGND VPWR VPWR booth_b22_m64 sky130_fd_sc_hd__xor2_1
XU$$2387 net1073 net561 net1065 net834 VGND VGND VPWR VPWR t$5625 sky130_fd_sc_hd__a22o_1
XU$$2398 t$5630 net1424 VGND VGND VPWR VPWR booth_b34_m31 sky130_fd_sc_hd__xor2_1
XFILLER_34_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1653 t$5250 net1466 VGND VGND VPWR VPWR booth_b24_m1 sky130_fd_sc_hd__xor2_1
XU$$1664 net1519 net602 net1511 net875 VGND VGND VPWR VPWR t$5256 sky130_fd_sc_hd__a22o_1
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1675 t$5261 net1469 VGND VGND VPWR VPWR booth_b24_m12 sky130_fd_sc_hd__xor2_1
XU$$1686 net1147 net602 net1138 net875 VGND VGND VPWR VPWR t$5267 sky130_fd_sc_hd__a22o_1
XU$$1697 t$5272 net1468 VGND VGND VPWR VPWR booth_b24_m23 sky130_fd_sc_hd__xor2_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1923_ clknet_leaf_80_clk booth_b14_m39 VGND VGND VPWR VPWR pp_row53_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_187_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_150_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_150_clk
+ sky130_fd_sc_hd__clkbuf_16
X_1854_ clknet_leaf_67_clk booth_b0_m51 VGND VGND VPWR VPWR pp_row51_0 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_95_1 s$3261 s$3263 s$3265 VGND VGND VPWR VPWR c$3778 s$3779 sky130_fd_sc_hd__fa_1
Xdadda_fa_3_112_0_1910 VGND VGND VPWR VPWR net1910 dadda_fa_3_112_0_1910/LO sky130_fd_sc_hd__conb_1
X_0805_ clknet_leaf_94_clk booth_b50_m41 VGND VGND VPWR VPWR pp_row91_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_128_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4457_1849 VGND VGND VPWR VPWR U$$4457_1849/HI net1849 sky130_fd_sc_hd__conb_1
X_1785_ clknet_leaf_222_clk booth_b38_m10 VGND VGND VPWR VPWR pp_row48_19 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_88_0 c$3212 c$3214 c$3216 VGND VGND VPWR VPWR c$3748 s$3749 sky130_fd_sc_hd__fa_2
XFILLER_7_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0736_ clknet_leaf_134_clk booth_b52_m36 VGND VGND VPWR VPWR pp_row88_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_144_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0667_ clknet_leaf_187_clk booth_b64_m21 VGND VGND VPWR VPWR pp_row85_22 sky130_fd_sc_hd__dfxtp_1
X_2406_ clknet_leaf_99_clk booth_b64_m2 VGND VGND VPWR VPWR pp_row66_32 sky130_fd_sc_hd__dfxtp_1
XFILLER_112_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0598_ clknet_leaf_188_clk booth_b38_m45 VGND VGND VPWR VPWR pp_row83_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_97_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2337_ clknet_leaf_127_clk booth_b48_m63 VGND VGND VPWR VPWR pp_row111_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_84_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$305 final_adder.p_new$304 final_adder.g_new$307 final_adder.g_new$305
+ VGND VGND VPWR VPWR final_adder.g_new$433 sky130_fd_sc_hd__a21o_1
XFILLER_97_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$316 final_adder.p_new$318 final_adder.p_new$316 VGND VGND VPWR VPWR
+ final_adder.p_new$444 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$327 final_adder.p_new$326 final_adder.g_new$329 final_adder.g_new$327
+ VGND VGND VPWR VPWR final_adder.g_new$455 sky130_fd_sc_hd__a21o_1
XTAP_3609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$338 final_adder.p_new$340 final_adder.p_new$338 VGND VGND VPWR VPWR
+ final_adder.p_new$466 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$349 final_adder.p_new$348 final_adder.g_new$351 final_adder.g_new$349
+ VGND VGND VPWR VPWR final_adder.g_new$477 sky130_fd_sc_hd__a21o_1
XFILLER_73_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2268_ clknet_leaf_214_clk booth_b16_m47 VGND VGND VPWR VPWR pp_row63_8 sky130_fd_sc_hd__dfxtp_1
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1219_ clknet_leaf_48_clk booth_b6_m17 VGND VGND VPWR VPWR pp_row23_3 sky130_fd_sc_hd__dfxtp_1
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2199_ clknet_leaf_228_clk booth_b22_m39 VGND VGND VPWR VPWR pp_row61_11 sky130_fd_sc_hd__dfxtp_1
XU$$4290 t$6597 net1256 VGND VGND VPWR VPWR booth_b62_m18 sky130_fd_sc_hd__xor2_1
XFILLER_65_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_884 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_141_clk clknet_5_25__leaf_clk VGND VGND VPWR VPWR clknet_leaf_141_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_166_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_90_0 s$1817 c$2550 c$2552 VGND VGND VPWR VPWR c$3230 s$3231 sky130_fd_sc_hd__fa_1
XFILLER_135_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_104_2 pp_row104_14 c$1950 c$1952 VGND VGND VPWR VPWR c$2674 s$2675 sky130_fd_sc_hd__fa_1
XFILLER_150_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_118_0 c$3864 c$3866 s$3869 VGND VGND VPWR VPWR c$4132 s$4133 sky130_fd_sc_hd__fa_1
XFILLER_64_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$700 t$4763 net1415 VGND VGND VPWR VPWR booth_b10_m4 sky130_fd_sc_hd__xor2_1
XFILLER_91_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$861 final_adder.p_new$892 final_adder.g_new$957 final_adder.g_new$893
+ VGND VGND VPWR VPWR final_adder.g_new$989 sky130_fd_sc_hd__a21o_2
XU$$711 net1499 net404 net1224 net670 VGND VGND VPWR VPWR t$4769 sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_38_3 s$1187 s$1189 s$1191 VGND VGND VPWR VPWR c$2148 s$2149 sky130_fd_sc_hd__fa_2
XU$$722 t$4774 net1412 VGND VGND VPWR VPWR booth_b10_m15 sky130_fd_sc_hd__xor2_1
XFILLER_90_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$883 final_adder.p_new$914 final_adder.g_new$747 final_adder.g_new$915
+ VGND VGND VPWR VPWR final_adder.g_new$1011 sky130_fd_sc_hd__a21o_1
XU$$733 net1114 net402 net1105 net668 VGND VGND VPWR VPWR t$4780 sky130_fd_sc_hd__a22o_1
XFILLER_72_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$744 t$4785 net1416 VGND VGND VPWR VPWR booth_b10_m26 sky130_fd_sc_hd__xor2_1
XU$$755 net1015 net401 net998 net667 VGND VGND VPWR VPWR t$4791 sky130_fd_sc_hd__a22o_1
XFILLER_44_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$766 t$4796 net1413 VGND VGND VPWR VPWR booth_b10_m37 sky130_fd_sc_hd__xor2_1
XFILLER_56_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_1115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$777 net1744 net405 net1736 net671 VGND VGND VPWR VPWR t$4802 sky130_fd_sc_hd__a22o_1
XU$$788 t$4807 net1419 VGND VGND VPWR VPWR booth_b10_m48 sky130_fd_sc_hd__xor2_1
XU$$799 net1630 net403 net1620 net669 VGND VGND VPWR VPWR t$4813 sky130_fd_sc_hd__a22o_1
XFILLER_25_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_132_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_132_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_185_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_5 c$4238 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1570_ clknet_leaf_19_clk booth_b36_m4 VGND VGND VPWR VPWR pp_row40_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_153_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0521_ clknet_leaf_159_clk booth_b50_m30 VGND VGND VPWR VPWR pp_row80_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0452_ clknet_leaf_158_clk booth_b32_m46 VGND VGND VPWR VPWR pp_row78_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_112_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_199_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_199_clk
+ sky130_fd_sc_hd__clkbuf_16
X_0383_ clknet_leaf_204_clk booth_b18_m58 VGND VGND VPWR VPWR pp_row76_4 sky130_fd_sc_hd__dfxtp_1
Xfanout1050 net1054 VGND VGND VPWR VPWR net1050 sky130_fd_sc_hd__buf_6
XFILLER_117_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1061 net1062 VGND VGND VPWR VPWR net1061 sky130_fd_sc_hd__buf_2
X_2122_ clknet_leaf_218_clk booth_b12_m47 VGND VGND VPWR VPWR pp_row59_6 sky130_fd_sc_hd__dfxtp_1
Xfanout1072 net1079 VGND VGND VPWR VPWR net1072 sky130_fd_sc_hd__clkbuf_4
XFILLER_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1083 net1084 VGND VGND VPWR VPWR net1083 sky130_fd_sc_hd__buf_4
Xfanout1094 net1096 VGND VGND VPWR VPWR net1094 sky130_fd_sc_hd__clkbuf_8
Xdadda_fa_2_40_3 pp_row40_20 pp_row40_21 pp_row40_22 VGND VGND VPWR VPWR c$1212 s$1213
+ sky130_fd_sc_hd__fa_1
XFILLER_54_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2053_ clknet_leaf_38_clk booth_b12_m45 VGND VGND VPWR VPWR pp_row57_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_33_2 pp_row33_6 pp_row33_7 pp_row33_8 VGND VGND VPWR VPWR c$1126 s$1127
+ sky130_fd_sc_hd__fa_1
X_1004_ clknet_leaf_117_clk booth_b48_m53 VGND VGND VPWR VPWR pp_row101_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_23_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2140 t$5498 net1446 VGND VGND VPWR VPWR booth_b30_m39 sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_10_1 c$2752 s$2755 s$2757 VGND VGND VPWR VPWR c$3438 s$3439 sky130_fd_sc_hd__fa_1
XU$$2151 net1722 net578 net1713 net851 VGND VGND VPWR VPWR t$5504 sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_26_1 pp_row26_3 pp_row26_4 pp_row26_5 VGND VGND VPWR VPWR c$1064 s$1065
+ sky130_fd_sc_hd__fa_1
XU$$2162 t$5509 net1444 VGND VGND VPWR VPWR booth_b30_m50 sky130_fd_sc_hd__xor2_1
XFILLER_179_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2173 net1613 net578 net1605 net851 VGND VGND VPWR VPWR t$5515 sky130_fd_sc_hd__a22o_1
XU$$2184 t$5520 net1446 VGND VGND VPWR VPWR booth_b30_m61 sky130_fd_sc_hd__xor2_1
XU$$2195 net1435 notblock$5525\[1\] VGND VGND VPWR VPWR t$5526 sky130_fd_sc_hd__and2_1
XU$$1450 net969 net630 net961 net903 VGND VGND VPWR VPWR t$5146 sky130_fd_sc_hd__a22o_1
XFILLER_34_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1461 t$5151 net1490 VGND VGND VPWR VPWR booth_b20_m42 sky130_fd_sc_hd__xor2_1
XFILLER_179_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1472 net1702 net634 net1692 net907 VGND VGND VPWR VPWR t$5157 sky130_fd_sc_hd__a22o_1
XU$$1483 t$5162 net1492 VGND VGND VPWR VPWR booth_b20_m53 sky130_fd_sc_hd__xor2_1
XFILLER_37_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1494 net1588 net633 net1579 net906 VGND VGND VPWR VPWR t$5168 sky130_fd_sc_hd__a22o_1
X_1906_ clknet_leaf_70_clk booth_b40_m12 VGND VGND VPWR VPWR pp_row52_20 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_123_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_123_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_31_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1837_ clknet_leaf_25_clk booth_b28_m22 VGND VGND VPWR VPWR pp_row50_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1768_ clknet_leaf_238_clk booth_b8_m40 VGND VGND VPWR VPWR pp_row48_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0719_ clknet_leaf_134_clk booth_b24_m64 VGND VGND VPWR VPWR pp_row88_1 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_85_5 pp_row85_15 pp_row85_16 pp_row85_17 VGND VGND VPWR VPWR c$976 s$977
+ sky130_fd_sc_hd__fa_1
X_1699_ clknet_leaf_23_clk booth_b34_m11 VGND VGND VPWR VPWR pp_row45_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_89_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_78_4 pp_row78_14 pp_row78_15 pp_row78_16 VGND VGND VPWR VPWR c$860 s$861
+ sky130_fd_sc_hd__fa_1
XFILLER_106_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$102 c$4354 s$4357 VGND VGND VPWR VPWR final_adder.$signal$206 final_adder.$signal$1192
+ sky130_fd_sc_hd__ha_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4511_1876 VGND VGND VPWR VPWR U$$4511_1876/HI net1876 sky130_fd_sc_hd__conb_1
XFILLER_112_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_1025 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$113 c$4376 s$4379 VGND VGND VPWR VPWR final_adder.$signal$228 final_adder.$signal$1203
+ sky130_fd_sc_hd__ha_1
XTAP_4129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_48_2 s$2225 s$2227 s$2229 VGND VGND VPWR VPWR c$2982 s$2983 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$124 c$4398 s$4401 VGND VGND VPWR VPWR final_adder.$signal$250 final_adder.$signal$1214
+ sky130_fd_sc_hd__ha_2
Xfinal_adder.U$$135 final_adder.$signal$1211 final_adder.$signal$242 final_adder.$signal$244
+ VGND VGND VPWR VPWR final_adder.g_new$263 sky130_fd_sc_hd__a21o_1
XTAP_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$146 final_adder.$signal$1198 final_adder.$signal$1199 VGND VGND VPWR
+ VPWR final_adder.p_new$274 sky130_fd_sc_hd__and2_1
XTAP_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$157 final_adder.$signal$1189 final_adder.$signal$198 final_adder.$signal$200
+ VGND VGND VPWR VPWR final_adder.g_new$285 sky130_fd_sc_hd__a21o_1
XTAP_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$168 final_adder.$signal$1176 final_adder.$signal$1177 VGND VGND VPWR
+ VPWR final_adder.p_new$296 sky130_fd_sc_hd__and2_1
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$179 final_adder.$signal$1167 final_adder.$signal$154 final_adder.$signal$156
+ VGND VGND VPWR VPWR final_adder.g_new$307 sky130_fd_sc_hd__a21o_1
XANTENNA_406 net1714 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_18_0 s$3471 c$3930 s$3933 VGND VGND VPWR VPWR c$4188 s$4189 sky130_fd_sc_hd__fa_2
XANTENNA_417 net408 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_428 net678 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_439 net949 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_114_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_114_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_16_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4479_1860 VGND VGND VPWR VPWR U$$4479_1860/HI net1860 sky130_fd_sc_hd__conb_1
XFILLER_154_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_607 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput120 b[5] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__buf_2
Xinput131 c[101] VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_50_2 c$1324 s$1327 s$1329 VGND VGND VPWR VPWR c$2242 s$2243 sky130_fd_sc_hd__fa_1
XFILLER_23_1128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput142 c[111] VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_1
Xinput153 c[121] VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_0_66_2 pp_row66_6 pp_row66_7 pp_row66_8 VGND VGND VPWR VPWR c$112 s$113
+ sky130_fd_sc_hd__fa_1
Xinput164 c[16] VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput175 c[26] VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_3_43_1 c$1234 c$1236 c$1238 VGND VGND VPWR VPWR c$2184 s$2185 sky130_fd_sc_hd__fa_1
Xinput186 c[36] VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_0_59_1 pp_row59_3 pp_row59_4 pp_row59_5 VGND VGND VPWR VPWR c$34 s$35 sky130_fd_sc_hd__fa_1
Xinput197 c[46] VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_6_20_0 c$3472 c$3474 s$3477 VGND VGND VPWR VPWR c$3936 s$3937 sky130_fd_sc_hd__fa_1
XTAP_3940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$680 final_adder.p_new$704 final_adder.p_new$688 VGND VGND VPWR VPWR
+ final_adder.p_new$808 sky130_fd_sc_hd__and2_1
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_36_0 s$211 c$1146 c$1148 VGND VGND VPWR VPWR c$2126 s$2127 sky130_fd_sc_hd__fa_1
XTAP_3962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$530 t$4675 net1246 VGND VGND VPWR VPWR booth_b6_m56 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$691 final_adder.p_new$698 final_adder.g_new$715 final_adder.g_new$699
+ VGND VGND VPWR VPWR final_adder.g_new$819 sky130_fd_sc_hd__a21o_1
XTAP_3973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$541 net1547 net432 net1539 net714 VGND VGND VPWR VPWR t$4681 sky130_fd_sc_hd__a22o_1
XTAP_3984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$552 notblock$4685\[2\] net63 net1246 t$4686 notblock$4685\[0\] VGND VGND VPWR
+ VPWR sel_0$4687 sky130_fd_sc_hd__a32o_1
XTAP_3995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$563 t$4693 net1240 VGND VGND VPWR VPWR booth_b8_m4 sky130_fd_sc_hd__xor2_1
XFILLER_60_911 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$574 net1496 net415 net1221 net681 VGND VGND VPWR VPWR t$4699 sky130_fd_sc_hd__a22o_1
XFILLER_44_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$585 t$4704 net1241 VGND VGND VPWR VPWR booth_b8_m15 sky130_fd_sc_hd__xor2_1
XU$$596 net1114 net409 net1105 net675 VGND VGND VPWR VPWR t$4710 sky130_fd_sc_hd__a22o_1
XFILLER_147_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_105_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_105_clk
+ sky130_fd_sc_hd__clkbuf_16
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_5_17__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_5_17__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_9_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1622_ clknet_leaf_5_clk booth_b38_m4 VGND VGND VPWR VPWR pp_row42_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_173_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_95_4 pp_row95_15 pp_row95_16 pp_row95_17 VGND VGND VPWR VPWR c$1874 s$1875
+ sky130_fd_sc_hd__fa_1
XFILLER_126_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1553_ clknet_leaf_5_clk booth_b4_m36 VGND VGND VPWR VPWR pp_row40_2 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_88_3 c$990 c$992 c$994 VGND VGND VPWR VPWR c$1788 s$1789 sky130_fd_sc_hd__fa_2
XFILLER_98_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0504_ clknet_leaf_157_clk booth_b18_m62 VGND VGND VPWR VPWR pp_row80_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_193_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1484_ clknet_leaf_45_clk booth_b6_m31 VGND VGND VPWR VPWR pp_row37_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_140_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_58_1 s$3039 s$3041 s$3043 VGND VGND VPWR VPWR c$3630 s$3631 sky130_fd_sc_hd__fa_1
X_0435_ clknet_leaf_153_clk booth_b54_m23 VGND VGND VPWR VPWR pp_row77_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0366_ clknet_leaf_125_clk booth_b56_m58 VGND VGND VPWR VPWR pp_row114_4 sky130_fd_sc_hd__dfxtp_1
X_2105_ clknet_leaf_137_clk booth_b50_m59 VGND VGND VPWR VPWR pp_row109_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_54_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0297_ clknet_leaf_201_clk booth_b34_m39 VGND VGND VPWR VPWR pp_row73_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_82_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2036_ clknet_leaf_72_clk booth_b44_m12 VGND VGND VPWR VPWR pp_row56_22 sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_104_1 pp_row104_3 pp_row104_4 pp_row104_5 VGND VGND VPWR VPWR c$1958 s$1959
+ sky130_fd_sc_hd__fa_1
XFILLER_35_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1280 t$5059 net1664 VGND VGND VPWR VPWR booth_b18_m20 sky130_fd_sc_hd__xor2_1
XU$$1291 net1073 net636 net1063 net909 VGND VGND VPWR VPWR t$5065 sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_125_0 pp_row125_0 pp_row125_1 pp_row125_2 VGND VGND VPWR VPWR c$3896 s$3897
+ sky130_fd_sc_hd__fa_2
XFILLER_148_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_83_2 pp_row83_6 pp_row83_7 pp_row83_8 VGND VGND VPWR VPWR c$942 s$943
+ sky130_fd_sc_hd__fa_1
XFILLER_104_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_1136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout810 net811 VGND VGND VPWR VPWR net810 sky130_fd_sc_hd__clkbuf_8
Xdadda_fa_4_60_1 c$2314 c$2316 s$2319 VGND VGND VPWR VPWR c$3052 s$3053 sky130_fd_sc_hd__fa_1
Xfanout821 net823 VGND VGND VPWR VPWR net821 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_76_1 pp_row76_8 pp_row76_9 pp_row76_10 VGND VGND VPWR VPWR c$818 s$819
+ sky130_fd_sc_hd__fa_1
Xfanout832 sel_1$5668 VGND VGND VPWR VPWR net832 sky130_fd_sc_hd__buf_4
Xfanout843 sel_1$5528 VGND VGND VPWR VPWR net843 sky130_fd_sc_hd__buf_8
Xdadda_fa_4_53_0 s$1373 c$2254 c$2256 VGND VGND VPWR VPWR c$3008 s$3009 sky130_fd_sc_hd__fa_1
XFILLER_86_830 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout854 net855 VGND VGND VPWR VPWR net854 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_69_0 pp_row69_15 pp_row69_16 pp_row69_17 VGND VGND VPWR VPWR c$690 s$691
+ sky130_fd_sc_hd__fa_2
Xfanout865 sel_1$5388 VGND VGND VPWR VPWR net865 sky130_fd_sc_hd__buf_6
Xfanout876 net877 VGND VGND VPWR VPWR net876 sky130_fd_sc_hd__clkbuf_4
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout887 net888 VGND VGND VPWR VPWR net887 sky130_fd_sc_hd__buf_2
Xfanout898 sel_1$4478 VGND VGND VPWR VPWR net898 sky130_fd_sc_hd__clkbuf_4
XTAP_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2909 net1208 net523 net1200 net796 VGND VGND VPWR VPWR t$5892 sky130_fd_sc_hd__a22o_1
XFILLER_22_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_203 net1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_214 net1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_225 net1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_236 net1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_247 net1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_258 net1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_269 net1732 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_98_2 c$1900 s$1903 s$1905 VGND VGND VPWR VPWR c$2626 s$2627 sky130_fd_sc_hd__fa_1
XFILLER_182_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_68_0 c$3664 c$3666 s$3669 VGND VGND VPWR VPWR c$4032 s$4033 sky130_fd_sc_hd__fa_1
Xdadda_fa_1_86_0_1899 VGND VGND VPWR VPWR net1899 dadda_fa_1_86_0_1899/LO sky130_fd_sc_hd__conb_1
Xdadda_fa_0_71_0 pp_row71_0 pp_row71_1 pp_row71_2 VGND VGND VPWR VPWR c$164 s$165
+ sky130_fd_sc_hd__fa_1
XFILLER_7_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0220_ clknet_leaf_199_clk booth_b16_m55 VGND VGND VPWR VPWR pp_row71_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_27_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_5_7_1 pp_row7_3 pp_row7_4 VGND VGND VPWR VPWR c$3426 s$3427 sky130_fd_sc_hd__ha_1
XTAP_3770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$360 net940 net529 net924 net802 VGND VGND VPWR VPWR t$4589 sky130_fd_sc_hd__a22o_1
XFILLER_17_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$371 t$4594 net1279 VGND VGND VPWR VPWR booth_b4_m45 sky130_fd_sc_hd__xor2_1
XU$$382 net1658 net533 net1650 net806 VGND VGND VPWR VPWR t$4600 sky130_fd_sc_hd__a22o_1
XFILLER_32_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$393 t$4605 net1276 VGND VGND VPWR VPWR booth_b4_m56 sky130_fd_sc_hd__xor2_1
XFILLER_20_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0984_ clknet_leaf_115_clk booth_b44_m56 VGND VGND VPWR VPWR pp_row100_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_164_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_559 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_93_1 pp_row93_9 pp_row93_10 pp_row93_11 VGND VGND VPWR VPWR c$1844 s$1845
+ sky130_fd_sc_hd__fa_1
XFILLER_173_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1605_ clknet_leaf_110_clk booth_b60_m45 VGND VGND VPWR VPWR pp_row105_10 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_70_0 c$3104 c$3106 c$3108 VGND VGND VPWR VPWR c$3676 s$3677 sky130_fd_sc_hd__fa_1
XFILLER_172_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_86_0 pp_row86_17 pp_row86_18 pp_row86_19 VGND VGND VPWR VPWR c$1758 s$1759
+ sky130_fd_sc_hd__fa_1
XFILLER_114_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1536_ clknet_leaf_8_clk booth_b16_m23 VGND VGND VPWR VPWR pp_row39_8 sky130_fd_sc_hd__dfxtp_1
Xdadda_ha_1_49_7 pp_row49_21 pp_row49_22 VGND VGND VPWR VPWR c$346 s$347 sky130_fd_sc_hd__ha_1
XFILLER_99_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1467_ clknet_leaf_40_clk booth_b18_m18 VGND VGND VPWR VPWR pp_row36_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_113_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_62_7 c$58 s$61 s$63 VGND VGND VPWR VPWR c$578 s$579 sky130_fd_sc_hd__fa_1
X_0418_ clknet_leaf_145_clk booth_b24_m53 VGND VGND VPWR VPWR pp_row77_6 sky130_fd_sc_hd__dfxtp_1
X_1398_ clknet_leaf_54_clk booth_b6_m27 VGND VGND VPWR VPWR pp_row33_3 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_55_6 pp_row55_23 pp_row55_24 pp_row55_25 VGND VGND VPWR VPWR c$450 s$451
+ sky130_fd_sc_hd__fa_1
X_0349_ clknet_leaf_200_clk booth_b12_m63 VGND VGND VPWR VPWR pp_row75_1 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_48_5 pp_row48_15 pp_row48_16 pp_row48_17 VGND VGND VPWR VPWR c$326 s$327
+ sky130_fd_sc_hd__fa_1
XFILLER_103_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_7_0 s$3427 c$3908 s$3911 VGND VGND VPWR VPWR c$4166 s$4167 sky130_fd_sc_hd__fa_1
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2019_ clknet_leaf_81_clk booth_b12_m44 VGND VGND VPWR VPWR pp_row56_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_85_0 s$3739 c$4064 s$4067 VGND VGND VPWR VPWR c$4322 s$4323 sky130_fd_sc_hd__fa_2
XFILLER_109_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_74_0_1894 VGND VGND VPWR VPWR net1894 dadda_fa_0_74_0_1894/LO sky130_fd_sc_hd__conb_1
XFILLER_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1605 net1606 VGND VGND VPWR VPWR net1605 sky130_fd_sc_hd__buf_4
XFILLER_78_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1616 net1619 VGND VGND VPWR VPWR net1616 sky130_fd_sc_hd__buf_4
Xfanout1627 net1628 VGND VGND VPWR VPWR net1627 sky130_fd_sc_hd__buf_4
XFILLER_120_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1086 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout640 net642 VGND VGND VPWR VPWR net640 sky130_fd_sc_hd__buf_4
Xfanout1638 net1640 VGND VGND VPWR VPWR net1638 sky130_fd_sc_hd__buf_6
Xfanout651 net652 VGND VGND VPWR VPWR net651 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1649 net111 VGND VGND VPWR VPWR net1649 sky130_fd_sc_hd__clkbuf_8
Xfanout662 net664 VGND VGND VPWR VPWR net662 sky130_fd_sc_hd__buf_4
XU$$4108 t$6503 net1284 VGND VGND VPWR VPWR booth_b58_m64 sky130_fd_sc_hd__xor2_1
XU$$4119 t$6510 net1263 VGND VGND VPWR VPWR booth_b60_m1 sky130_fd_sc_hd__xor2_1
Xfanout673 net674 VGND VGND VPWR VPWR net673 sky130_fd_sc_hd__buf_6
Xfanout684 net692 VGND VGND VPWR VPWR net684 sky130_fd_sc_hd__buf_4
XFILLER_46_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout695 sel_1$6648 VGND VGND VPWR VPWR net695 sky130_fd_sc_hd__buf_4
XFILLER_74_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3407 t$6145 net1344 VGND VGND VPWR VPWR booth_b48_m56 sky130_fd_sc_hd__xor2_1
XTAP_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3418 net1548 net495 net1540 net768 VGND VGND VPWR VPWR t$6151 sky130_fd_sc_hd__a22o_1
XTAP_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_100_0 c$3792 c$3794 s$3797 VGND VGND VPWR VPWR c$4096 s$4097 sky130_fd_sc_hd__fa_1
XU$$3429 notblock$6155\[2\] net46 net1342 t$6156 notblock$6155\[0\] VGND VGND VPWR
+ VPWR sel_0$6157 sky130_fd_sc_hd__a32o_2
XTAP_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2706 t$5787 net1396 VGND VGND VPWR VPWR booth_b38_m48 sky130_fd_sc_hd__xor2_1
XFILLER_37_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2717 net1635 net547 net1627 net820 VGND VGND VPWR VPWR t$5793 sky130_fd_sc_hd__a22o_1
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2728 t$5798 net1400 VGND VGND VPWR VPWR booth_b38_m59 sky130_fd_sc_hd__xor2_1
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2739 net1401 VGND VGND VPWR VPWR notsign$5804 sky130_fd_sc_hd__inv_1
XTAP_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2370_ clknet_leaf_127_clk booth_b54_m57 VGND VGND VPWR VPWR pp_row111_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_155_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_882 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1321_ clknet_leaf_0_clk booth_b10_m19 VGND VGND VPWR VPWR pp_row29_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_150_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_65_5 s$629 s$631 s$633 VGND VGND VPWR VPWR c$1516 s$1517 sky130_fd_sc_hd__fa_1
X_1252_ clknet_leaf_10_clk booth_b10_m15 VGND VGND VPWR VPWR pp_row25_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_77_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_58_4 s$497 s$499 s$501 VGND VGND VPWR VPWR c$1430 s$1431 sky130_fd_sc_hd__fa_1
XFILLER_83_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0203_ clknet_leaf_153_clk booth_b46_m24 VGND VGND VPWR VPWR pp_row70_21 sky130_fd_sc_hd__dfxtp_1
X_1183_ clknet_leaf_124_clk booth_b40_m63 VGND VGND VPWR VPWR pp_row103_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_76_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3930 net1734 net466 net1726 net739 VGND VGND VPWR VPWR t$6413 sky130_fd_sc_hd__a22o_1
XU$$3941 t$6418 net1298 VGND VGND VPWR VPWR booth_b56_m49 sky130_fd_sc_hd__xor2_1
XTAP_4290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3952 net1624 net465 net1616 net738 VGND VGND VPWR VPWR t$6424 sky130_fd_sc_hd__a22o_1
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3963 t$6429 net1297 VGND VGND VPWR VPWR booth_b56_m60 sky130_fd_sc_hd__xor2_1
XU$$3974 net54 VGND VGND VPWR VPWR notblock$6435\[1\] sky130_fd_sc_hd__inv_1
XU$$3985 net1034 net451 net935 net724 VGND VGND VPWR VPWR t$6442 sky130_fd_sc_hd__a22o_1
XU$$3996 t$6447 net1287 VGND VGND VPWR VPWR booth_b58_m8 sky130_fd_sc_hd__xor2_1
XFILLER_75_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$190 t$4502 net1386 VGND VGND VPWR VPWR booth_b2_m23 sky130_fd_sc_hd__xor2_1
XFILLER_178_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0967_ clknet_leaf_116_clk booth_b44_m55 VGND VGND VPWR VPWR pp_row99_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_174_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0898_ clknet_leaf_101_clk booth_b62_m33 VGND VGND VPWR VPWR pp_row95_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_127_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput265 net265 VGND VGND VPWR VPWR o[107] sky130_fd_sc_hd__buf_2
Xoutput276 net276 VGND VGND VPWR VPWR o[117] sky130_fd_sc_hd__buf_2
XFILLER_88_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput287 net287 VGND VGND VPWR VPWR o[127] sky130_fd_sc_hd__buf_2
Xoutput298 net298 VGND VGND VPWR VPWR o[21] sky130_fd_sc_hd__buf_2
X_1519_ clknet_leaf_246_clk booth_b28_m10 VGND VGND VPWR VPWR pp_row38_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_101_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2499_ clknet_leaf_97_clk booth_b38_m31 VGND VGND VPWR VPWR pp_row69_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_59_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_60_4 pp_row60_26 pp_row60_27 pp_row60_28 VGND VGND VPWR VPWR c$536 s$537
+ sky130_fd_sc_hd__fa_1
XFILLER_56_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_53_3 pp_row53_11 pp_row53_12 pp_row53_13 VGND VGND VPWR VPWR c$408 s$409
+ sky130_fd_sc_hd__fa_1
Xclkbuf_leaf_94_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_94_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_55_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_30_2 s$2081 s$2083 s$2085 VGND VGND VPWR VPWR c$2874 s$2875 sky130_fd_sc_hd__fa_1
Xdadda_fa_1_46_2 pp_row46_6 pp_row46_7 pp_row46_8 VGND VGND VPWR VPWR c$292 s$293
+ sky130_fd_sc_hd__fa_2
XFILLER_83_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_23_1 c$2018 c$2020 s$2023 VGND VGND VPWR VPWR c$2830 s$2831 sky130_fd_sc_hd__fa_1
Xdadda_fa_1_39_1 pp_row39_3 pp_row39_4 pp_row39_5 VGND VGND VPWR VPWR c$224 s$225
+ sky130_fd_sc_hd__fa_1
Xdadda_fa_4_16_0 pp_row16_5 pp_row16_6 pp_row16_7 VGND VGND VPWR VPWR c$2786 s$2787
+ sky130_fd_sc_hd__fa_1
XFILLER_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_1025 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1402 net33 VGND VGND VPWR VPWR net1402 sky130_fd_sc_hd__buf_6
Xfanout1413 net3 VGND VGND VPWR VPWR net1413 sky130_fd_sc_hd__buf_4
Xdadda_fa_3_68_3 s$1547 s$1549 s$1551 VGND VGND VPWR VPWR c$2388 s$2389 sky130_fd_sc_hd__fa_1
Xfanout1424 net1429 VGND VGND VPWR VPWR net1424 sky130_fd_sc_hd__buf_4
Xfanout1435 net1436 VGND VGND VPWR VPWR net1435 sky130_fd_sc_hd__buf_6
Xfanout1446 net1447 VGND VGND VPWR VPWR net1446 sky130_fd_sc_hd__buf_8
Xfanout1457 net1459 VGND VGND VPWR VPWR net1457 sky130_fd_sc_hd__buf_6
Xfanout1468 net18 VGND VGND VPWR VPWR net1468 sky130_fd_sc_hd__buf_6
Xfanout470 net471 VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__clkbuf_4
Xfanout481 sel_0$6227 VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__buf_4
XFILLER_120_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1479 net1480 VGND VGND VPWR VPWR net1479 sky130_fd_sc_hd__clkbuf_4
Xfanout492 sel_0$6157 VGND VGND VPWR VPWR net492 sky130_fd_sc_hd__clkbuf_8
XU$$3204 t$6042 net1354 VGND VGND VPWR VPWR booth_b46_m23 sky130_fd_sc_hd__xor2_1
XFILLER_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3215 net1051 net503 net1043 net776 VGND VGND VPWR VPWR t$6048 sky130_fd_sc_hd__a22o_1
XFILLER_46_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3226 t$6053 net1350 VGND VGND VPWR VPWR booth_b46_m34 sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_85_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_85_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_74_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3237 net942 net503 net926 net776 VGND VGND VPWR VPWR t$6059 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$19 c$4188 s$4191 VGND VGND VPWR VPWR final_adder.$signal$40 final_adder.$signal$1109
+ sky130_fd_sc_hd__ha_1
XFILLER_185_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2503 t$5684 net1406 VGND VGND VPWR VPWR booth_b36_m15 sky130_fd_sc_hd__xor2_1
XU$$3248 t$6064 net1355 VGND VGND VPWR VPWR booth_b46_m45 sky130_fd_sc_hd__xor2_1
XFILLER_47_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3259 net1660 net507 net1652 net780 VGND VGND VPWR VPWR t$6070 sky130_fd_sc_hd__a22o_1
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2514 net1118 net552 net1109 net825 VGND VGND VPWR VPWR t$5690 sky130_fd_sc_hd__a22o_1
XU$$2525 t$5695 net1405 VGND VGND VPWR VPWR booth_b36_m26 sky130_fd_sc_hd__xor2_1
XU$$2536 net1021 net557 net1004 net830 VGND VGND VPWR VPWR t$5701 sky130_fd_sc_hd__a22o_1
XU$$1802 t$5326 net1460 VGND VGND VPWR VPWR booth_b26_m7 sky130_fd_sc_hd__xor2_1
XU$$2547 t$5706 net1405 VGND VGND VPWR VPWR booth_b36_m37 sky130_fd_sc_hd__xor2_1
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1813 net1203 net594 net1194 net867 VGND VGND VPWR VPWR t$5332 sky130_fd_sc_hd__a22o_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2558 net1739 net555 net1731 net828 VGND VGND VPWR VPWR t$5712 sky130_fd_sc_hd__a22o_1
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2569 t$5717 net1408 VGND VGND VPWR VPWR booth_b36_m48 sky130_fd_sc_hd__xor2_1
XFILLER_62_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1824 t$5337 net1458 VGND VGND VPWR VPWR booth_b26_m18 sky130_fd_sc_hd__xor2_1
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1835 net1090 net596 net1084 net869 VGND VGND VPWR VPWR t$5343 sky130_fd_sc_hd__a22o_1
XU$$1846 t$5348 net1461 VGND VGND VPWR VPWR booth_b26_m29 sky130_fd_sc_hd__xor2_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1857 net982 net595 net973 net868 VGND VGND VPWR VPWR t$5354 sky130_fd_sc_hd__a22o_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1868 t$5359 net1462 VGND VGND VPWR VPWR booth_b26_m40 sky130_fd_sc_hd__xor2_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1879 net1712 net598 net1705 net871 VGND VGND VPWR VPWR t$5365 sky130_fd_sc_hd__a22o_1
XFILLER_70_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1870_ clknet_leaf_68_clk booth_b30_m21 VGND VGND VPWR VPWR pp_row51_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_175_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0821_ clknet_leaf_164_clk booth_b60_m59 VGND VGND VPWR VPWR pp_row119_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_128_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0752_ clknet_leaf_160_clk booth_b38_m51 VGND VGND VPWR VPWR pp_row89_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_116_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0683_ clknet_leaf_176_clk booth_b48_m38 VGND VGND VPWR VPWR pp_row86_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_115_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2422_ clknet_leaf_142_clk booth_b26_m41 VGND VGND VPWR VPWR pp_row67_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_143_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_70_3 c$706 s$709 s$711 VGND VGND VPWR VPWR c$1572 s$1573 sky130_fd_sc_hd__fa_1
XFILLER_124_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2353_ clknet_leaf_77_clk booth_b36_m29 VGND VGND VPWR VPWR pp_row65_18 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_63_2 c$574 c$576 c$578 VGND VGND VPWR VPWR c$1486 s$1487 sky130_fd_sc_hd__fa_2
X_1304_ clknet_leaf_1_clk booth_b14_m14 VGND VGND VPWR VPWR pp_row28_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_85_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2284_ clknet_leaf_152_clk booth_b42_m21 VGND VGND VPWR VPWR pp_row63_21 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$509 final_adder.p_new$512 final_adder.g_new$521 final_adder.g_new$513
+ VGND VGND VPWR VPWR final_adder.g_new$637 sky130_fd_sc_hd__a21o_1
XFILLER_38_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_40_1 s$2931 s$2933 s$2935 VGND VGND VPWR VPWR c$3558 s$3559 sky130_fd_sc_hd__fa_2
Xdadda_fa_2_56_1 c$442 c$444 c$446 VGND VGND VPWR VPWR c$1400 s$1401 sky130_fd_sc_hd__fa_2
X_1235_ clknet_leaf_13_clk booth_b10_m14 VGND VGND VPWR VPWR pp_row24_5 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_33_0 c$2882 c$2884 c$2886 VGND VGND VPWR VPWR c$3528 s$3529 sky130_fd_sc_hd__fa_2
Xclkbuf_leaf_76_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_76_clk sky130_fd_sc_hd__clkbuf_16
XU$$4450 net1046 sel_0$6647 net1029 net698 VGND VGND VPWR VPWR t$6679 sky130_fd_sc_hd__a22o_1
XU$$4461 t$6684 net1851 VGND VGND VPWR VPWR booth_b64_m35 sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_49_0 pp_row49_23 pp_row49_24 pp_row49_25 VGND VGND VPWR VPWR c$1314 s$1315
+ sky130_fd_sc_hd__fa_1
XU$$4472 net930 sel_0$6647 net1751 net697 VGND VGND VPWR VPWR t$6690 sky130_fd_sc_hd__a22o_1
XFILLER_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1166_ clknet_leaf_46_clk booth_b12_m7 VGND VGND VPWR VPWR pp_row19_6 sky130_fd_sc_hd__dfxtp_1
XU$$4483 t$6695 net1862 VGND VGND VPWR VPWR booth_b64_m46 sky130_fd_sc_hd__xor2_1
XU$$4494 net1653 sel_0$6647 net1645 net697 VGND VGND VPWR VPWR t$6701 sky130_fd_sc_hd__a22o_1
XU$$3760 t$6326 net1303 VGND VGND VPWR VPWR booth_b54_m27 sky130_fd_sc_hd__xor2_1
XFILLER_37_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3771 net1003 net469 net995 net742 VGND VGND VPWR VPWR t$6332 sky130_fd_sc_hd__a22o_1
XU$$3782 t$6337 net1307 VGND VGND VPWR VPWR booth_b54_m38 sky130_fd_sc_hd__xor2_1
XU$$3793 net1734 net475 net1726 net748 VGND VGND VPWR VPWR t$6343 sky130_fd_sc_hd__a22o_1
X_1097_ clknet_leaf_59_clk booth_b6_m7 VGND VGND VPWR VPWR pp_row13_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1999_ clknet_leaf_62_clk booth_b34_m21 VGND VGND VPWR VPWR pp_row55_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_165_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_78_2 s$2465 s$2467 s$2469 VGND VGND VPWR VPWR c$3162 s$3163 sky130_fd_sc_hd__fa_1
XFILLER_192_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_48_0 s$3591 c$3990 s$3993 VGND VGND VPWR VPWR c$4248 s$4249 sky130_fd_sc_hd__fa_2
XFILLER_125_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_51_0 pp_row51_0 pp_row51_1 pp_row51_2 VGND VGND VPWR VPWR c$366 s$367
+ sky130_fd_sc_hd__fa_1
XFILLER_75_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_67_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_67_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_91_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$904 net960 net398 net952 net664 VGND VGND VPWR VPWR t$4867 sky130_fd_sc_hd__a22o_1
XFILLER_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$915 t$4872 net1315 VGND VGND VPWR VPWR booth_b12_m43 sky130_fd_sc_hd__xor2_1
XU$$926 net1687 net395 net1679 net661 VGND VGND VPWR VPWR t$4878 sky130_fd_sc_hd__a22o_1
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$937 t$4883 net1318 VGND VGND VPWR VPWR booth_b12_m54 sky130_fd_sc_hd__xor2_1
XFILLER_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$948 net1581 net395 net1552 net661 VGND VGND VPWR VPWR t$4889 sky130_fd_sc_hd__a22o_1
XU$$959 net1316 VGND VGND VPWR VPWR notblock$4895\[0\] sky130_fd_sc_hd__inv_1
XFILLER_44_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1109 t$4972 net1009 VGND VGND VPWR VPWR booth_b16_m3 sky130_fd_sc_hd__xor2_1
XFILLER_188_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_911 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_80_2 c$1684 s$1687 s$1689 VGND VGND VPWR VPWR c$2482 s$2483 sky130_fd_sc_hd__fa_1
XFILLER_98_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_73_1 c$1594 c$1596 c$1598 VGND VGND VPWR VPWR c$2424 s$2425 sky130_fd_sc_hd__fa_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_50_0 c$3592 c$3594 s$3597 VGND VGND VPWR VPWR c$3996 s$3997 sky130_fd_sc_hd__fa_2
Xfanout1210 net1213 VGND VGND VPWR VPWR net1210 sky130_fd_sc_hd__buf_4
Xdadda_fa_3_66_0 s$653 c$1506 c$1508 VGND VGND VPWR VPWR c$2366 s$2367 sky130_fd_sc_hd__fa_1
Xfanout1221 net1223 VGND VGND VPWR VPWR net1221 sky130_fd_sc_hd__buf_4
Xfanout1232 net1234 VGND VGND VPWR VPWR net1232 sky130_fd_sc_hd__buf_4
Xfanout1243 net64 VGND VGND VPWR VPWR net1243 sky130_fd_sc_hd__buf_6
Xfanout1254 net1258 VGND VGND VPWR VPWR net1254 sky130_fd_sc_hd__buf_6
Xfanout1265 net1266 VGND VGND VPWR VPWR net1265 sky130_fd_sc_hd__buf_4
XFILLER_113_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1276 net1281 VGND VGND VPWR VPWR net1276 sky130_fd_sc_hd__buf_8
Xfanout1287 net1290 VGND VGND VPWR VPWR net1287 sky130_fd_sc_hd__buf_6
XU$$3001 net1592 net525 net1584 net798 VGND VGND VPWR VPWR t$5938 sky130_fd_sc_hd__a22o_1
XFILLER_8_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_58_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_58_clk sky130_fd_sc_hd__clkbuf_16
Xfanout1298 net1299 VGND VGND VPWR VPWR net1298 sky130_fd_sc_hd__buf_4
XFILLER_47_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3012 t$5943 net1374 VGND VGND VPWR VPWR booth_b42_m64 sky130_fd_sc_hd__xor2_1
X_1020_ clknet_leaf_60_clk booth_b0_m1 VGND VGND VPWR VPWR pp_row1_0 sky130_fd_sc_hd__dfxtp_1
XU$$3023 t$5950 net1358 VGND VGND VPWR VPWR booth_b44_m1 sky130_fd_sc_hd__xor2_1
XU$$3034 net1524 net514 net1516 net787 VGND VGND VPWR VPWR t$5956 sky130_fd_sc_hd__a22o_1
XU$$3045 t$5961 net1362 VGND VGND VPWR VPWR booth_b44_m12 sky130_fd_sc_hd__xor2_1
XU$$2300 net1655 net573 net1647 net846 VGND VGND VPWR VPWR t$5580 sky130_fd_sc_hd__a22o_1
XFILLER_47_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3056 net1151 net511 net1142 net784 VGND VGND VPWR VPWR t$5967 sky130_fd_sc_hd__a22o_1
XU$$2311 t$5585 net1434 VGND VGND VPWR VPWR booth_b32_m56 sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_102_1 c$2650 c$2652 s$2655 VGND VGND VPWR VPWR c$3304 s$3305 sky130_fd_sc_hd__fa_1
XFILLER_62_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2322 net1547 net575 net1539 net848 VGND VGND VPWR VPWR t$5591 sky130_fd_sc_hd__a22o_1
XU$$3067 t$5972 net1363 VGND VGND VPWR VPWR booth_b44_m23 sky130_fd_sc_hd__xor2_1
XU$$3078 net1048 net510 net1040 net783 VGND VGND VPWR VPWR t$5978 sky130_fd_sc_hd__a22o_1
XU$$2333 notblock$5595\[2\] net28 net1435 t$5596 notblock$5595\[0\] VGND VGND VPWR
+ VPWR sel_0$5597 sky130_fd_sc_hd__a32o_1
XU$$2344 t$5603 net1420 VGND VGND VPWR VPWR booth_b34_m4 sky130_fd_sc_hd__xor2_1
XU$$3089 t$5983 net1359 VGND VGND VPWR VPWR booth_b44_m34 sky130_fd_sc_hd__xor2_1
XU$$2355 net1494 net560 net1219 net833 VGND VGND VPWR VPWR t$5609 sky130_fd_sc_hd__a22o_1
XU$$1610 t$5227 net1484 VGND VGND VPWR VPWR booth_b22_m48 sky130_fd_sc_hd__xor2_1
XU$$1621 net1629 net616 net1621 net889 VGND VGND VPWR VPWR t$5233 sky130_fd_sc_hd__a22o_1
XFILLER_62_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2366 t$5614 net1421 VGND VGND VPWR VPWR booth_b34_m15 sky130_fd_sc_hd__xor2_1
XFILLER_90_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1632 t$5238 net1482 VGND VGND VPWR VPWR booth_b22_m59 sky130_fd_sc_hd__xor2_1
XU$$2377 net1118 net563 net1109 net836 VGND VGND VPWR VPWR t$5620 sky130_fd_sc_hd__a22o_1
XU$$1643 net1481 VGND VGND VPWR VPWR notsign$5244 sky130_fd_sc_hd__inv_1
XU$$2388 t$5625 net1421 VGND VGND VPWR VPWR booth_b34_m26 sky130_fd_sc_hd__xor2_1
XFILLER_90_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2399 net1018 net564 net1001 net837 VGND VGND VPWR VPWR t$5631 sky130_fd_sc_hd__a22o_1
XU$$1654 net1123 net603 net1032 net876 VGND VGND VPWR VPWR t$5251 sky130_fd_sc_hd__a22o_1
XU$$1665 t$5256 net1466 VGND VGND VPWR VPWR booth_b24_m7 sky130_fd_sc_hd__xor2_1
XFILLER_72_1135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1676 net1206 net605 net1198 net878 VGND VGND VPWR VPWR t$5262 sky130_fd_sc_hd__a22o_1
XU$$1687 t$5267 net1466 VGND VGND VPWR VPWR booth_b24_m18 sky130_fd_sc_hd__xor2_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_123_0 s$3891 c$4140 s$4143 VGND VGND VPWR VPWR c$4398 s$4399 sky130_fd_sc_hd__fa_1
X_1922_ clknet_leaf_80_clk booth_b12_m41 VGND VGND VPWR VPWR pp_row53_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_175_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1698 net1090 net604 net1082 net877 VGND VGND VPWR VPWR t$5273 sky130_fd_sc_hd__a22o_1
XFILLER_33_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1853_ clknet_leaf_232_clk net202 VGND VGND VPWR VPWR pp_row50_27 sky130_fd_sc_hd__dfxtp_2
X_0804_ clknet_leaf_94_clk booth_b48_m43 VGND VGND VPWR VPWR pp_row91_11 sky130_fd_sc_hd__dfxtp_1
X_1784_ clknet_leaf_222_clk booth_b36_m12 VGND VGND VPWR VPWR pp_row48_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_129_996 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_88_1 s$3219 s$3221 s$3223 VGND VGND VPWR VPWR c$3750 s$3751 sky130_fd_sc_hd__fa_1
X_0735_ clknet_leaf_162_clk booth_b50_m38 VGND VGND VPWR VPWR pp_row88_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_171_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0666_ clknet_leaf_131_clk booth_b60_m57 VGND VGND VPWR VPWR pp_row117_4 sky130_fd_sc_hd__dfxtp_1
X_2405_ clknet_leaf_99_clk booth_b62_m4 VGND VGND VPWR VPWR pp_row66_31 sky130_fd_sc_hd__dfxtp_1
X_0597_ clknet_leaf_188_clk booth_b36_m47 VGND VGND VPWR VPWR pp_row83_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_112_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2336_ clknet_leaf_89_clk booth_b6_m59 VGND VGND VPWR VPWR pp_row65_3 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$306 final_adder.p_new$308 final_adder.p_new$306 VGND VGND VPWR VPWR
+ final_adder.p_new$434 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$317 final_adder.p_new$316 final_adder.g_new$319 final_adder.g_new$317
+ VGND VGND VPWR VPWR final_adder.g_new$445 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$328 final_adder.p_new$330 final_adder.p_new$328 VGND VGND VPWR VPWR
+ final_adder.p_new$456 sky130_fd_sc_hd__and2_1
XFILLER_57_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2267_ clknet_leaf_214_clk booth_b14_m49 VGND VGND VPWR VPWR pp_row63_7 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$339 final_adder.p_new$338 final_adder.g_new$341 final_adder.g_new$339
+ VGND VGND VPWR VPWR final_adder.g_new$467 sky130_fd_sc_hd__a21o_1
XFILLER_73_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_49_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_49_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_38_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1218_ clknet_leaf_48_clk booth_b4_m19 VGND VGND VPWR VPWR pp_row23_2 sky130_fd_sc_hd__dfxtp_1
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4280 t$6592 net1254 VGND VGND VPWR VPWR booth_b62_m13 sky130_fd_sc_hd__xor2_1
X_2198_ clknet_leaf_228_clk booth_b20_m41 VGND VGND VPWR VPWR pp_row61_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_81_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4291 net1141 net418 net1135 net700 VGND VGND VPWR VPWR t$6598 sky130_fd_sc_hd__a22o_1
XFILLER_77_1035 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1149_ clknet_leaf_119_clk booth_b64_m38 VGND VGND VPWR VPWR pp_row102_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_81_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3590 net1222 net476 net1215 net749 VGND VGND VPWR VPWR t$6240 sky130_fd_sc_hd__a22o_1
XFILLER_179_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_90_1 c$2554 c$2556 s$2559 VGND VGND VPWR VPWR c$3232 s$3233 sky130_fd_sc_hd__fa_1
XFILLER_193_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_83_0 s$1733 c$2494 c$2496 VGND VGND VPWR VPWR c$3188 s$3189 sky130_fd_sc_hd__fa_1
Xdadda_fa_3_104_3 c$1954 s$1957 s$1959 VGND VGND VPWR VPWR c$2676 s$2677 sky130_fd_sc_hd__fa_1
XFILLER_101_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_124_0_1914 VGND VGND VPWR VPWR net1914 dadda_fa_5_124_0_1914/LO sky130_fd_sc_hd__conb_1
XFILLER_88_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$851 final_adder.p_new$882 final_adder.g_new$947 final_adder.g_new$883
+ VGND VGND VPWR VPWR final_adder.g_new$979 sky130_fd_sc_hd__a21o_2
XU$$701 net1672 net406 net1561 net672 VGND VGND VPWR VPWR t$4764 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$873 final_adder.p_new$904 final_adder.g_new$857 final_adder.g_new$905
+ VGND VGND VPWR VPWR final_adder.g_new$1001 sky130_fd_sc_hd__a21o_1
XU$$712 t$4769 net1414 VGND VGND VPWR VPWR booth_b10_m10 sky130_fd_sc_hd__xor2_1
XU$$723 net1164 net401 net1155 net667 VGND VGND VPWR VPWR t$4775 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$895 final_adder.p_new$926 final_adder.g_new$509 final_adder.g_new$927
+ VGND VGND VPWR VPWR final_adder.g_new$1023 sky130_fd_sc_hd__a21o_1
XU$$734 t$4780 net1412 VGND VGND VPWR VPWR booth_b10_m21 sky130_fd_sc_hd__xor2_1
XU$$745 net1066 net406 net1057 net672 VGND VGND VPWR VPWR t$4786 sky130_fd_sc_hd__a22o_1
XU$$756 t$4791 net1413 VGND VGND VPWR VPWR booth_b10_m32 sky130_fd_sc_hd__xor2_1
XFILLER_182_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$767 net956 net401 net948 net667 VGND VGND VPWR VPWR t$4797 sky130_fd_sc_hd__a22o_1
XFILLER_56_1119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$778 t$4802 net1416 VGND VGND VPWR VPWR booth_b10_m43 sky130_fd_sc_hd__xor2_1
XFILLER_182_1127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$789 net1689 net408 net1679 net674 VGND VGND VPWR VPWR t$4808 sky130_fd_sc_hd__a22o_1
XFILLER_72_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_98_0 c$3784 c$3786 s$3789 VGND VGND VPWR VPWR c$4092 s$4093 sky130_fd_sc_hd__fa_1
XFILLER_61_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_911 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_6 c$4240 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0520_ clknet_leaf_166_clk booth_b48_m32 VGND VGND VPWR VPWR pp_row80_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_152_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0451_ clknet_leaf_158_clk booth_b30_m48 VGND VGND VPWR VPWR pp_row78_9 sky130_fd_sc_hd__dfxtp_1
X_0382_ clknet_leaf_204_clk booth_b16_m60 VGND VGND VPWR VPWR pp_row76_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_117_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1040 net1046 VGND VGND VPWR VPWR net1040 sky130_fd_sc_hd__buf_6
XFILLER_67_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1051 net1053 VGND VGND VPWR VPWR net1051 sky130_fd_sc_hd__buf_4
XFILLER_0_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2121_ clknet_leaf_218_clk booth_b10_m49 VGND VGND VPWR VPWR pp_row59_5 sky130_fd_sc_hd__dfxtp_1
Xfanout1062 net84 VGND VGND VPWR VPWR net1062 sky130_fd_sc_hd__buf_6
XFILLER_39_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1073 net1079 VGND VGND VPWR VPWR net1073 sky130_fd_sc_hd__buf_4
Xfanout1084 net81 VGND VGND VPWR VPWR net1084 sky130_fd_sc_hd__clkbuf_8
Xfanout1095 net1096 VGND VGND VPWR VPWR net1095 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_40_4 c$222 c$224 c$226 VGND VGND VPWR VPWR c$1214 s$1215 sky130_fd_sc_hd__fa_1
X_2052_ clknet_leaf_38_clk booth_b10_m47 VGND VGND VPWR VPWR pp_row57_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_35_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1003_ clknet_leaf_118_clk booth_b46_m55 VGND VGND VPWR VPWR pp_row101_5 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_33_3 pp_row33_9 pp_row33_10 pp_row33_11 VGND VGND VPWR VPWR c$1128 s$1129
+ sky130_fd_sc_hd__fa_1
XU$$2130 t$5493 net1442 VGND VGND VPWR VPWR booth_b30_m34 sky130_fd_sc_hd__xor2_1
XFILLER_34_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2141 net946 net582 net930 net855 VGND VGND VPWR VPWR t$5499 sky130_fd_sc_hd__a22o_1
XU$$2152 t$5504 net1445 VGND VGND VPWR VPWR booth_b30_m45 sky130_fd_sc_hd__xor2_1
XU$$2163 net1655 net579 net1647 net852 VGND VGND VPWR VPWR t$5510 sky130_fd_sc_hd__a22o_1
XU$$2174 t$5515 net1444 VGND VGND VPWR VPWR booth_b30_m56 sky130_fd_sc_hd__xor2_1
XFILLER_62_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1440 net1017 net629 net1000 net902 VGND VGND VPWR VPWR t$5141 sky130_fd_sc_hd__a22o_1
XFILLER_23_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2185 net1548 net582 net1540 net855 VGND VGND VPWR VPWR t$5521 sky130_fd_sc_hd__a22o_1
XU$$1451 t$5146 net1489 VGND VGND VPWR VPWR booth_b20_m37 sky130_fd_sc_hd__xor2_1
XU$$2196 notblock$5525\[2\] net26 net1444 t$5526 notblock$5525\[0\] VGND VGND VPWR
+ VPWR sel_0$5527 sky130_fd_sc_hd__a32o_4
XU$$1462 net1738 net632 net1730 net905 VGND VGND VPWR VPWR t$5152 sky130_fd_sc_hd__a22o_1
XFILLER_76_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1473 t$5157 net1493 VGND VGND VPWR VPWR booth_b20_m48 sky130_fd_sc_hd__xor2_1
XU$$1484 net1629 net632 net1620 net905 VGND VGND VPWR VPWR t$5163 sky130_fd_sc_hd__a22o_1
XFILLER_50_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1495 t$5168 net1491 VGND VGND VPWR VPWR booth_b20_m59 sky130_fd_sc_hd__xor2_1
XFILLER_188_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1905_ clknet_leaf_138_clk booth_b62_m45 VGND VGND VPWR VPWR pp_row107_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_30_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1836_ clknet_leaf_25_clk booth_b26_m24 VGND VGND VPWR VPWR pp_row50_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_135_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1767_ clknet_leaf_237_clk booth_b6_m42 VGND VGND VPWR VPWR pp_row48_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0718_ clknet_leaf_184_clk net242 VGND VGND VPWR VPWR pp_row87_22 sky130_fd_sc_hd__dfxtp_1
XFILLER_117_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1698_ clknet_leaf_19_clk booth_b32_m13 VGND VGND VPWR VPWR pp_row45_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_89_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0649_ clknet_leaf_165_clk booth_b32_m53 VGND VGND VPWR VPWR pp_row85_6 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_78_5 pp_row78_17 pp_row78_18 pp_row78_19 VGND VGND VPWR VPWR c$862 s$863
+ sky130_fd_sc_hd__fa_1
XFILLER_83_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$103 c$4356 s$4359 VGND VGND VPWR VPWR final_adder.$signal$208 final_adder.$signal$1193
+ sky130_fd_sc_hd__ha_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$114 c$4378 s$4381 VGND VGND VPWR VPWR final_adder.$signal$230 final_adder.$signal$1204
+ sky130_fd_sc_hd__ha_1
X_2319_ clknet_leaf_77_clk booth_b40_m24 VGND VGND VPWR VPWR pp_row64_20 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$125 c$4400 s$4403 VGND VGND VPWR VPWR final_adder.$signal$252 final_adder.$signal$1215
+ sky130_fd_sc_hd__ha_2
XFILLER_131_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$136 final_adder.$signal$1208 final_adder.$signal$1209 VGND VGND VPWR
+ VPWR final_adder.p_new$264 sky130_fd_sc_hd__and2_1
XTAP_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$147 final_adder.$signal$1199 final_adder.$signal$218 final_adder.$signal$220
+ VGND VGND VPWR VPWR final_adder.g_new$275 sky130_fd_sc_hd__a21o_1
XFILLER_79_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$158 final_adder.$signal$1186 final_adder.$signal$1187 VGND VGND VPWR
+ VPWR final_adder.p_new$286 sky130_fd_sc_hd__and2_1
XTAP_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$169 final_adder.$signal$1177 final_adder.$signal$174 final_adder.$signal$176
+ VGND VGND VPWR VPWR final_adder.g_new$297 sky130_fd_sc_hd__a21o_1
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_407 net1714 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_418 net455 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_429 net681 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_118_0_1912 VGND VGND VPWR VPWR net1912 dadda_fa_4_118_0_1912/LO sky130_fd_sc_hd__conb_1
Xdadda_fa_3_102_0 pp_row102_11 pp_row102_12 pp_row102_13 VGND VGND VPWR VPWR c$2654
+ s$2655 sky130_fd_sc_hd__fa_1
XFILLER_162_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_861 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput110 b[50] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__buf_6
Xinput121 b[60] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput132 c[102] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_1
Xinput143 c[112] VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_747 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_50_3 s$1331 s$1333 s$1335 VGND VGND VPWR VPWR c$2244 s$2245 sky130_fd_sc_hd__fa_1
XFILLER_88_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput154 c[122] VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_0_66_3 pp_row66_9 pp_row66_10 pp_row66_11 VGND VGND VPWR VPWR c$114 s$115
+ sky130_fd_sc_hd__fa_1
Xinput165 c[17] VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__clkbuf_1
Xinput176 c[27] VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_3_43_2 c$1240 s$1243 s$1245 VGND VGND VPWR VPWR c$2186 s$2187 sky130_fd_sc_hd__fa_1
XFILLER_76_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput187 c[37] VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_1
Xinput198 c[47] VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_0_59_2 pp_row59_6 pp_row59_7 pp_row59_8 VGND VGND VPWR VPWR c$36 s$37 sky130_fd_sc_hd__fa_1
XTAP_3930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$670 final_adder.p_new$694 final_adder.p_new$678 VGND VGND VPWR VPWR
+ final_adder.p_new$798 sky130_fd_sc_hd__and2_1
XTAP_3952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$681 final_adder.p_new$688 final_adder.g_new$705 final_adder.g_new$689
+ VGND VGND VPWR VPWR final_adder.g_new$809 sky130_fd_sc_hd__a21o_1
Xdadda_fa_3_36_1 c$1150 c$1152 c$1154 VGND VGND VPWR VPWR c$2128 s$2129 sky130_fd_sc_hd__fa_1
XU$$520 t$4670 net1251 VGND VGND VPWR VPWR booth_b6_m51 sky130_fd_sc_hd__xor2_1
XTAP_3963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$531 net1604 net433 net1595 net715 VGND VGND VPWR VPWR t$4676 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$692 final_adder.p_new$716 final_adder.p_new$700 VGND VGND VPWR VPWR
+ final_adder.p_new$820 sky130_fd_sc_hd__and2_1
XTAP_3974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$542 t$4681 net1251 VGND VGND VPWR VPWR booth_b6_m62 sky130_fd_sc_hd__xor2_1
Xdadda_fa_6_13_0 c$3444 c$3446 s$3449 VGND VGND VPWR VPWR c$3922 s$3923 sky130_fd_sc_hd__fa_1
XFILLER_186_1060 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$553 net63 net1247 VGND VGND VPWR VPWR sel_1$4688 sky130_fd_sc_hd__xor2_1
XTAP_3996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_29_0 pp_row29_11 pp_row29_12 pp_row29_13 VGND VGND VPWR VPWR c$2070 s$2071
+ sky130_fd_sc_hd__fa_1
XU$$564 net1676 net414 net1564 net680 VGND VGND VPWR VPWR t$4694 sky130_fd_sc_hd__a22o_1
XU$$575 t$4699 net1241 VGND VGND VPWR VPWR booth_b8_m10 sky130_fd_sc_hd__xor2_1
XFILLER_60_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$586 net1166 net409 net1157 net675 VGND VGND VPWR VPWR t$4705 sky130_fd_sc_hd__a22o_1
XU$$597 t$4710 net1235 VGND VGND VPWR VPWR booth_b8_m21 sky130_fd_sc_hd__xor2_1
XFILLER_60_967 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1621_ clknet_leaf_5_clk booth_b36_m6 VGND VGND VPWR VPWR pp_row42_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_184_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_95_5 pp_row95_18 c$1042 c$1044 VGND VGND VPWR VPWR c$1876 s$1877 sky130_fd_sc_hd__fa_1
XFILLER_193_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1552_ clknet_leaf_5_clk booth_b2_m38 VGND VGND VPWR VPWR pp_row40_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_114_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_88_4 c$996 c$998 s$1001 VGND VGND VPWR VPWR c$1790 s$1791 sky130_fd_sc_hd__fa_1
XFILLER_193_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0503_ clknet_leaf_206_clk booth_b16_m64 VGND VGND VPWR VPWR pp_row80_1 sky130_fd_sc_hd__dfxtp_1
X_1483_ clknet_leaf_184_clk net134 VGND VGND VPWR VPWR pp_row104_14 sky130_fd_sc_hd__dfxtp_2
XFILLER_87_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0434_ clknet_leaf_154_clk booth_b52_m25 VGND VGND VPWR VPWR pp_row77_20 sky130_fd_sc_hd__dfxtp_1
XFILLER_39_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0365_ clknet_leaf_204_clk booth_b42_m33 VGND VGND VPWR VPWR pp_row75_16 sky130_fd_sc_hd__dfxtp_1
Xdadda_ha_2_25_1 pp_row25_3 pp_row25_4 VGND VGND VPWR VPWR c$1060 s$1061 sky130_fd_sc_hd__ha_1
XFILLER_67_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2104_ clknet_leaf_30_clk booth_b44_m14 VGND VGND VPWR VPWR pp_row58_22 sky130_fd_sc_hd__dfxtp_1
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0296_ clknet_leaf_201_clk booth_b32_m41 VGND VGND VPWR VPWR pp_row73_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_54_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2035_ clknet_leaf_73_clk booth_b42_m14 VGND VGND VPWR VPWR pp_row56_21 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_31_0 pp_row31_0 pp_row31_1 pp_row31_2 VGND VGND VPWR VPWR c$1100 s$1101
+ sky130_fd_sc_hd__fa_1
XFILLER_35_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1270 t$5054 net1665 VGND VGND VPWR VPWR booth_b18_m15 sky130_fd_sc_hd__xor2_1
XU$$1281 net1115 net635 net1106 net908 VGND VGND VPWR VPWR t$5060 sky130_fd_sc_hd__a22o_1
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1292 t$5065 net1663 VGND VGND VPWR VPWR booth_b18_m26 sky130_fd_sc_hd__xor2_1
XFILLER_10_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_118_0 c$3392 c$3394 c$3396 VGND VGND VPWR VPWR c$3868 s$3869 sky130_fd_sc_hd__fa_1
XFILLER_136_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1819_ clknet_leaf_220_clk booth_b46_m3 VGND VGND VPWR VPWR pp_row49_23 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_83_3 pp_row83_9 pp_row83_10 pp_row83_11 VGND VGND VPWR VPWR c$944 s$945
+ sky130_fd_sc_hd__fa_1
XFILLER_117_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout800 net803 VGND VGND VPWR VPWR net800 sky130_fd_sc_hd__buf_4
Xfanout811 net815 VGND VGND VPWR VPWR net811 sky130_fd_sc_hd__buf_4
Xdadda_fa_4_60_2 s$2321 s$2323 s$2325 VGND VGND VPWR VPWR c$3054 s$3055 sky130_fd_sc_hd__fa_1
XFILLER_120_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout822 net823 VGND VGND VPWR VPWR net822 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_76_2 pp_row76_11 pp_row76_12 pp_row76_13 VGND VGND VPWR VPWR c$820 s$821
+ sky130_fd_sc_hd__fa_1
Xfanout833 net835 VGND VGND VPWR VPWR net833 sky130_fd_sc_hd__buf_4
Xfanout844 net845 VGND VGND VPWR VPWR net844 sky130_fd_sc_hd__buf_4
Xdadda_fa_4_53_1 c$2258 c$2260 s$2263 VGND VGND VPWR VPWR c$3010 s$3011 sky130_fd_sc_hd__fa_1
Xfanout855 net856 VGND VGND VPWR VPWR net855 sky130_fd_sc_hd__buf_6
Xfanout866 net868 VGND VGND VPWR VPWR net866 sky130_fd_sc_hd__buf_4
XFILLER_98_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_69_1 pp_row69_18 pp_row69_19 pp_row69_20 VGND VGND VPWR VPWR c$692 s$693
+ sky130_fd_sc_hd__fa_1
XFILLER_133_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout877 sel_1$5248 VGND VGND VPWR VPWR net877 sky130_fd_sc_hd__buf_4
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_30_0 s$3519 c$3954 s$3957 VGND VGND VPWR VPWR c$4212 s$4213 sky130_fd_sc_hd__fa_2
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout888 sel_1$5178 VGND VGND VPWR VPWR net888 sky130_fd_sc_hd__buf_4
Xdadda_fa_4_46_0 s$1289 c$2198 c$2200 VGND VGND VPWR VPWR c$2966 s$2967 sky130_fd_sc_hd__fa_1
Xfanout899 sel_1$4478 VGND VGND VPWR VPWR net899 sky130_fd_sc_hd__buf_4
XTAP_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_204 net1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_23__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_5_23__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA_215 net1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_226 net1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_237 net1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_248 net1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_259 net1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_98_3 s$1907 s$1909 s$1911 VGND VGND VPWR VPWR c$2628 s$2629 sky130_fd_sc_hd__fa_1
Xdadda_ha_0_72_3 pp_row72_9 pp_row72_10 VGND VGND VPWR VPWR c$178 s$179 sky130_fd_sc_hd__ha_1
XFILLER_182_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_0_71_1 pp_row71_3 pp_row71_4 pp_row71_5 VGND VGND VPWR VPWR c$166 s$167
+ sky130_fd_sc_hd__fa_1
XFILLER_89_691 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_0_64_0 pp_row64_0 pp_row64_1 pp_row64_2 VGND VGND VPWR VPWR c$84 s$85 sky130_fd_sc_hd__fa_2
XFILLER_3_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_834 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$350 net986 net532 net974 net805 VGND VGND VPWR VPWR t$4584 sky130_fd_sc_hd__a22o_1
XTAP_3782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_997 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$361 t$4589 net1276 VGND VGND VPWR VPWR booth_b4_m40 sky130_fd_sc_hd__xor2_1
XU$$372 net1711 net529 net1703 net802 VGND VGND VPWR VPWR t$4595 sky130_fd_sc_hd__a22o_1
XU$$383 t$4600 net1280 VGND VGND VPWR VPWR booth_b4_m51 sky130_fd_sc_hd__xor2_1
XU$$394 net1604 net529 net1595 net802 VGND VGND VPWR VPWR t$4606 sky130_fd_sc_hd__a22o_1
XFILLER_17_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0983_ clknet_leaf_118_clk booth_b42_m58 VGND VGND VPWR VPWR pp_row100_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_1047 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_93_2 pp_row93_12 pp_row93_13 pp_row93_14 VGND VGND VPWR VPWR c$1846 s$1847
+ sky130_fd_sc_hd__fa_1
XFILLER_172_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1604_ clknet_leaf_240_clk booth_b8_m34 VGND VGND VPWR VPWR pp_row42_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_160_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_70_1 s$3111 s$3113 s$3115 VGND VGND VPWR VPWR c$3678 s$3679 sky130_fd_sc_hd__fa_1
Xdadda_fa_2_86_1 pp_row86_20 pp_row86_21 pp_row86_22 VGND VGND VPWR VPWR c$1760 s$1761
+ sky130_fd_sc_hd__fa_1
XFILLER_99_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1535_ clknet_leaf_16_clk booth_b14_m25 VGND VGND VPWR VPWR pp_row39_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_113_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_63_0 c$3062 c$3064 c$3066 VGND VGND VPWR VPWR c$3648 s$3649 sky130_fd_sc_hd__fa_1
XFILLER_102_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_79_0 c$202 c$852 c$854 VGND VGND VPWR VPWR c$1674 s$1675 sky130_fd_sc_hd__fa_1
XFILLER_87_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1466_ clknet_leaf_40_clk booth_b16_m20 VGND VGND VPWR VPWR pp_row36_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_68_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4389_1814 VGND VGND VPWR VPWR U$$4389_1814/HI net1814 sky130_fd_sc_hd__conb_1
Xdadda_fa_1_62_8 s$65 s$67 s$69 VGND VGND VPWR VPWR c$580 s$581 sky130_fd_sc_hd__fa_2
X_0417_ clknet_leaf_155_clk booth_b22_m55 VGND VGND VPWR VPWR pp_row77_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1397_ clknet_leaf_54_clk booth_b4_m29 VGND VGND VPWR VPWR pp_row33_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_28_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_55_7 pp_row55_26 pp_row55_27 pp_row55_28 VGND VGND VPWR VPWR c$452 s$453
+ sky130_fd_sc_hd__fa_1
XFILLER_80_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0348_ clknet_leaf_203_clk notsign$4824 VGND VGND VPWR VPWR pp_row75_0 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_48_6 pp_row48_18 pp_row48_19 pp_row48_20 VGND VGND VPWR VPWR c$328 s$329
+ sky130_fd_sc_hd__fa_1
X_0279_ clknet_leaf_201_clk booth_b60_m12 VGND VGND VPWR VPWR pp_row72_27 sky130_fd_sc_hd__dfxtp_1
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2018_ clknet_leaf_81_clk booth_b10_m46 VGND VGND VPWR VPWR pp_row56_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_169_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_78_0 s$3711 c$4050 s$4053 VGND VGND VPWR VPWR c$4308 s$4309 sky130_fd_sc_hd__fa_2
XFILLER_191_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_81_0 pp_row81_0 pp_row81_1 pp_row81_2 VGND VGND VPWR VPWR c$906 s$907
+ sky130_fd_sc_hd__fa_1
XFILLER_144_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1606 net116 VGND VGND VPWR VPWR net1606 sky130_fd_sc_hd__buf_6
XFILLER_137_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1617 net1619 VGND VGND VPWR VPWR net1617 sky130_fd_sc_hd__clkbuf_2
Xfanout630 net631 VGND VGND VPWR VPWR net630 sky130_fd_sc_hd__buf_6
Xfanout1628 net114 VGND VGND VPWR VPWR net1628 sky130_fd_sc_hd__buf_4
XFILLER_104_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout641 net642 VGND VGND VPWR VPWR net641 sky130_fd_sc_hd__clkbuf_4
Xfanout1639 net1640 VGND VGND VPWR VPWR net1639 sky130_fd_sc_hd__buf_6
XFILLER_120_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout652 net658 VGND VGND VPWR VPWR net652 sky130_fd_sc_hd__buf_4
XFILLER_59_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4109 net1284 VGND VGND VPWR VPWR notsign$6504 sky130_fd_sc_hd__inv_1
Xfanout663 net664 VGND VGND VPWR VPWR net663 sky130_fd_sc_hd__buf_4
Xfanout674 sel_1$4758 VGND VGND VPWR VPWR net674 sky130_fd_sc_hd__buf_6
Xfanout685 net692 VGND VGND VPWR VPWR net685 sky130_fd_sc_hd__buf_2
Xfanout696 net699 VGND VGND VPWR VPWR net696 sky130_fd_sc_hd__buf_4
XTAP_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3408 net1609 net499 net1603 net772 VGND VGND VPWR VPWR t$6146 sky130_fd_sc_hd__a22o_1
XFILLER_46_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3419 t$6151 net1340 VGND VGND VPWR VPWR booth_b48_m62 sky130_fd_sc_hd__xor2_1
XTAP_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2707 net1688 net545 net1680 net818 VGND VGND VPWR VPWR t$5788 sky130_fd_sc_hd__a22o_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2718 t$5793 net1400 VGND VGND VPWR VPWR booth_b38_m54 sky130_fd_sc_hd__xor2_1
XFILLER_46_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2729 net1584 net547 net1557 net820 VGND VGND VPWR VPWR t$5799 sky130_fd_sc_hd__a22o_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_80_0 c$3712 c$3714 s$3717 VGND VGND VPWR VPWR c$4056 s$4057 sky130_fd_sc_hd__fa_1
Xdadda_fa_3_96_0 s$1049 c$1866 c$1868 VGND VGND VPWR VPWR c$2606 s$2607 sky130_fd_sc_hd__fa_1
XFILLER_185_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_244_clk clknet_5_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_244_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_64_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1320_ clknet_leaf_250_clk booth_b8_m21 VGND VGND VPWR VPWR pp_row29_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_151_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1251_ clknet_leaf_10_clk booth_b8_m17 VGND VGND VPWR VPWR pp_row25_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_68_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_58_5 s$503 s$505 s$507 VGND VGND VPWR VPWR c$1432 s$1433 sky130_fd_sc_hd__fa_1
XFILLER_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0202_ clknet_leaf_152_clk booth_b44_m26 VGND VGND VPWR VPWR pp_row70_20 sky130_fd_sc_hd__dfxtp_1
X_1182_ clknet_leaf_53_clk booth_b18_m2 VGND VGND VPWR VPWR pp_row20_9 sky130_fd_sc_hd__dfxtp_1
XU$$3920 net953 net464 net947 net737 VGND VGND VPWR VPWR t$6408 sky130_fd_sc_hd__a22o_1
XFILLER_76_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3931 t$6413 net1298 VGND VGND VPWR VPWR booth_b56_m44 sky130_fd_sc_hd__xor2_1
XU$$3942 net1684 net465 net1660 net738 VGND VGND VPWR VPWR t$6419 sky130_fd_sc_hd__a22o_1
XTAP_4291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3953 t$6424 net1297 VGND VGND VPWR VPWR booth_b56_m55 sky130_fd_sc_hd__xor2_1
XU$$3964 net1554 net463 net1545 net736 VGND VGND VPWR VPWR t$6430 sky130_fd_sc_hd__a22o_1
XU$$3975 net1284 VGND VGND VPWR VPWR notblock$6435\[2\] sky130_fd_sc_hd__inv_1
XFILLER_18_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3986 t$6442 net1282 VGND VGND VPWR VPWR booth_b58_m3 sky130_fd_sc_hd__xor2_1
XU$$3997 net1510 net455 net1501 net728 VGND VGND VPWR VPWR t$6448 sky130_fd_sc_hd__a22o_1
XU$$180 t$4497 net1389 VGND VGND VPWR VPWR booth_b2_m18 sky130_fd_sc_hd__xor2_1
XU$$191 net1088 net619 net1080 net892 VGND VGND VPWR VPWR t$4503 sky130_fd_sc_hd__a22o_1
XFILLER_162_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0966_ clknet_leaf_180_clk booth_b62_m59 VGND VGND VPWR VPWR pp_row121_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_118_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0897_ clknet_leaf_101_clk booth_b60_m35 VGND VGND VPWR VPWR pp_row95_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput266 net266 VGND VGND VPWR VPWR o[108] sky130_fd_sc_hd__buf_2
XFILLER_0_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_235_clk clknet_5_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_235_clk
+ sky130_fd_sc_hd__clkbuf_16
Xoutput277 net277 VGND VGND VPWR VPWR o[118] sky130_fd_sc_hd__buf_2
Xoutput288 net288 VGND VGND VPWR VPWR o[12] sky130_fd_sc_hd__buf_2
XFILLER_87_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput299 net299 VGND VGND VPWR VPWR o[22] sky130_fd_sc_hd__buf_2
X_1518_ clknet_leaf_17_clk booth_b26_m12 VGND VGND VPWR VPWR pp_row38_13 sky130_fd_sc_hd__dfxtp_1
X_2498_ clknet_leaf_97_clk booth_b36_m33 VGND VGND VPWR VPWR pp_row69_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_141_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_60_5 pp_row60_29 pp_row60_30 pp_row60_31 VGND VGND VPWR VPWR c$538 s$539
+ sky130_fd_sc_hd__fa_1
X_1449_ clknet_leaf_65_clk booth_b24_m11 VGND VGND VPWR VPWR pp_row35_12 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_53_4 pp_row53_14 pp_row53_15 pp_row53_16 VGND VGND VPWR VPWR c$410 s$411
+ sky130_fd_sc_hd__fa_1
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_46_3 pp_row46_9 pp_row46_10 pp_row46_11 VGND VGND VPWR VPWR c$294 s$295
+ sky130_fd_sc_hd__fa_1
Xdadda_fa_4_23_2 s$2025 s$2027 s$2029 VGND VGND VPWR VPWR c$2832 s$2833 sky130_fd_sc_hd__fa_1
XFILLER_71_848 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_16_1 pp_row16_8 pp_row16_9 pp_row16_10 VGND VGND VPWR VPWR c$2788 s$2789
+ sky130_fd_sc_hd__fa_1
XFILLER_130_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_226_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_226_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_105_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1403 net1405 VGND VGND VPWR VPWR net1403 sky130_fd_sc_hd__buf_6
Xfanout1414 net1415 VGND VGND VPWR VPWR net1414 sky130_fd_sc_hd__clkbuf_8
Xfanout1425 net1427 VGND VGND VPWR VPWR net1425 sky130_fd_sc_hd__buf_6
XFILLER_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1436 net1437 VGND VGND VPWR VPWR net1436 sky130_fd_sc_hd__buf_4
XFILLER_94_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1447 net25 VGND VGND VPWR VPWR net1447 sky130_fd_sc_hd__buf_8
XFILLER_47_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1458 net1459 VGND VGND VPWR VPWR net1458 sky130_fd_sc_hd__clkbuf_4
Xfanout460 net461 VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__buf_4
Xfanout471 sel_0$6297 VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__clkbuf_4
Xfanout1469 net1470 VGND VGND VPWR VPWR net1469 sky130_fd_sc_hd__buf_6
Xfanout482 net483 VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__buf_4
XFILLER_4_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout493 net496 VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__buf_4
XU$$3205 net1094 net504 net1086 net777 VGND VGND VPWR VPWR t$6043 sky130_fd_sc_hd__a22o_1
XFILLER_93_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_791 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3216 t$6048 net1351 VGND VGND VPWR VPWR booth_b46_m29 sky130_fd_sc_hd__xor2_1
XFILLER_46_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3227 net985 net503 net976 net776 VGND VGND VPWR VPWR t$6054 sky130_fd_sc_hd__a22o_1
XFILLER_19_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3238 t$6059 net1351 VGND VGND VPWR VPWR booth_b46_m40 sky130_fd_sc_hd__xor2_1
XU$$2504 net1171 net554 net1162 net827 VGND VGND VPWR VPWR t$5685 sky130_fd_sc_hd__a22o_1
XU$$3249 net1717 net507 net1708 net780 VGND VGND VPWR VPWR t$6065 sky130_fd_sc_hd__a22o_1
XFILLER_74_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2515 t$5690 net1404 VGND VGND VPWR VPWR booth_b36_m21 sky130_fd_sc_hd__xor2_1
XFILLER_73_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2526 net1068 net553 net1060 net826 VGND VGND VPWR VPWR t$5696 sky130_fd_sc_hd__a22o_1
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2537 t$5701 net1410 VGND VGND VPWR VPWR booth_b36_m32 sky130_fd_sc_hd__xor2_1
XU$$1803 net1516 net596 net1509 net869 VGND VGND VPWR VPWR t$5327 sky130_fd_sc_hd__a22o_1
XU$$2548 net957 net553 net949 net826 VGND VGND VPWR VPWR t$5707 sky130_fd_sc_hd__a22o_1
XFILLER_61_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1814 t$5332 net1457 VGND VGND VPWR VPWR booth_b26_m13 sky130_fd_sc_hd__xor2_1
XU$$2559 t$5712 net1409 VGND VGND VPWR VPWR booth_b36_m43 sky130_fd_sc_hd__xor2_1
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1825 net1139 net593 net1132 net866 VGND VGND VPWR VPWR t$5338 sky130_fd_sc_hd__a22o_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1836 t$5343 net1460 VGND VGND VPWR VPWR booth_b26_m24 sky130_fd_sc_hd__xor2_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1847 net1041 net601 net1025 net874 VGND VGND VPWR VPWR t$5349 sky130_fd_sc_hd__a22o_1
XU$$1858 t$5354 net1459 VGND VGND VPWR VPWR booth_b26_m35 sky130_fd_sc_hd__xor2_1
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1869 net930 net600 net1751 net873 VGND VGND VPWR VPWR t$5360 sky130_fd_sc_hd__a22o_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0820_ clknet_leaf_106_clk booth_b38_m54 VGND VGND VPWR VPWR pp_row92_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_127_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0751_ clknet_leaf_160_clk booth_b36_m53 VGND VGND VPWR VPWR pp_row89_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_171_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0682_ clknet_leaf_176_clk booth_b46_m40 VGND VGND VPWR VPWR pp_row86_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_192_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2421_ clknet_leaf_142_clk booth_b24_m43 VGND VGND VPWR VPWR pp_row67_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_124_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_217_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_217_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2352_ clknet_leaf_77_clk booth_b34_m31 VGND VGND VPWR VPWR pp_row65_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_70_4 s$713 s$715 s$717 VGND VGND VPWR VPWR c$1574 s$1575 sky130_fd_sc_hd__fa_2
XFILLER_123_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1303_ clknet_leaf_1_clk booth_b12_m16 VGND VGND VPWR VPWR pp_row28_6 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_63_3 c$580 s$583 s$585 VGND VGND VPWR VPWR c$1488 s$1489 sky130_fd_sc_hd__fa_1
X_2283_ clknet_leaf_181_clk net156 VGND VGND VPWR VPWR pp_row124_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_97_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_56_2 c$448 c$450 c$452 VGND VGND VPWR VPWR c$1402 s$1403 sky130_fd_sc_hd__fa_1
XFILLER_56_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1234_ clknet_leaf_13_clk booth_b8_m16 VGND VGND VPWR VPWR pp_row24_4 sky130_fd_sc_hd__dfxtp_1
XU$$4440 net1086 sel_0$6647 net1076 net695 VGND VGND VPWR VPWR t$6674 sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_33_1 s$2889 s$2891 s$2893 VGND VGND VPWR VPWR c$3530 s$3531 sky130_fd_sc_hd__fa_1
XFILLER_93_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4451 t$6679 net1846 VGND VGND VPWR VPWR booth_b64_m30 sky130_fd_sc_hd__xor2_1
XU$$4462 net980 sel_0$6647 net971 net697 VGND VGND VPWR VPWR t$6685 sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_49_1 c$316 c$318 c$320 VGND VGND VPWR VPWR c$1316 s$1317 sky130_fd_sc_hd__fa_1
X_1165_ clknet_leaf_50_clk booth_b10_m9 VGND VGND VPWR VPWR pp_row19_5 sky130_fd_sc_hd__dfxtp_1
XU$$4473 t$6690 net1857 VGND VGND VPWR VPWR booth_b64_m41 sky130_fd_sc_hd__xor2_1
XU$$4484 net1710 sel_0$6647 net1702 net696 VGND VGND VPWR VPWR t$6696 sky130_fd_sc_hd__a22o_1
XU$$3750 t$6321 net1300 VGND VGND VPWR VPWR booth_b54_m22 sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_26_0 c$2840 c$2842 c$2844 VGND VGND VPWR VPWR c$3500 s$3501 sky130_fd_sc_hd__fa_1
XU$$4495 t$6701 net1868 VGND VGND VPWR VPWR booth_b64_m52 sky130_fd_sc_hd__xor2_1
XU$$3761 net1060 net469 net1051 net742 VGND VGND VPWR VPWR t$6327 sky130_fd_sc_hd__a22o_1
XU$$3772 t$6332 net1301 VGND VGND VPWR VPWR booth_b54_m33 sky130_fd_sc_hd__xor2_1
X_1096_ clknet_leaf_60_clk booth_b4_m9 VGND VGND VPWR VPWR pp_row13_2 sky130_fd_sc_hd__dfxtp_1
XU$$3783 net954 net470 net946 net743 VGND VGND VPWR VPWR t$6338 sky130_fd_sc_hd__a22o_1
XU$$3794 t$6343 net1307 VGND VGND VPWR VPWR booth_b54_m44 sky130_fd_sc_hd__xor2_1
XFILLER_33_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1998_ clknet_leaf_69_clk booth_b32_m23 VGND VGND VPWR VPWR pp_row55_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_147_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0949_ clknet_leaf_113_clk booth_b46_m52 VGND VGND VPWR VPWR pp_row98_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_107_817 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_100_0 c$3284 c$3286 c$3288 VGND VGND VPWR VPWR c$3796 s$3797 sky130_fd_sc_hd__fa_1
XFILLER_162_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_208_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_208_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_88_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_872 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_51_1 pp_row51_3 pp_row51_4 pp_row51_5 VGND VGND VPWR VPWR c$368 s$369
+ sky130_fd_sc_hd__fa_1
XU$$905 t$4867 net1314 VGND VGND VPWR VPWR booth_b12_m38 sky130_fd_sc_hd__xor2_1
XFILLER_141_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$916 net1733 net399 net1724 net665 VGND VGND VPWR VPWR t$4873 sky130_fd_sc_hd__a22o_1
XU$$927 t$4878 net1317 VGND VGND VPWR VPWR booth_b12_m49 sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_44_0 pp_row44_0 pp_row44_1 pp_row44_2 VGND VGND VPWR VPWR c$264 s$265
+ sky130_fd_sc_hd__fa_1
XFILLER_83_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$938 net1623 net399 net1615 net665 VGND VGND VPWR VPWR t$4884 sky130_fd_sc_hd__a22o_1
XFILLER_55_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$949 t$4889 net1317 VGND VGND VPWR VPWR booth_b12_m60 sky130_fd_sc_hd__xor2_1
XFILLER_189_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1085 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_923 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_80_3 s$1691 s$1693 s$1695 VGND VGND VPWR VPWR c$2484 s$2485 sky130_fd_sc_hd__fa_1
XFILLER_166_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_978 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_73_2 c$1600 s$1603 s$1605 VGND VGND VPWR VPWR c$2426 s$2427 sky130_fd_sc_hd__fa_1
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1200 net69 VGND VGND VPWR VPWR net1200 sky130_fd_sc_hd__buf_4
XFILLER_3_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1211 net1212 VGND VGND VPWR VPWR net1211 sky130_fd_sc_hd__buf_4
XFILLER_105_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_66_1 c$1510 c$1512 c$1514 VGND VGND VPWR VPWR c$2368 s$2369 sky130_fd_sc_hd__fa_1
XFILLER_39_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1222 net1223 VGND VGND VPWR VPWR net1222 sky130_fd_sc_hd__buf_6
XFILLER_26_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1233 net1234 VGND VGND VPWR VPWR net1233 sky130_fd_sc_hd__buf_6
XFILLER_182_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1244 net1245 VGND VGND VPWR VPWR net1244 sky130_fd_sc_hd__buf_6
Xdadda_fa_6_43_0 c$3564 c$3566 s$3569 VGND VGND VPWR VPWR c$3982 s$3983 sky130_fd_sc_hd__fa_1
Xfanout1255 net1257 VGND VGND VPWR VPWR net1255 sky130_fd_sc_hd__clkbuf_8
Xdadda_fa_3_59_0 s$527 c$1422 c$1424 VGND VGND VPWR VPWR c$2310 s$2311 sky130_fd_sc_hd__fa_1
Xfanout1266 net1267 VGND VGND VPWR VPWR net1266 sky130_fd_sc_hd__buf_2
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1277 net1278 VGND VGND VPWR VPWR net1277 sky130_fd_sc_hd__buf_6
Xfanout1288 net1290 VGND VGND VPWR VPWR net1288 sky130_fd_sc_hd__buf_6
XU$$3002 t$5938 net1373 VGND VGND VPWR VPWR booth_b42_m59 sky130_fd_sc_hd__xor2_1
Xfanout1299 net53 VGND VGND VPWR VPWR net1299 sky130_fd_sc_hd__buf_6
XU$$3013 net1374 VGND VGND VPWR VPWR notsign$5944 sky130_fd_sc_hd__inv_1
XFILLER_47_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3024 net1125 net511 net1034 net784 VGND VGND VPWR VPWR t$5951 sky130_fd_sc_hd__a22o_1
XFILLER_19_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3035 t$5956 net1362 VGND VGND VPWR VPWR booth_b44_m7 sky130_fd_sc_hd__xor2_1
XFILLER_46_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2301 t$5580 net1434 VGND VGND VPWR VPWR booth_b32_m51 sky130_fd_sc_hd__xor2_1
XU$$3046 net1206 net517 net1198 net790 VGND VGND VPWR VPWR t$5962 sky130_fd_sc_hd__a22o_1
XU$$2312 net1606 net574 net1598 net847 VGND VGND VPWR VPWR t$5586 sky130_fd_sc_hd__a22o_1
XU$$3057 t$5967 net1358 VGND VGND VPWR VPWR booth_b44_m18 sky130_fd_sc_hd__xor2_1
XU$$2323 t$5591 net1437 VGND VGND VPWR VPWR booth_b32_m62 sky130_fd_sc_hd__xor2_1
XU$$3068 net1096 net515 net1087 net788 VGND VGND VPWR VPWR t$5973 sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_102_2 s$2657 s$2659 s$2661 VGND VGND VPWR VPWR c$3306 s$3307 sky130_fd_sc_hd__fa_1
XFILLER_35_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2334 net28 net1435 VGND VGND VPWR VPWR sel_1$5598 sky130_fd_sc_hd__xor2_2
XFILLER_62_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3079 t$5978 net1357 VGND VGND VPWR VPWR booth_b44_m29 sky130_fd_sc_hd__xor2_1
XFILLER_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1600 t$5222 net1480 VGND VGND VPWR VPWR booth_b22_m43 sky130_fd_sc_hd__xor2_1
XU$$2345 net1672 net561 net1561 net834 VGND VGND VPWR VPWR t$5604 sky130_fd_sc_hd__a22o_1
XU$$2356 t$5609 net1420 VGND VGND VPWR VPWR booth_b34_m10 sky130_fd_sc_hd__xor2_1
XU$$1611 net1687 net616 net1679 net889 VGND VGND VPWR VPWR t$5228 sky130_fd_sc_hd__a22o_1
XU$$2367 net1170 net563 net1161 net836 VGND VGND VPWR VPWR t$5615 sky130_fd_sc_hd__a22o_1
XU$$1622 t$5233 net1483 VGND VGND VPWR VPWR booth_b22_m54 sky130_fd_sc_hd__xor2_1
XU$$2378 t$5620 net1424 VGND VGND VPWR VPWR booth_b34_m21 sky130_fd_sc_hd__xor2_1
XU$$1633 net1579 net617 net1553 net890 VGND VGND VPWR VPWR t$5239 sky130_fd_sc_hd__a22o_1
XU$$1644 net1481 VGND VGND VPWR VPWR notblock$5245\[0\] sky130_fd_sc_hd__inv_1
XU$$2389 net1065 net562 net1059 net835 VGND VGND VPWR VPWR t$5626 sky130_fd_sc_hd__a22o_1
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1655 t$5251 net1467 VGND VGND VPWR VPWR booth_b24_m2 sky130_fd_sc_hd__xor2_1
XFILLER_61_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1666 net1515 net605 net1508 net878 VGND VGND VPWR VPWR t$5257 sky130_fd_sc_hd__a22o_1
XU$$1677 t$5262 net1469 VGND VGND VPWR VPWR booth_b24_m13 sky130_fd_sc_hd__xor2_1
X_1921_ clknet_leaf_80_clk booth_b10_m43 VGND VGND VPWR VPWR pp_row53_5 sky130_fd_sc_hd__dfxtp_1
XU$$1688 net1138 net602 net1130 net875 VGND VGND VPWR VPWR t$5268 sky130_fd_sc_hd__a22o_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1699 t$5273 net1468 VGND VGND VPWR VPWR booth_b24_m24 sky130_fd_sc_hd__xor2_1
XFILLER_187_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1852_ clknet_leaf_25_clk net1332 VGND VGND VPWR VPWR pp_row50_26 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_7_116_0 s$3863 c$4126 s$4129 VGND VGND VPWR VPWR c$4384 s$4385 sky130_fd_sc_hd__fa_1
XFILLER_129_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0803_ clknet_leaf_94_clk booth_b46_m45 VGND VGND VPWR VPWR pp_row91_10 sky130_fd_sc_hd__dfxtp_1
X_1783_ clknet_leaf_184_clk net136 VGND VGND VPWR VPWR pp_row106_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_155_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0734_ clknet_leaf_163_clk booth_b48_m40 VGND VGND VPWR VPWR pp_row88_13 sky130_fd_sc_hd__dfxtp_1
X_0665_ clknet_leaf_187_clk booth_b62_m23 VGND VGND VPWR VPWR pp_row85_21 sky130_fd_sc_hd__dfxtp_1
X_2404_ clknet_leaf_99_clk booth_b60_m6 VGND VGND VPWR VPWR pp_row66_30 sky130_fd_sc_hd__dfxtp_1
XFILLER_130_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0596_ clknet_leaf_193_clk booth_b34_m49 VGND VGND VPWR VPWR pp_row83_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_69_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2335_ clknet_leaf_86_clk booth_b4_m61 VGND VGND VPWR VPWR pp_row65_2 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_61_0 s$59 c$528 c$530 VGND VGND VPWR VPWR c$1458 s$1459 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$307 final_adder.p_new$306 final_adder.g_new$309 final_adder.g_new$307
+ VGND VGND VPWR VPWR final_adder.g_new$435 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$318 final_adder.p_new$320 final_adder.p_new$318 VGND VGND VPWR VPWR
+ final_adder.p_new$446 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$329 final_adder.p_new$328 final_adder.g_new$331 final_adder.g_new$329
+ VGND VGND VPWR VPWR final_adder.g_new$457 sky130_fd_sc_hd__a21o_1
XFILLER_38_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2266_ clknet_leaf_214_clk booth_b12_m51 VGND VGND VPWR VPWR pp_row63_6 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_5_4__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_5_4__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_1217_ clknet_leaf_47_clk booth_b2_m21 VGND VGND VPWR VPWR pp_row23_1 sky130_fd_sc_hd__dfxtp_1
X_2197_ clknet_leaf_228_clk booth_b18_m43 VGND VGND VPWR VPWR pp_row61_9 sky130_fd_sc_hd__dfxtp_1
XU$$4270 t$6587 net1254 VGND VGND VPWR VPWR booth_b62_m8 sky130_fd_sc_hd__xor2_1
XFILLER_168_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4281 net1196 net418 net1177 net700 VGND VGND VPWR VPWR t$6593 sky130_fd_sc_hd__a22o_1
XFILLER_53_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4292 t$6598 net1255 VGND VGND VPWR VPWR booth_b62_m19 sky130_fd_sc_hd__xor2_1
XFILLER_77_1047 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1148_ clknet_leaf_15_clk booth_b4_m14 VGND VGND VPWR VPWR pp_row18_2 sky130_fd_sc_hd__dfxtp_1
XU$$3580 net1566 net481 net1525 net754 VGND VGND VPWR VPWR t$6235 sky130_fd_sc_hd__a22o_1
XU$$3591 t$6240 net1320 VGND VGND VPWR VPWR booth_b52_m11 sky130_fd_sc_hd__xor2_1
XFILLER_81_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_818 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1079_ clknet_leaf_52_clk booth_b6_m5 VGND VGND VPWR VPWR pp_row11_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_52_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2890 t$5882 net1368 VGND VGND VPWR VPWR booth_b42_m3 sky130_fd_sc_hd__xor2_1
XFILLER_179_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_90_2 s$2561 s$2563 s$2565 VGND VGND VPWR VPWR c$3234 s$3235 sky130_fd_sc_hd__fa_1
XFILLER_146_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_83_1 c$2498 c$2500 s$2503 VGND VGND VPWR VPWR c$3190 s$3191 sky130_fd_sc_hd__fa_1
XFILLER_101_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_60_0 s$3639 c$4014 s$4017 VGND VGND VPWR VPWR c$4272 s$4273 sky130_fd_sc_hd__fa_1
XFILLER_175_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_76_0 s$1649 c$2438 c$2440 VGND VGND VPWR VPWR c$3146 s$3147 sky130_fd_sc_hd__fa_1
XFILLER_134_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$841 final_adder.p_new$872 final_adder.g_new$937 final_adder.g_new$873
+ VGND VGND VPWR VPWR final_adder.g_new$969 sky130_fd_sc_hd__a21o_2
Xfinal_adder.U$$863 final_adder.p_new$894 final_adder.g_new$959 final_adder.g_new$895
+ VGND VGND VPWR VPWR final_adder.g_new$991 sky130_fd_sc_hd__a21o_2
XU$$702 t$4764 net1415 VGND VGND VPWR VPWR booth_b10_m5 sky130_fd_sc_hd__xor2_1
XFILLER_1_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$713 net1224 net404 net1216 net670 VGND VGND VPWR VPWR t$4770 sky130_fd_sc_hd__a22o_1
XU$$724 t$4775 net1412 VGND VGND VPWR VPWR booth_b10_m16 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$885 final_adder.p_new$916 final_adder.g_new$749 final_adder.g_new$917
+ VGND VGND VPWR VPWR final_adder.g_new$1013 sky130_fd_sc_hd__a21o_1
XU$$735 net1106 net402 net1099 net668 VGND VGND VPWR VPWR t$4781 sky130_fd_sc_hd__a22o_1
XFILLER_16_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$746 t$4786 net1416 VGND VGND VPWR VPWR booth_b10_m27 sky130_fd_sc_hd__xor2_1
XU$$757 net998 net402 net990 net668 VGND VGND VPWR VPWR t$4792 sky130_fd_sc_hd__a22o_1
XFILLER_43_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$768 t$4797 net1413 VGND VGND VPWR VPWR booth_b10_m38 sky130_fd_sc_hd__xor2_1
XU$$779 net1736 net405 net1725 net671 VGND VGND VPWR VPWR t$4803 sky130_fd_sc_hd__a22o_1
XFILLER_182_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_7 c$628 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0450_ clknet_leaf_158_clk booth_b28_m50 VGND VGND VPWR VPWR pp_row78_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_113_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0381_ clknet_leaf_204_clk booth_b14_m62 VGND VGND VPWR VPWR pp_row76_2 sky130_fd_sc_hd__dfxtp_1
Xfanout1030 net88 VGND VGND VPWR VPWR net1030 sky130_fd_sc_hd__buf_6
Xfanout1041 net1042 VGND VGND VPWR VPWR net1041 sky130_fd_sc_hd__buf_4
XFILLER_39_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2120_ clknet_leaf_218_clk booth_b8_m51 VGND VGND VPWR VPWR pp_row59_4 sky130_fd_sc_hd__dfxtp_1
Xfanout1052 net1053 VGND VGND VPWR VPWR net1052 sky130_fd_sc_hd__buf_2
Xfanout1063 net1064 VGND VGND VPWR VPWR net1063 sky130_fd_sc_hd__buf_4
Xfanout1074 net1075 VGND VGND VPWR VPWR net1074 sky130_fd_sc_hd__buf_4
Xfanout1085 net1086 VGND VGND VPWR VPWR net1085 sky130_fd_sc_hd__buf_4
Xfanout1096 net80 VGND VGND VPWR VPWR net1096 sky130_fd_sc_hd__clkbuf_8
X_2051_ clknet_leaf_38_clk booth_b8_m49 VGND VGND VPWR VPWR pp_row57_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_94_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_40_5 s$229 s$231 s$233 VGND VGND VPWR VPWR c$1216 s$1217 sky130_fd_sc_hd__fa_1
X_1002_ clknet_leaf_118_clk booth_b44_m57 VGND VGND VPWR VPWR pp_row101_4 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_33_4 pp_row33_12 pp_row33_13 pp_row33_14 VGND VGND VPWR VPWR c$1130 s$1131
+ sky130_fd_sc_hd__fa_1
XFILLER_19_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2120 t$5488 net1442 VGND VGND VPWR VPWR booth_b30_m29 sky130_fd_sc_hd__xor2_1
XU$$2131 net989 net580 net978 net853 VGND VGND VPWR VPWR t$5494 sky130_fd_sc_hd__a22o_1
XU$$2142 t$5499 net1446 VGND VGND VPWR VPWR booth_b30_m40 sky130_fd_sc_hd__xor2_1
XFILLER_179_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2153 net1713 net578 net1704 net851 VGND VGND VPWR VPWR t$5505 sky130_fd_sc_hd__a22o_1
XU$$2164 t$5510 net1446 VGND VGND VPWR VPWR booth_b30_m51 sky130_fd_sc_hd__xor2_1
XU$$2175 net1605 net578 net1597 net851 VGND VGND VPWR VPWR t$5516 sky130_fd_sc_hd__a22o_1
XU$$1430 net1064 net628 net1056 net901 VGND VGND VPWR VPWR t$5136 sky130_fd_sc_hd__a22o_1
XU$$1441 t$5141 net1488 VGND VGND VPWR VPWR booth_b20_m32 sky130_fd_sc_hd__xor2_1
XU$$2186 t$5521 net1446 VGND VGND VPWR VPWR booth_b30_m62 sky130_fd_sc_hd__xor2_1
XFILLER_179_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2197 net26 net1444 VGND VGND VPWR VPWR sel_1$5528 sky130_fd_sc_hd__xor2_4
XU$$1452 net961 net631 net955 net904 VGND VGND VPWR VPWR t$5147 sky130_fd_sc_hd__a22o_1
XU$$1463 t$5152 net1492 VGND VGND VPWR VPWR booth_b20_m43 sky130_fd_sc_hd__xor2_1
XU$$1474 net1690 net634 net1682 net907 VGND VGND VPWR VPWR t$5158 sky130_fd_sc_hd__a22o_1
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1485 t$5163 net1492 VGND VGND VPWR VPWR booth_b20_m54 sky130_fd_sc_hd__xor2_1
XU$$1496 net1579 net633 net1553 net906 VGND VGND VPWR VPWR t$5169 sky130_fd_sc_hd__a22o_1
X_1904_ clknet_leaf_71_clk booth_b38_m14 VGND VGND VPWR VPWR pp_row52_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_187_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1835_ clknet_leaf_25_clk booth_b24_m26 VGND VGND VPWR VPWR pp_row50_12 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_93_0 c$3242 c$3244 c$3246 VGND VGND VPWR VPWR c$3768 s$3769 sky130_fd_sc_hd__fa_1
XFILLER_159_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1766_ clknet_leaf_236_clk booth_b4_m44 VGND VGND VPWR VPWR pp_row48_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_116_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0717_ clknet_leaf_179_clk booth_b64_m23 VGND VGND VPWR VPWR pp_row87_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_171_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1697_ clknet_leaf_19_clk booth_b30_m15 VGND VGND VPWR VPWR pp_row45_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_116_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0648_ clknet_leaf_183_clk booth_b30_m55 VGND VGND VPWR VPWR pp_row85_5 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_78_6 pp_row78_20 pp_row78_21 pp_row78_22 VGND VGND VPWR VPWR c$864 s$865
+ sky130_fd_sc_hd__fa_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0579_ clknet_leaf_205_clk booth_b52_m30 VGND VGND VPWR VPWR pp_row82_18 sky130_fd_sc_hd__dfxtp_1
XTAP_4109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$104 c$4358 s$4361 VGND VGND VPWR VPWR final_adder.$signal$210 final_adder.$signal$1194
+ sky130_fd_sc_hd__ha_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2318_ clknet_leaf_77_clk booth_b38_m26 VGND VGND VPWR VPWR pp_row64_19 sky130_fd_sc_hd__dfxtp_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$115 c$4380 s$4383 VGND VGND VPWR VPWR final_adder.$signal$232 final_adder.$signal$1205
+ sky130_fd_sc_hd__ha_1
XFILLER_39_940 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$126 c$4402 s$4405 VGND VGND VPWR VPWR final_adder.$signal$254 final_adder.$signal$1216
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$137 final_adder.$signal$1209 final_adder.$signal$238 final_adder.$signal$240
+ VGND VGND VPWR VPWR final_adder.g_new$265 sky130_fd_sc_hd__a21o_1
XTAP_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$148 final_adder.$signal$1196 final_adder.$signal$1197 VGND VGND VPWR
+ VPWR final_adder.p_new$276 sky130_fd_sc_hd__and2_1
XTAP_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$159 final_adder.$signal$1187 final_adder.$signal$194 final_adder.$signal$196
+ VGND VGND VPWR VPWR final_adder.g_new$287 sky130_fd_sc_hd__a21o_1
XFILLER_45_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2249_ clknet_leaf_136_clk booth_b54_m56 VGND VGND VPWR VPWR pp_row110_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_26_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_408 net1714 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_419 net492 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_102_1 pp_row102_14 pp_row102_15 c$1934 VGND VGND VPWR VPWR c$2656 s$2657
+ sky130_fd_sc_hd__fa_1
XFILLER_150_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput100 b[41] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_873 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput111 b[51] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__buf_6
XFILLER_88_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput122 b[61] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__buf_6
Xdadda_fa_6_123_0 c$3884 c$3886 s$3889 VGND VGND VPWR VPWR c$4142 s$4143 sky130_fd_sc_hd__fa_1
Xinput133 c[103] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_1
Xinput144 c[113] VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_759 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput155 c[123] VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_0_66_4 pp_row66_12 pp_row66_13 pp_row66_14 VGND VGND VPWR VPWR c$116 s$117
+ sky130_fd_sc_hd__fa_1
Xinput166 c[18] VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_1
Xinput177 c[28] VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_3_43_3 s$1247 s$1249 s$1251 VGND VGND VPWR VPWR c$2188 s$2189 sky130_fd_sc_hd__fa_1
XFILLER_76_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput188 c[38] VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_1
XFILLER_56_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput199 c[48] VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$660 final_adder.p_new$684 final_adder.p_new$668 VGND VGND VPWR VPWR
+ final_adder.p_new$788 sky130_fd_sc_hd__and2_1
XTAP_3942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1084 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$510 t$4665 net1252 VGND VGND VPWR VPWR booth_b6_m46 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$671 final_adder.p_new$678 final_adder.g_new$695 final_adder.g_new$679
+ VGND VGND VPWR VPWR final_adder.g_new$799 sky130_fd_sc_hd__a21o_1
XTAP_3953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$682 final_adder.p_new$706 final_adder.p_new$690 VGND VGND VPWR VPWR
+ final_adder.p_new$810 sky130_fd_sc_hd__and2_1
XU$$521 net1649 net432 net1641 net714 VGND VGND VPWR VPWR t$4671 sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_36_2 c$1156 s$1159 s$1161 VGND VGND VPWR VPWR c$2130 s$2131 sky130_fd_sc_hd__fa_1
XTAP_3964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$532 t$4676 net1246 VGND VGND VPWR VPWR booth_b6_m57 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$693 final_adder.p_new$700 final_adder.g_new$717 final_adder.g_new$701
+ VGND VGND VPWR VPWR final_adder.g_new$821 sky130_fd_sc_hd__a21o_1
XTAP_3975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$543 net1539 net432 net1531 net714 VGND VGND VPWR VPWR t$4682 sky130_fd_sc_hd__a22o_1
XFILLER_56_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_29_1 pp_row29_14 pp_row29_15 c$1074 VGND VGND VPWR VPWR c$2072 s$2073
+ sky130_fd_sc_hd__fa_1
XU$$554 net1882 net413 net1231 net679 VGND VGND VPWR VPWR t$4689 sky130_fd_sc_hd__a22o_1
XFILLER_186_1072 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$565 t$4694 net1240 VGND VGND VPWR VPWR booth_b8_m5 sky130_fd_sc_hd__xor2_1
XU$$576 net1224 net413 net1216 net679 VGND VGND VPWR VPWR t$4700 sky130_fd_sc_hd__a22o_1
XU$$587 t$4705 net1241 VGND VGND VPWR VPWR booth_b8_m16 sky130_fd_sc_hd__xor2_1
XFILLER_189_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$598 net1105 net409 net1097 net675 VGND VGND VPWR VPWR t$4711 sky130_fd_sc_hd__a22o_1
XFILLER_60_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1620_ clknet_leaf_5_clk booth_b34_m8 VGND VGND VPWR VPWR pp_row42_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_126_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1551_ clknet_leaf_240_clk booth_b0_m40 VGND VGND VPWR VPWR pp_row40_0 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_88_5 s$1003 s$1005 s$1007 VGND VGND VPWR VPWR c$1792 s$1793 sky130_fd_sc_hd__fa_1
X_0502_ clknet_leaf_195_clk net233 VGND VGND VPWR VPWR pp_row79_26 sky130_fd_sc_hd__dfxtp_1
XFILLER_114_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1482_ clknet_leaf_241_clk booth_b4_m33 VGND VGND VPWR VPWR pp_row37_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_113_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0433_ clknet_leaf_131_clk notsign$6224 VGND VGND VPWR VPWR pp_row115_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_98_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0364_ clknet_leaf_204_clk booth_b40_m35 VGND VGND VPWR VPWR pp_row75_15 sky130_fd_sc_hd__dfxtp_1
X_2103_ clknet_leaf_30_clk booth_b42_m16 VGND VGND VPWR VPWR pp_row58_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_95_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0295_ clknet_leaf_199_clk booth_b30_m43 VGND VGND VPWR VPWR pp_row73_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_54_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2034_ clknet_leaf_73_clk booth_b40_m16 VGND VGND VPWR VPWR pp_row56_20 sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_31_1 pp_row31_3 pp_row31_4 pp_row31_5 VGND VGND VPWR VPWR c$1102 s$1103
+ sky130_fd_sc_hd__fa_1
XFILLER_130_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_24_0 pp_row24_0 pp_row24_1 pp_row24_2 VGND VGND VPWR VPWR c$1054 s$1055
+ sky130_fd_sc_hd__fa_1
XFILLER_161_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1260 t$5049 net1662 VGND VGND VPWR VPWR booth_b18_m10 sky130_fd_sc_hd__xor2_1
XFILLER_50_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1271 net1170 net638 net1161 net911 VGND VGND VPWR VPWR t$5055 sky130_fd_sc_hd__a22o_1
XU$$1282 t$5060 net1662 VGND VGND VPWR VPWR booth_b18_m21 sky130_fd_sc_hd__xor2_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1293 net1064 net639 net1055 net912 VGND VGND VPWR VPWR t$5066 sky130_fd_sc_hd__a22o_1
Xdadda_ha_1_84_6 pp_row84_18 pp_row84_19 VGND VGND VPWR VPWR c$964 s$965 sky130_fd_sc_hd__ha_1
Xdadda_fa_5_118_1 s$3399 s$3401 s$3403 VGND VGND VPWR VPWR c$3870 s$3871 sky130_fd_sc_hd__fa_2
XFILLER_11_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1376_1760 VGND VGND VPWR VPWR U$$1376_1760/HI net1760 sky130_fd_sc_hd__conb_1
X_1818_ clknet_leaf_222_clk booth_b44_m5 VGND VGND VPWR VPWR pp_row49_22 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1749_ clknet_leaf_234_clk booth_b24_m23 VGND VGND VPWR VPWR pp_row47_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_2_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_83_4 pp_row83_12 pp_row83_13 pp_row83_14 VGND VGND VPWR VPWR c$946 s$947
+ sky130_fd_sc_hd__fa_1
XFILLER_117_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout801 net803 VGND VGND VPWR VPWR net801 sky130_fd_sc_hd__buf_2
Xfanout812 net815 VGND VGND VPWR VPWR net812 sky130_fd_sc_hd__buf_4
Xfanout823 sel_1$5738 VGND VGND VPWR VPWR net823 sky130_fd_sc_hd__buf_6
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_76_3 pp_row76_14 pp_row76_15 pp_row76_16 VGND VGND VPWR VPWR c$822 s$823
+ sky130_fd_sc_hd__fa_1
Xfanout834 net835 VGND VGND VPWR VPWR net834 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout845 sel_1$5528 VGND VGND VPWR VPWR net845 sky130_fd_sc_hd__buf_6
Xdadda_fa_4_53_2 s$2265 s$2267 s$2269 VGND VGND VPWR VPWR c$3012 s$3013 sky130_fd_sc_hd__fa_1
Xfanout856 sel_1$5458 VGND VGND VPWR VPWR net856 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_69_2 pp_row69_21 pp_row69_22 pp_row69_23 VGND VGND VPWR VPWR c$694 s$695
+ sky130_fd_sc_hd__fa_1
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout867 net868 VGND VGND VPWR VPWR net867 sky130_fd_sc_hd__clkbuf_2
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout878 net879 VGND VGND VPWR VPWR net878 sky130_fd_sc_hd__buf_4
XFILLER_85_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout889 net891 VGND VGND VPWR VPWR net889 sky130_fd_sc_hd__buf_4
Xdadda_fa_4_46_1 c$2202 c$2204 s$2207 VGND VGND VPWR VPWR c$2968 s$2969 sky130_fd_sc_hd__fa_1
XFILLER_100_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_23_0 s$3491 c$3940 s$3943 VGND VGND VPWR VPWR c$4198 s$4199 sky130_fd_sc_hd__fa_1
XTAP_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_39_0 s$1205 c$2142 c$2144 VGND VGND VPWR VPWR c$2924 s$2925 sky130_fd_sc_hd__fa_1
XTAP_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_205 net1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_216 net1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_227 net1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_238 net1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_249 net1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_0_71_2 pp_row71_6 pp_row71_7 pp_row71_8 VGND VGND VPWR VPWR c$168 s$169
+ sky130_fd_sc_hd__fa_1
XFILLER_122_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_0_64_1 pp_row64_3 pp_row64_4 pp_row64_5 VGND VGND VPWR VPWR c$86 s$87 sky130_fd_sc_hd__fa_2
XFILLER_76_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_41_0 s$243 c$1206 c$1208 VGND VGND VPWR VPWR c$2166 s$2167 sky130_fd_sc_hd__fa_1
XFILLER_190_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_0_57_0 pp_row57_0 pp_row57_1 pp_row57_2 VGND VGND VPWR VPWR c$18 s$19 sky130_fd_sc_hd__fa_1
XFILLER_92_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_1099 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$0_1753 VGND VGND VPWR VPWR U$$0_1753/HI net1753 sky130_fd_sc_hd__conb_1
XFILLER_64_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$490 final_adder.p_new$496 final_adder.p_new$492 VGND VGND VPWR VPWR
+ final_adder.p_new$618 sky130_fd_sc_hd__and2_1
XTAP_3772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$340 net1042 net534 net1026 net807 VGND VGND VPWR VPWR t$4579 sky130_fd_sc_hd__a22o_1
XFILLER_18_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$351 t$4584 net1279 VGND VGND VPWR VPWR booth_b4_m35 sky130_fd_sc_hd__xor2_1
XTAP_3794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$362 net925 net530 net1746 net803 VGND VGND VPWR VPWR t$4590 sky130_fd_sc_hd__a22o_1
XFILLER_91_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$373 t$4595 net1275 VGND VGND VPWR VPWR booth_b4_m46 sky130_fd_sc_hd__xor2_1
XFILLER_44_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$384 net1649 net534 net1641 net807 VGND VGND VPWR VPWR t$4601 sky130_fd_sc_hd__a22o_1
XU$$395 t$4606 net1275 VGND VGND VPWR VPWR booth_b4_m57 sky130_fd_sc_hd__xor2_1
XFILLER_32_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0982_ clknet_leaf_115_clk booth_b40_m60 VGND VGND VPWR VPWR pp_row100_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_158_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1603_ clknet_leaf_240_clk booth_b6_m36 VGND VGND VPWR VPWR pp_row42_3 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_93_3 pp_row93_15 pp_row93_16 pp_row93_17 VGND VGND VPWR VPWR c$1848 s$1849
+ sky130_fd_sc_hd__fa_1
XFILLER_172_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_86_2 pp_row86_23 c$966 c$968 VGND VGND VPWR VPWR c$1762 s$1763 sky130_fd_sc_hd__fa_2
X_1534_ clknet_leaf_16_clk booth_b12_m27 VGND VGND VPWR VPWR pp_row39_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_99_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_63_1 s$3069 s$3071 s$3073 VGND VGND VPWR VPWR c$3650 s$3651 sky130_fd_sc_hd__fa_1
XFILLER_113_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_79_1 c$856 c$858 c$860 VGND VGND VPWR VPWR c$1676 s$1677 sky130_fd_sc_hd__fa_1
XFILLER_114_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1465_ clknet_leaf_39_clk booth_b14_m22 VGND VGND VPWR VPWR pp_row36_7 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_56_0 c$3020 c$3022 c$3024 VGND VGND VPWR VPWR c$3620 s$3621 sky130_fd_sc_hd__fa_1
XFILLER_68_832 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0416_ clknet_leaf_155_clk booth_b20_m57 VGND VGND VPWR VPWR pp_row77_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_41_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1396_ clknet_leaf_54_clk booth_b2_m31 VGND VGND VPWR VPWR pp_row33_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1367_1759 VGND VGND VPWR VPWR U$$1367_1759/HI net1759 sky130_fd_sc_hd__conb_1
Xdadda_fa_1_55_8 c$4 c$6 s$9 VGND VGND VPWR VPWR c$454 s$455 sky130_fd_sc_hd__fa_1
X_0347_ clknet_leaf_197_clk net228 VGND VGND VPWR VPWR pp_row74_29 sky130_fd_sc_hd__dfxtp_1
X_0278_ clknet_leaf_179_clk booth_b64_m61 VGND VGND VPWR VPWR pp_row125_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_42_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2017_ clknet_leaf_81_clk booth_b8_m48 VGND VGND VPWR VPWR pp_row56_4 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_102_0 net1905 pp_row102_1 pp_row102_2 VGND VGND VPWR VPWR c$1942 s$1943
+ sky130_fd_sc_hd__fa_1
XFILLER_168_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_940 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1090 t$4961 net1188 VGND VGND VPWR VPWR booth_b14_m62 sky130_fd_sc_hd__xor2_1
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2326_1774 VGND VGND VPWR VPWR U$$2326_1774/HI net1774 sky130_fd_sc_hd__conb_1
XFILLER_164_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_81_1 pp_row81_3 pp_row81_4 pp_row81_5 VGND VGND VPWR VPWR c$908 s$909
+ sky130_fd_sc_hd__fa_1
XFILLER_104_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1607 net1611 VGND VGND VPWR VPWR net1607 sky130_fd_sc_hd__buf_4
Xfanout1618 net1619 VGND VGND VPWR VPWR net1618 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_74_0 pp_row74_8 pp_row74_9 pp_row74_10 VGND VGND VPWR VPWR c$780 s$781
+ sky130_fd_sc_hd__fa_1
Xfanout620 net622 VGND VGND VPWR VPWR net620 sky130_fd_sc_hd__clkbuf_4
XFILLER_144_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout631 sel_0$5107 VGND VGND VPWR VPWR net631 sky130_fd_sc_hd__buf_4
Xfanout1629 net1630 VGND VGND VPWR VPWR net1629 sky130_fd_sc_hd__buf_4
XFILLER_99_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout642 sel_0$5037 VGND VGND VPWR VPWR net642 sky130_fd_sc_hd__buf_6
Xfanout653 net655 VGND VGND VPWR VPWR net653 sky130_fd_sc_hd__buf_4
Xfanout664 net665 VGND VGND VPWR VPWR net664 sky130_fd_sc_hd__clkbuf_4
Xfanout675 net678 VGND VGND VPWR VPWR net675 sky130_fd_sc_hd__buf_4
Xfanout686 net687 VGND VGND VPWR VPWR net686 sky130_fd_sc_hd__buf_4
XFILLER_100_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout697 net699 VGND VGND VPWR VPWR net697 sky130_fd_sc_hd__clkbuf_4
XTAP_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3409 t$6146 net1345 VGND VGND VPWR VPWR booth_b48_m57 sky130_fd_sc_hd__xor2_1
XTAP_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2708 t$5788 net1398 VGND VGND VPWR VPWR booth_b38_m49 sky130_fd_sc_hd__xor2_1
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2719 net1627 net547 net1619 net820 VGND VGND VPWR VPWR t$5794 sky130_fd_sc_hd__a22o_1
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_96_1 c$1870 c$1872 c$1874 VGND VGND VPWR VPWR c$2608 s$2609 sky130_fd_sc_hd__fa_1
Xdadda_fa_6_73_0 c$3684 c$3686 s$3689 VGND VGND VPWR VPWR c$4042 s$4043 sky130_fd_sc_hd__fa_1
XFILLER_120_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_89_0 s$1017 c$1782 c$1784 VGND VGND VPWR VPWR c$2550 s$2551 sky130_fd_sc_hd__fa_2
XFILLER_135_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1250_ clknet_leaf_10_clk booth_b6_m19 VGND VGND VPWR VPWR pp_row25_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_96_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0201_ clknet_leaf_153_clk booth_b42_m28 VGND VGND VPWR VPWR pp_row70_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_77_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1181_ clknet_leaf_49_clk booth_b16_m4 VGND VGND VPWR VPWR pp_row20_8 sky130_fd_sc_hd__dfxtp_1
XU$$3910 net997 net465 net988 net738 VGND VGND VPWR VPWR t$6403 sky130_fd_sc_hd__a22o_1
XU$$3921 t$6408 net1299 VGND VGND VPWR VPWR booth_b56_m39 sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_118_0 net1912 pp_row118_1 pp_row118_2 VGND VGND VPWR VPWR c$3398 s$3399
+ sky130_fd_sc_hd__fa_1
XTAP_4270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3932 net1726 net466 net1718 net739 VGND VGND VPWR VPWR t$6414 sky130_fd_sc_hd__a22o_1
XTAP_4281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3943 t$6419 net1297 VGND VGND VPWR VPWR booth_b56_m50 sky130_fd_sc_hd__xor2_1
XTAP_4292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3954 net1616 net465 net1608 net738 VGND VGND VPWR VPWR t$6425 sky130_fd_sc_hd__a22o_1
Xdadda_ha_5_5_0 pp_row5_0 pp_row5_1 VGND VGND VPWR VPWR c$3418 s$3419 sky130_fd_sc_hd__ha_1
XFILLER_40_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3965 t$6430 net1292 VGND VGND VPWR VPWR booth_b56_m61 sky130_fd_sc_hd__xor2_1
XU$$3976 net1284 notblock$6435\[1\] VGND VGND VPWR VPWR t$6436 sky130_fd_sc_hd__and2_1
XTAP_3580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3987 net935 net452 net1674 net725 VGND VGND VPWR VPWR t$6443 sky130_fd_sc_hd__a22o_1
XU$$3998 t$6448 net1287 VGND VGND VPWR VPWR booth_b58_m9 sky130_fd_sc_hd__xor2_1
XTAP_3591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$170 t$4492 net1386 VGND VGND VPWR VPWR booth_b2_m13 sky130_fd_sc_hd__xor2_1
XU$$181 net1143 net623 net1133 net896 VGND VGND VPWR VPWR t$4498 sky130_fd_sc_hd__a22o_1
XFILLER_32_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$192 t$4503 net1385 VGND VGND VPWR VPWR booth_b2_m24 sky130_fd_sc_hd__xor2_1
XFILLER_162_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_180_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_180_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_193_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0965_ clknet_leaf_116_clk booth_b42_m57 VGND VGND VPWR VPWR pp_row99_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0896_ clknet_leaf_100_clk booth_b58_m37 VGND VGND VPWR VPWR pp_row95_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_134_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_91_0 pp_row91_9 pp_row91_10 pp_row91_11 VGND VGND VPWR VPWR c$1818 s$1819
+ sky130_fd_sc_hd__fa_1
XFILLER_114_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput267 net267 VGND VGND VPWR VPWR o[109] sky130_fd_sc_hd__buf_2
XFILLER_88_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput278 net278 VGND VGND VPWR VPWR o[119] sky130_fd_sc_hd__buf_2
X_1517_ clknet_leaf_121_clk booth_b44_m61 VGND VGND VPWR VPWR pp_row105_2 sky130_fd_sc_hd__dfxtp_1
Xoutput289 net289 VGND VGND VPWR VPWR o[13] sky130_fd_sc_hd__buf_2
XFILLER_82_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2497_ clknet_leaf_97_clk booth_b34_m35 VGND VGND VPWR VPWR pp_row69_15 sky130_fd_sc_hd__dfxtp_1
Xdadda_ha_1_47_6 pp_row47_18 pp_row47_19 VGND VGND VPWR VPWR c$314 s$315 sky130_fd_sc_hd__ha_1
XFILLER_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1448_ clknet_leaf_56_clk booth_b22_m13 VGND VGND VPWR VPWR pp_row35_11 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_60_6 pp_row60_32 c$32 c$34 VGND VGND VPWR VPWR c$540 s$541 sky130_fd_sc_hd__fa_1
XU$$1230_1756 VGND VGND VPWR VPWR U$$1230_1756/HI net1756 sky130_fd_sc_hd__conb_1
XFILLER_56_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_53_5 pp_row53_17 pp_row53_18 pp_row53_19 VGND VGND VPWR VPWR c$412 s$413
+ sky130_fd_sc_hd__fa_1
X_1379_ clknet_leaf_35_clk booth_b14_m18 VGND VGND VPWR VPWR pp_row32_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_56_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_46_4 pp_row46_12 pp_row46_13 pp_row46_14 VGND VGND VPWR VPWR c$296 s$297
+ sky130_fd_sc_hd__fa_1
XFILLER_55_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_16_2 c$1976 s$1979 s$1981 VGND VGND VPWR VPWR c$2790 s$2791 sky130_fd_sc_hd__fa_1
XFILLER_12_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4443_1842 VGND VGND VPWR VPWR U$$4443_1842/HI net1842 sky130_fd_sc_hd__conb_1
XFILLER_90_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_171_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_171_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_23_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_90_0 s$3759 c$4074 s$4077 VGND VGND VPWR VPWR c$4332 s$4333 sky130_fd_sc_hd__fa_1
XFILLER_183_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1404 net1405 VGND VGND VPWR VPWR net1404 sky130_fd_sc_hd__buf_4
XFILLER_132_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1415 net1416 VGND VGND VPWR VPWR net1415 sky130_fd_sc_hd__buf_6
Xfanout1426 net1427 VGND VGND VPWR VPWR net1426 sky130_fd_sc_hd__buf_4
Xfanout1437 net1438 VGND VGND VPWR VPWR net1437 sky130_fd_sc_hd__clkbuf_16
Xfanout450 sel_0 VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__buf_6
Xfanout1448 net1450 VGND VGND VPWR VPWR net1448 sky130_fd_sc_hd__buf_6
Xfanout1459 net20 VGND VGND VPWR VPWR net1459 sky130_fd_sc_hd__buf_6
Xfanout461 sel_0$6367 VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__clkbuf_4
Xfanout472 net475 VGND VGND VPWR VPWR net472 sky130_fd_sc_hd__buf_6
XFILLER_47_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout483 sel_0$6227 VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__buf_4
XFILLER_115_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout494 net495 VGND VGND VPWR VPWR net494 sky130_fd_sc_hd__buf_4
XFILLER_48_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3206 t$6043 net1350 VGND VGND VPWR VPWR booth_b46_m24 sky130_fd_sc_hd__xor2_1
XU$$3217 net1043 net503 net1027 net776 VGND VGND VPWR VPWR t$6049 sky130_fd_sc_hd__a22o_1
XFILLER_4_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3228 t$6054 net1351 VGND VGND VPWR VPWR booth_b46_m35 sky130_fd_sc_hd__xor2_1
XFILLER_111_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3239 net927 net503 net1748 net776 VGND VGND VPWR VPWR t$6060 sky130_fd_sc_hd__a22o_1
XFILLER_73_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2505 t$5685 net1406 VGND VGND VPWR VPWR booth_b36_m16 sky130_fd_sc_hd__xor2_1
XFILLER_59_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2516 net1109 net552 net1101 net825 VGND VGND VPWR VPWR t$5691 sky130_fd_sc_hd__a22o_1
XU$$2527 t$5696 net1405 VGND VGND VPWR VPWR booth_b36_m27 sky130_fd_sc_hd__xor2_1
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2538 net1004 net557 net996 net830 VGND VGND VPWR VPWR t$5702 sky130_fd_sc_hd__a22o_1
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1804 t$5327 net1460 VGND VGND VPWR VPWR booth_b26_m8 sky130_fd_sc_hd__xor2_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2549 t$5707 net1405 VGND VGND VPWR VPWR booth_b36_m38 sky130_fd_sc_hd__xor2_1
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1815 net1192 net594 net1173 net867 VGND VGND VPWR VPWR t$5333 sky130_fd_sc_hd__a22o_1
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1826 t$5338 net1458 VGND VGND VPWR VPWR booth_b26_m19 sky130_fd_sc_hd__xor2_1
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1837 net1083 net596 net1074 net869 VGND VGND VPWR VPWR t$5344 sky130_fd_sc_hd__a22o_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1848 t$5349 net1460 VGND VGND VPWR VPWR booth_b26_m30 sky130_fd_sc_hd__xor2_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1859 net974 net595 net965 net868 VGND VGND VPWR VPWR t$5355 sky130_fd_sc_hd__a22o_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_162_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_162_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0750_ clknet_leaf_160_clk booth_b34_m55 VGND VGND VPWR VPWR pp_row89_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_128_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0681_ clknet_leaf_169_clk booth_b44_m42 VGND VGND VPWR VPWR pp_row86_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_115_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2420_ clknet_leaf_145_clk booth_b22_m45 VGND VGND VPWR VPWR pp_row67_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_124_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2351_ clknet_leaf_77_clk booth_b32_m33 VGND VGND VPWR VPWR pp_row65_16 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_70_5 s$719 s$721 s$723 VGND VGND VPWR VPWR c$1576 s$1577 sky130_fd_sc_hd__fa_2
XFILLER_151_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1302_ clknet_leaf_250_clk booth_b10_m18 VGND VGND VPWR VPWR pp_row28_5 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_63_4 s$587 s$589 s$591 VGND VGND VPWR VPWR c$1490 s$1491 sky130_fd_sc_hd__fa_1
X_2282_ clknet_leaf_129_clk booth_b60_m50 VGND VGND VPWR VPWR pp_row110_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_56_3 c$454 s$457 s$459 VGND VGND VPWR VPWR c$1404 s$1405 sky130_fd_sc_hd__fa_1
X_1233_ clknet_leaf_13_clk booth_b6_m18 VGND VGND VPWR VPWR pp_row24_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_78_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4430 net1135 sel_0$6647 net1119 net694 VGND VGND VPWR VPWR t$6669 sky130_fd_sc_hd__a22o_1
XU$$4441 t$6674 net1841 VGND VGND VPWR VPWR booth_b64_m25 sky130_fd_sc_hd__xor2_1
XU$$4452 net1030 sel_0$6647 net1022 net698 VGND VGND VPWR VPWR t$6680 sky130_fd_sc_hd__a22o_1
XFILLER_37_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_49_2 c$322 c$324 c$326 VGND VGND VPWR VPWR c$1318 s$1319 sky130_fd_sc_hd__fa_1
XU$$4463 t$6685 net1852 VGND VGND VPWR VPWR booth_b64_m36 sky130_fd_sc_hd__xor2_1
X_1164_ clknet_leaf_50_clk booth_b8_m11 VGND VGND VPWR VPWR pp_row19_4 sky130_fd_sc_hd__dfxtp_1
XU$$4474 net1747 sel_0$6647 net1739 net693 VGND VGND VPWR VPWR t$6691 sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_26_1 s$2847 s$2849 s$2851 VGND VGND VPWR VPWR c$3502 s$3503 sky130_fd_sc_hd__fa_2
XU$$3740 t$6316 net1301 VGND VGND VPWR VPWR booth_b54_m17 sky130_fd_sc_hd__xor2_1
XFILLER_93_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4485 t$6696 net1863 VGND VGND VPWR VPWR booth_b64_m47 sky130_fd_sc_hd__xor2_1
XU$$3751 net1102 net470 net1094 net743 VGND VGND VPWR VPWR t$6322 sky130_fd_sc_hd__a22o_1
XU$$4496 net1640 sel_0$6647 net1632 net695 VGND VGND VPWR VPWR t$6702 sky130_fd_sc_hd__a22o_1
XU$$3762 t$6327 net1303 VGND VGND VPWR VPWR booth_b54_m28 sky130_fd_sc_hd__xor2_1
X_1095_ clknet_leaf_59_clk booth_b2_m11 VGND VGND VPWR VPWR pp_row13_1 sky130_fd_sc_hd__dfxtp_1
XU$$3773 net997 net470 net988 net743 VGND VGND VPWR VPWR t$6333 sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_19_0 c$2798 c$2800 c$2802 VGND VGND VPWR VPWR c$3472 s$3473 sky130_fd_sc_hd__fa_1
XU$$3784 t$6338 net1301 VGND VGND VPWR VPWR booth_b54_m39 sky130_fd_sc_hd__xor2_1
XU$$3795 net1726 net474 net1717 net747 VGND VGND VPWR VPWR t$6344 sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_153_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_153_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_178_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1997_ clknet_leaf_69_clk booth_b30_m25 VGND VGND VPWR VPWR pp_row55_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_159_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0948_ clknet_leaf_113_clk booth_b44_m54 VGND VGND VPWR VPWR pp_row98_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_109_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_100_1 s$3291 s$3293 s$3295 VGND VGND VPWR VPWR c$3798 s$3799 sky130_fd_sc_hd__fa_2
XFILLER_107_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0879_ clknet_leaf_93_clk booth_b64_m30 VGND VGND VPWR VPWR pp_row94_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_133_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4473_1857 VGND VGND VPWR VPWR U$$4473_1857/HI net1857 sky130_fd_sc_hd__conb_1
Xdadda_ha_4_122_0 net1919 pp_row122_1 VGND VGND VPWR VPWR c$3414 s$3415 sky130_fd_sc_hd__ha_1
XFILLER_133_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_884 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_1_38_2 pp_row38_6 pp_row38_7 VGND VGND VPWR VPWR c$220 s$221 sky130_fd_sc_hd__ha_1
XFILLER_102_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_51_2 pp_row51_6 pp_row51_7 pp_row51_8 VGND VGND VPWR VPWR c$370 s$371
+ sky130_fd_sc_hd__fa_1
XFILLER_56_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_952 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$906 net955 net397 net947 net663 VGND VGND VPWR VPWR t$4868 sky130_fd_sc_hd__a22o_1
XU$$917 t$4873 net1318 VGND VGND VPWR VPWR booth_b12_m44 sky130_fd_sc_hd__xor2_1
XFILLER_141_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$928 net1679 net395 net1654 net661 VGND VGND VPWR VPWR t$4879 sky130_fd_sc_hd__a22o_1
Xdadda_fa_1_44_1 pp_row44_3 pp_row44_4 pp_row44_5 VGND VGND VPWR VPWR c$266 s$267
+ sky130_fd_sc_hd__fa_1
XFILLER_55_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$939 t$4884 net1318 VGND VGND VPWR VPWR booth_b12_m55 sky130_fd_sc_hd__xor2_1
XFILLER_141_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_21_0 pp_row21_11 c$1998 c$2000 VGND VGND VPWR VPWR c$2816 s$2817 sky130_fd_sc_hd__fa_1
Xdadda_fa_1_37_0 pp_row37_0 pp_row37_1 pp_row37_2 VGND VGND VPWR VPWR c$212 s$213
+ sky130_fd_sc_hd__fa_2
XFILLER_43_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1080 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_144_clk clknet_5_25__leaf_clk VGND VGND VPWR VPWR clknet_leaf_144_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_19_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1097 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_702 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_73_3 s$1607 s$1609 s$1611 VGND VGND VPWR VPWR c$2428 s$2429 sky130_fd_sc_hd__fa_1
XFILLER_121_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1201 net1202 VGND VGND VPWR VPWR net1201 sky130_fd_sc_hd__buf_4
XFILLER_182_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1212 net1213 VGND VGND VPWR VPWR net1212 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_3_66_2 c$1516 s$1519 s$1521 VGND VGND VPWR VPWR c$2370 s$2371 sky130_fd_sc_hd__fa_1
Xfanout1223 net66 VGND VGND VPWR VPWR net1223 sky130_fd_sc_hd__clkbuf_8
Xfanout1234 net65 VGND VGND VPWR VPWR net1234 sky130_fd_sc_hd__clkbuf_8
Xfanout1245 net1253 VGND VGND VPWR VPWR net1245 sky130_fd_sc_hd__buf_6
XFILLER_182_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1256 net1257 VGND VGND VPWR VPWR net1256 sky130_fd_sc_hd__buf_6
Xdadda_fa_3_59_1 c$1426 c$1428 c$1430 VGND VGND VPWR VPWR c$2312 s$2313 sky130_fd_sc_hd__fa_1
Xfanout1267 net1268 VGND VGND VPWR VPWR net1267 sky130_fd_sc_hd__buf_4
Xfanout1278 net1281 VGND VGND VPWR VPWR net1278 sky130_fd_sc_hd__buf_4
Xdadda_fa_6_36_0 c$3536 c$3538 s$3541 VGND VGND VPWR VPWR c$3968 s$3969 sky130_fd_sc_hd__fa_1
Xfanout1289 net1290 VGND VGND VPWR VPWR net1289 sky130_fd_sc_hd__buf_6
XFILLER_8_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3003 net1585 net524 net1558 net797 VGND VGND VPWR VPWR t$5939 sky130_fd_sc_hd__a22o_1
XU$$3014 net1369 VGND VGND VPWR VPWR notblock$5945\[0\] sky130_fd_sc_hd__inv_1
XU$$3025 t$5951 net1358 VGND VGND VPWR VPWR booth_b44_m2 sky130_fd_sc_hd__xor2_1
XU$$3036 net1516 net514 net1509 net787 VGND VGND VPWR VPWR t$5957 sky130_fd_sc_hd__a22o_1
XFILLER_47_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2302 net1647 net574 net1639 net847 VGND VGND VPWR VPWR t$5581 sky130_fd_sc_hd__a22o_1
XFILLER_46_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3047 t$5962 net1363 VGND VGND VPWR VPWR booth_b44_m13 sky130_fd_sc_hd__xor2_1
XU$$2313 t$5586 net1436 VGND VGND VPWR VPWR booth_b32_m57 sky130_fd_sc_hd__xor2_1
XU$$3058 net1142 net513 net1135 net786 VGND VGND VPWR VPWR t$5968 sky130_fd_sc_hd__a22o_1
XU$$2324 net1542 net575 net1534 net848 VGND VGND VPWR VPWR t$5592 sky130_fd_sc_hd__a22o_1
XU$$3069 t$5973 net1363 VGND VGND VPWR VPWR booth_b44_m24 sky130_fd_sc_hd__xor2_1
XU$$2335 net1775 net563 net1230 net836 VGND VGND VPWR VPWR t$5599 sky130_fd_sc_hd__a22o_1
XFILLER_34_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2346 t$5604 net1420 VGND VGND VPWR VPWR booth_b34_m5 sky130_fd_sc_hd__xor2_1
XFILLER_90_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1601 net1733 net615 net1724 net888 VGND VGND VPWR VPWR t$5223 sky130_fd_sc_hd__a22o_1
XU$$1612 t$5228 net1483 VGND VGND VPWR VPWR booth_b22_m49 sky130_fd_sc_hd__xor2_1
XU$$2357 net1220 net560 net1213 net833 VGND VGND VPWR VPWR t$5610 sky130_fd_sc_hd__a22o_1
XU$$1623 net1621 net616 net1614 net889 VGND VGND VPWR VPWR t$5234 sky130_fd_sc_hd__a22o_1
XU$$2368 t$5615 net1423 VGND VGND VPWR VPWR booth_b34_m16 sky130_fd_sc_hd__xor2_1
XU$$2379 net1109 net564 net1101 net837 VGND VGND VPWR VPWR t$5621 sky130_fd_sc_hd__a22o_1
XU$$1634 t$5239 net1481 VGND VGND VPWR VPWR booth_b22_m60 sky130_fd_sc_hd__xor2_1
XU$$1645 net17 VGND VGND VPWR VPWR notblock$5245\[1\] sky130_fd_sc_hd__inv_1
XU$$1656 net1031 net602 net932 net875 VGND VGND VPWR VPWR t$5252 sky130_fd_sc_hd__a22o_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1667 t$5257 net1469 VGND VGND VPWR VPWR booth_b24_m8 sky130_fd_sc_hd__xor2_1
X_1920_ clknet_leaf_81_clk booth_b8_m45 VGND VGND VPWR VPWR pp_row53_4 sky130_fd_sc_hd__dfxtp_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1678 net1194 net605 net1175 net878 VGND VGND VPWR VPWR t$5263 sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_135_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_135_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1689 t$5268 net1466 VGND VGND VPWR VPWR booth_b24_m19 sky130_fd_sc_hd__xor2_1
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1851_ clknet_leaf_25_clk booth_b50_m0 VGND VGND VPWR VPWR pp_row50_25 sky130_fd_sc_hd__dfxtp_1
XFILLER_175_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0802_ clknet_leaf_94_clk booth_b44_m47 VGND VGND VPWR VPWR pp_row91_9 sky130_fd_sc_hd__dfxtp_1
X_1782_ clknet_leaf_222_clk booth_b34_m14 VGND VGND VPWR VPWR pp_row48_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_129_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_109_0 s$3835 c$4112 s$4115 VGND VGND VPWR VPWR c$4370 s$4371 sky130_fd_sc_hd__fa_1
X_0733_ clknet_leaf_132_clk booth_b58_m60 VGND VGND VPWR VPWR pp_row118_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_116_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0664_ clknet_leaf_169_clk booth_b60_m25 VGND VGND VPWR VPWR pp_row85_20 sky130_fd_sc_hd__dfxtp_1
XFILLER_115_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2403_ clknet_leaf_127_clk booth_b60_m51 VGND VGND VPWR VPWR pp_row111_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_112_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0595_ clknet_leaf_193_clk booth_b32_m51 VGND VGND VPWR VPWR pp_row83_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2334_ clknet_leaf_86_clk booth_b2_m63 VGND VGND VPWR VPWR pp_row65_1 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_61_1 c$532 c$534 c$536 VGND VGND VPWR VPWR c$1460 s$1461 sky130_fd_sc_hd__fa_1
XFILLER_29_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$308 final_adder.p_new$310 final_adder.p_new$308 VGND VGND VPWR VPWR
+ final_adder.p_new$436 sky130_fd_sc_hd__and2_1
XFILLER_57_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2265_ clknet_leaf_230_clk booth_b10_m53 VGND VGND VPWR VPWR pp_row63_5 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$319 final_adder.p_new$318 final_adder.g_new$321 final_adder.g_new$319
+ VGND VGND VPWR VPWR final_adder.g_new$447 sky130_fd_sc_hd__a21o_1
Xdadda_fa_2_54_0 s$7 c$402 c$404 VGND VGND VPWR VPWR c$1374 s$1375 sky130_fd_sc_hd__fa_1
XFILLER_37_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1216_ clknet_leaf_143_clk booth_b46_m57 VGND VGND VPWR VPWR pp_row103_4 sky130_fd_sc_hd__dfxtp_1
XU$$4260 t$6582 net1259 VGND VGND VPWR VPWR booth_b62_m3 sky130_fd_sc_hd__xor2_1
X_2196_ clknet_leaf_223_clk booth_b16_m45 VGND VGND VPWR VPWR pp_row61_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_38_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4271 net1507 net418 net1498 net700 VGND VGND VPWR VPWR t$6588 sky130_fd_sc_hd__a22o_1
XU$$4282 t$6593 net1254 VGND VGND VPWR VPWR booth_b62_m14 sky130_fd_sc_hd__xor2_1
XFILLER_65_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4293 net1135 net419 net1119 net701 VGND VGND VPWR VPWR t$6599 sky130_fd_sc_hd__a22o_1
X_1147_ clknet_leaf_15_clk booth_b2_m16 VGND VGND VPWR VPWR pp_row18_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3570 net1233 net480 net1129 net753 VGND VGND VPWR VPWR t$6230 sky130_fd_sc_hd__a22o_1
XU$$3559_1794 VGND VGND VPWR VPWR U$$3559_1794/HI net1794 sky130_fd_sc_hd__conb_1
XFILLER_77_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3581 t$6235 net1325 VGND VGND VPWR VPWR booth_b52_m6 sky130_fd_sc_hd__xor2_1
XU$$3592 net1217 net480 net1208 net753 VGND VGND VPWR VPWR t$6241 sky130_fd_sc_hd__a22o_1
X_1078_ clknet_leaf_52_clk booth_b4_m7 VGND VGND VPWR VPWR pp_row11_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_8_0 pp_row8_2 pp_row8_3 pp_row8_4 VGND VGND VPWR VPWR c$3428 s$3429 sky130_fd_sc_hd__fa_1
XU$$2880 net1369 notblock$5875\[1\] VGND VGND VPWR VPWR t$5876 sky130_fd_sc_hd__and2_1
XFILLER_52_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2891 net935 net520 net1673 net793 VGND VGND VPWR VPWR t$5883 sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_126_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_126_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_178_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_83_2 s$2505 s$2507 s$2509 VGND VGND VPWR VPWR c$3192 s$3193 sky130_fd_sc_hd__fa_1
XFILLER_146_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_76_1 c$2442 c$2444 s$2447 VGND VGND VPWR VPWR c$3148 s$3149 sky130_fd_sc_hd__fa_1
XFILLER_136_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_53_0 s$3611 c$4000 s$4003 VGND VGND VPWR VPWR c$4258 s$4259 sky130_fd_sc_hd__fa_1
Xdadda_fa_4_69_0 s$1565 c$2382 c$2384 VGND VGND VPWR VPWR c$3104 s$3105 sky130_fd_sc_hd__fa_1
XFILLER_0_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_876 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$831 final_adder.p_new$846 final_adder.g_new$509 final_adder.g_new$847
+ VGND VGND VPWR VPWR final_adder.g_new$959 sky130_fd_sc_hd__a21o_2
Xfinal_adder.U$$853 final_adder.p_new$884 final_adder.g_new$949 final_adder.g_new$885
+ VGND VGND VPWR VPWR final_adder.g_new$981 sky130_fd_sc_hd__a21o_1
XFILLER_91_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$703 net1561 net402 net1522 net668 VGND VGND VPWR VPWR t$4765 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$875 final_adder.p_new$906 final_adder.g_new$859 final_adder.g_new$907
+ VGND VGND VPWR VPWR final_adder.g_new$1003 sky130_fd_sc_hd__a21o_1
XFILLER_21_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$714 t$4770 net1414 VGND VGND VPWR VPWR booth_b10_m11 sky130_fd_sc_hd__xor2_1
XU$$725 net1155 net401 net1146 net667 VGND VGND VPWR VPWR t$4776 sky130_fd_sc_hd__a22o_1
XFILLER_44_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$897 final_adder.p_new$928 final_adder.g_new$383 final_adder.g_new$929
+ VGND VGND VPWR VPWR final_adder.g_new$1025 sky130_fd_sc_hd__a21o_1
XU$$736 t$4781 net1413 VGND VGND VPWR VPWR booth_b10_m22 sky130_fd_sc_hd__xor2_1
XFILLER_44_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$747 net1056 net406 net1048 net672 VGND VGND VPWR VPWR t$4787 sky130_fd_sc_hd__a22o_1
XFILLER_16_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$758 t$4792 net1413 VGND VGND VPWR VPWR booth_b10_m33 sky130_fd_sc_hd__xor2_1
XU$$769 net949 net403 net941 net669 VGND VGND VPWR VPWR t$4798 sky130_fd_sc_hd__a22o_1
XFILLER_189_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_117_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_117_clk
+ sky130_fd_sc_hd__clkbuf_16
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_1132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_8 final_adder.g_new$855 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_71_0 s$743 c$1566 c$1568 VGND VGND VPWR VPWR c$2406 s$2407 sky130_fd_sc_hd__fa_1
XFILLER_3_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0380_ clknet_leaf_204_clk booth_b12_m64 VGND VGND VPWR VPWR pp_row76_1 sky130_fd_sc_hd__dfxtp_1
Xfanout1020 net1021 VGND VGND VPWR VPWR net1020 sky130_fd_sc_hd__buf_4
Xfanout1031 net1033 VGND VGND VPWR VPWR net1031 sky130_fd_sc_hd__clkbuf_4
Xfanout1042 net1046 VGND VGND VPWR VPWR net1042 sky130_fd_sc_hd__buf_6
XFILLER_67_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1053 net1054 VGND VGND VPWR VPWR net1053 sky130_fd_sc_hd__buf_6
Xfanout1064 net83 VGND VGND VPWR VPWR net1064 sky130_fd_sc_hd__buf_4
XFILLER_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1075 net1079 VGND VGND VPWR VPWR net1075 sky130_fd_sc_hd__buf_4
XFILLER_120_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1086 net1087 VGND VGND VPWR VPWR net1086 sky130_fd_sc_hd__buf_4
XFILLER_120_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1097 net1099 VGND VGND VPWR VPWR net1097 sky130_fd_sc_hd__buf_4
X_2050_ clknet_leaf_38_clk booth_b6_m51 VGND VGND VPWR VPWR pp_row57_3 sky130_fd_sc_hd__dfxtp_1
X_1001_ clknet_leaf_119_clk booth_b42_m59 VGND VGND VPWR VPWR pp_row101_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_75_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2110 t$5483 net1442 VGND VGND VPWR VPWR booth_b30_m24 sky130_fd_sc_hd__xor2_1
XFILLER_63_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_100_0 s$1933 c$2630 c$2632 VGND VGND VPWR VPWR c$3290 s$3291 sky130_fd_sc_hd__fa_1
XU$$2121 net1040 net577 net1024 net850 VGND VGND VPWR VPWR t$5489 sky130_fd_sc_hd__a22o_1
XU$$2132 t$5494 net1442 VGND VGND VPWR VPWR booth_b30_m35 sky130_fd_sc_hd__xor2_1
XFILLER_90_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2143 net926 net579 net1748 net852 VGND VGND VPWR VPWR t$5500 sky130_fd_sc_hd__a22o_1
XU$$2154 t$5505 net1445 VGND VGND VPWR VPWR booth_b30_m46 sky130_fd_sc_hd__xor2_1
XU$$2165 net1647 net578 net1639 net851 VGND VGND VPWR VPWR t$5511 sky130_fd_sc_hd__a22o_1
XU$$1420 net1107 net628 net1098 net901 VGND VGND VPWR VPWR t$5131 sky130_fd_sc_hd__a22o_1
XU$$2176 t$5516 net1444 VGND VGND VPWR VPWR booth_b30_m57 sky130_fd_sc_hd__xor2_1
XU$$1431 t$5136 net1486 VGND VGND VPWR VPWR booth_b20_m27 sky130_fd_sc_hd__xor2_1
XU$$1442 net1000 net630 net992 net903 VGND VGND VPWR VPWR t$5142 sky130_fd_sc_hd__a22o_1
XFILLER_62_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2187 net1539 net582 net1531 net855 VGND VGND VPWR VPWR t$5522 sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_108_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_108_clk
+ sky130_fd_sc_hd__clkbuf_16
XU$$2198 net1773 net571 net1230 net844 VGND VGND VPWR VPWR t$5529 sky130_fd_sc_hd__a22o_1
XU$$1453 t$5147 net1489 VGND VGND VPWR VPWR booth_b20_m38 sky130_fd_sc_hd__xor2_1
XFILLER_96_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1464 net1733 net634 net1724 net907 VGND VGND VPWR VPWR t$5153 sky130_fd_sc_hd__a22o_1
XU$$1475 t$5158 net1493 VGND VGND VPWR VPWR booth_b20_m49 sky130_fd_sc_hd__xor2_1
XFILLER_176_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1486 net1620 net632 net1612 net905 VGND VGND VPWR VPWR t$5164 sky130_fd_sc_hd__a22o_1
X_1903_ clknet_leaf_71_clk booth_b36_m16 VGND VGND VPWR VPWR pp_row52_18 sky130_fd_sc_hd__dfxtp_1
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1497 t$5169 net1493 VGND VGND VPWR VPWR booth_b20_m60 sky130_fd_sc_hd__xor2_1
XFILLER_187_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1834_ clknet_leaf_18_clk booth_b22_m28 VGND VGND VPWR VPWR pp_row50_11 sky130_fd_sc_hd__dfxtp_1
XU$$2463_1776 VGND VGND VPWR VPWR U$$2463_1776/HI net1776 sky130_fd_sc_hd__conb_1
Xdadda_fa_5_93_1 s$3249 s$3251 s$3253 VGND VGND VPWR VPWR c$3770 s$3771 sky130_fd_sc_hd__fa_1
XFILLER_175_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1765_ clknet_leaf_234_clk booth_b2_m46 VGND VGND VPWR VPWR pp_row48_1 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_86_0 c$3200 c$3202 c$3204 VGND VGND VPWR VPWR c$3740 s$3741 sky130_fd_sc_hd__fa_1
X_0716_ clknet_leaf_165_clk booth_b62_m25 VGND VGND VPWR VPWR pp_row87_20 sky130_fd_sc_hd__dfxtp_1
XFILLER_116_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1696_ clknet_leaf_18_clk booth_b28_m17 VGND VGND VPWR VPWR pp_row45_14 sky130_fd_sc_hd__dfxtp_1
XU$$417_1806 VGND VGND VPWR VPWR U$$417_1806/HI net1806 sky130_fd_sc_hd__conb_1
X_0647_ clknet_leaf_183_clk booth_b28_m57 VGND VGND VPWR VPWR pp_row85_4 sky130_fd_sc_hd__dfxtp_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_78_7 pp_row78_23 pp_row78_24 pp_row78_25 VGND VGND VPWR VPWR c$866 s$867
+ sky130_fd_sc_hd__fa_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0578_ clknet_leaf_189_clk booth_b50_m32 VGND VGND VPWR VPWR pp_row82_17 sky130_fd_sc_hd__dfxtp_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2317_ clknet_leaf_96_clk booth_b36_m28 VGND VGND VPWR VPWR pp_row64_18 sky130_fd_sc_hd__dfxtp_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$105 c$4360 s$4363 VGND VGND VPWR VPWR final_adder.$signal$212 final_adder.$signal$1195
+ sky130_fd_sc_hd__ha_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$116 c$4382 s$4385 VGND VGND VPWR VPWR final_adder.$signal$234 final_adder.$signal$1206
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$127 c$4404 s$4407 VGND VGND VPWR VPWR final_adder.U$$127/COUT final_adder.$signal$1217
+ sky130_fd_sc_hd__ha_2
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$138 final_adder.$signal$1206 final_adder.$signal$1207 VGND VGND VPWR
+ VPWR final_adder.p_new$266 sky130_fd_sc_hd__and2_1
XTAP_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$149 final_adder.$signal$1197 final_adder.$signal$214 final_adder.$signal$216
+ VGND VGND VPWR VPWR final_adder.g_new$277 sky130_fd_sc_hd__a21o_1
XFILLER_57_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2248_ clknet_leaf_149_clk booth_b48_m14 VGND VGND VPWR VPWR pp_row62_24 sky130_fd_sc_hd__dfxtp_1
XFILLER_122_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_409 net1732 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2179_ clknet_leaf_218_clk booth_b52_m8 VGND VGND VPWR VPWR pp_row60_26 sky130_fd_sc_hd__dfxtp_1
XU$$4090 t$6494 net1288 VGND VGND VPWR VPWR booth_b58_m55 sky130_fd_sc_hd__xor2_1
XFILLER_80_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_102_2 c$1936 c$1938 c$1940 VGND VGND VPWR VPWR c$2658 s$2659 sky130_fd_sc_hd__fa_1
XFILLER_135_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput101 b[42] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__buf_4
XFILLER_1_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput112 b[52] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__buf_4
XFILLER_49_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput123 b[62] VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__buf_4
XFILLER_163_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput134 c[104] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput145 c[114] VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_1
XFILLER_163_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_66_5 pp_row66_15 pp_row66_16 pp_row66_17 VGND VGND VPWR VPWR c$118 s$119
+ sky130_fd_sc_hd__fa_2
Xinput156 c[124] VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_1
XFILLER_56_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput167 c[19] VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_6_116_0 c$3856 c$3858 s$3861 VGND VGND VPWR VPWR c$4128 s$4129 sky130_fd_sc_hd__fa_1
Xinput178 c[29] VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_1
XTAP_3910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput189 c[39] VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_719 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$650 final_adder.p_new$674 final_adder.p_new$658 VGND VGND VPWR VPWR
+ final_adder.p_new$778 sky130_fd_sc_hd__and2_1
XFILLER_5_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$500 t$4660 net1244 VGND VGND VPWR VPWR booth_b6_m41 sky130_fd_sc_hd__xor2_1
XFILLER_45_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$661 final_adder.p_new$668 final_adder.g_new$685 final_adder.g_new$669
+ VGND VGND VPWR VPWR final_adder.g_new$789 sky130_fd_sc_hd__a21o_1
XTAP_3943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$672 final_adder.p_new$696 final_adder.p_new$680 VGND VGND VPWR VPWR
+ final_adder.p_new$800 sky130_fd_sc_hd__and2_1
XFILLER_63_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$511 net1707 net430 net1699 net712 VGND VGND VPWR VPWR t$4666 sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_36_3 s$1163 s$1165 s$1167 VGND VGND VPWR VPWR c$2132 s$2133 sky130_fd_sc_hd__fa_1
XTAP_3954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$683 final_adder.p_new$690 final_adder.g_new$707 final_adder.g_new$691
+ VGND VGND VPWR VPWR final_adder.g_new$811 sky130_fd_sc_hd__a21o_1
XFILLER_5_1096 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$522 t$4671 net1251 VGND VGND VPWR VPWR booth_b6_m52 sky130_fd_sc_hd__xor2_1
XTAP_3965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$533 net1595 net428 net1586 net710 VGND VGND VPWR VPWR t$4677 sky130_fd_sc_hd__a22o_1
XFILLER_44_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$694 final_adder.p_new$718 final_adder.p_new$702 VGND VGND VPWR VPWR
+ final_adder.p_new$822 sky130_fd_sc_hd__and2_1
XTAP_3976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$544 t$4682 net1251 VGND VGND VPWR VPWR booth_b6_m63 sky130_fd_sc_hd__xor2_1
XTAP_3987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$555 t$4689 net1239 VGND VGND VPWR VPWR booth_b8_m0 sky130_fd_sc_hd__xor2_1
XTAP_3998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_29_2 c$1076 c$1078 c$1080 VGND VGND VPWR VPWR c$2074 s$2075 sky130_fd_sc_hd__fa_1
XU$$566 net1561 net415 net1521 net681 VGND VGND VPWR VPWR t$4695 sky130_fd_sc_hd__a22o_1
XFILLER_186_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$577 t$4700 net1239 VGND VGND VPWR VPWR booth_b8_m11 sky130_fd_sc_hd__xor2_1
XU$$588 net1155 net410 net1146 net676 VGND VGND VPWR VPWR t$4706 sky130_fd_sc_hd__a22o_1
XFILLER_112_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$599 t$4711 net1235 VGND VGND VPWR VPWR booth_b8_m22 sky130_fd_sc_hd__xor2_1
XFILLER_72_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1550_ clknet_leaf_121_clk booth_b50_m55 VGND VGND VPWR VPWR pp_row105_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_193_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0501_ clknet_leaf_208_clk booth_b64_m15 VGND VGND VPWR VPWR pp_row79_25 sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1481_ clknet_leaf_246_clk booth_b2_m35 VGND VGND VPWR VPWR pp_row37_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_113_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0432_ clknet_leaf_154_clk booth_b50_m27 VGND VGND VPWR VPWR pp_row77_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_79_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0363_ clknet_leaf_204_clk booth_b38_m37 VGND VGND VPWR VPWR pp_row75_14 sky130_fd_sc_hd__dfxtp_1
X_2102_ clknet_leaf_29_clk booth_b40_m18 VGND VGND VPWR VPWR pp_row58_20 sky130_fd_sc_hd__dfxtp_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0294_ clknet_leaf_199_clk booth_b28_m45 VGND VGND VPWR VPWR pp_row73_10 sky130_fd_sc_hd__dfxtp_1
X_2033_ clknet_leaf_72_clk booth_b38_m18 VGND VGND VPWR VPWR pp_row56_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_35_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_31_2 pp_row31_6 pp_row31_7 pp_row31_8 VGND VGND VPWR VPWR c$1104 s$1105
+ sky130_fd_sc_hd__fa_1
XFILLER_90_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1250 t$5044 net1664 VGND VGND VPWR VPWR booth_b18_m5 sky130_fd_sc_hd__xor2_1
XU$$1261 net1219 net635 net1210 net908 VGND VGND VPWR VPWR t$5050 sky130_fd_sc_hd__a22o_1
XFILLER_22_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1272 t$5055 net1665 VGND VGND VPWR VPWR booth_b18_m16 sky130_fd_sc_hd__xor2_1
XU$$1283 net1105 net635 net1097 net908 VGND VGND VPWR VPWR t$5061 sky130_fd_sc_hd__a22o_1
XFILLER_31_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1294 t$5066 net1663 VGND VGND VPWR VPWR booth_b18_m27 sky130_fd_sc_hd__xor2_1
XFILLER_176_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1817_ clknet_leaf_224_clk booth_b42_m7 VGND VGND VPWR VPWR pp_row49_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_117_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1748_ clknet_leaf_238_clk booth_b22_m25 VGND VGND VPWR VPWR pp_row47_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1679_ clknet_leaf_235_clk net195 VGND VGND VPWR VPWR pp_row44_24 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_83_5 pp_row83_15 pp_row83_16 pp_row83_17 VGND VGND VPWR VPWR c$948 s$949
+ sky130_fd_sc_hd__fa_1
Xfanout802 net803 VGND VGND VPWR VPWR net802 sky130_fd_sc_hd__buf_4
XFILLER_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout813 net814 VGND VGND VPWR VPWR net813 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_76_4 pp_row76_17 pp_row76_18 pp_row76_19 VGND VGND VPWR VPWR c$824 s$825
+ sky130_fd_sc_hd__fa_1
Xfanout824 net826 VGND VGND VPWR VPWR net824 sky130_fd_sc_hd__buf_4
Xfanout835 net841 VGND VGND VPWR VPWR net835 sky130_fd_sc_hd__buf_4
XFILLER_86_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout846 net847 VGND VGND VPWR VPWR net846 sky130_fd_sc_hd__buf_4
Xfanout857 net859 VGND VGND VPWR VPWR net857 sky130_fd_sc_hd__buf_4
XFILLER_113_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_69_3 pp_row69_24 pp_row69_25 pp_row69_26 VGND VGND VPWR VPWR c$696 s$697
+ sky130_fd_sc_hd__fa_1
Xfanout868 net874 VGND VGND VPWR VPWR net868 sky130_fd_sc_hd__buf_2
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout879 sel_1$5248 VGND VGND VPWR VPWR net879 sky130_fd_sc_hd__buf_6
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_46_2 s$2209 s$2211 s$2213 VGND VGND VPWR VPWR c$2970 s$2971 sky130_fd_sc_hd__fa_1
XTAP_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_39_1 c$2146 c$2148 s$2151 VGND VGND VPWR VPWR c$2926 s$2927 sky130_fd_sc_hd__fa_1
XTAP_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_16_0 s$3463 c$3926 s$3929 VGND VGND VPWR VPWR c$4184 s$4185 sky130_fd_sc_hd__fa_2
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_206 net1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_217 net1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_228 net1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_239 net1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4407_1824 VGND VGND VPWR VPWR U$$4407_1824/HI net1824 sky130_fd_sc_hd__conb_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_ha_0_58_3 pp_row58_9 pp_row58_10 VGND VGND VPWR VPWR c$30 s$31 sky130_fd_sc_hd__ha_1
XFILLER_89_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_71_3 pp_row71_9 pp_row71_10 pp_row71_11 VGND VGND VPWR VPWR c$170 s$171
+ sky130_fd_sc_hd__fa_2
XFILLER_107_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_0_64_2 pp_row64_6 pp_row64_7 pp_row64_8 VGND VGND VPWR VPWR c$88 s$89 sky130_fd_sc_hd__fa_1
XFILLER_190_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_41_1 c$1210 c$1212 c$1214 VGND VGND VPWR VPWR c$2168 s$2169 sky130_fd_sc_hd__fa_1
XFILLER_190_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_0_57_1 pp_row57_3 pp_row57_4 pp_row57_5 VGND VGND VPWR VPWR c$20 s$21 sky130_fd_sc_hd__fa_1
XTAP_3740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_34_0 s$205 c$1122 c$1124 VGND VGND VPWR VPWR c$2110 s$2111 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$480 final_adder.p_new$486 final_adder.p_new$482 VGND VGND VPWR VPWR
+ final_adder.p_new$608 sky130_fd_sc_hd__and2_1
XTAP_3762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$330 net1080 net527 net1071 net800 VGND VGND VPWR VPWR t$4574 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$491 final_adder.p_new$492 final_adder.g_new$497 final_adder.g_new$493
+ VGND VGND VPWR VPWR final_adder.g_new$619 sky130_fd_sc_hd__a21o_1
XFILLER_91_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$341 t$4579 net1278 VGND VGND VPWR VPWR booth_b4_m30 sky130_fd_sc_hd__xor2_1
XFILLER_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$352 net973 net527 net964 net800 VGND VGND VPWR VPWR t$4585 sky130_fd_sc_hd__a22o_1
XTAP_3795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$363 t$4590 net1276 VGND VGND VPWR VPWR booth_b4_m41 sky130_fd_sc_hd__xor2_1
XFILLER_83_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$374 net1706 net533 net1699 net806 VGND VGND VPWR VPWR t$4596 sky130_fd_sc_hd__a22o_1
XFILLER_45_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$385 t$4601 net1280 VGND VGND VPWR VPWR booth_b4_m52 sky130_fd_sc_hd__xor2_1
XFILLER_60_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$396 net1595 net529 net1586 net802 VGND VGND VPWR VPWR t$4607 sky130_fd_sc_hd__a22o_1
XFILLER_32_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0981_ clknet_leaf_114_clk booth_b38_m62 VGND VGND VPWR VPWR pp_row100_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1602_ clknet_leaf_243_clk booth_b4_m38 VGND VGND VPWR VPWR pp_row42_2 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_93_4 pp_row93_18 pp_row93_19 c$1032 VGND VGND VPWR VPWR c$1850 s$1851
+ sky130_fd_sc_hd__fa_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1533_ clknet_leaf_44_clk booth_b10_m29 VGND VGND VPWR VPWR pp_row39_5 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_86_3 c$970 c$972 c$974 VGND VGND VPWR VPWR c$1764 s$1765 sky130_fd_sc_hd__fa_1
XFILLER_141_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_79_2 c$862 c$864 c$866 VGND VGND VPWR VPWR c$1678 s$1679 sky130_fd_sc_hd__fa_1
X_1464_ clknet_leaf_40_clk booth_b12_m24 VGND VGND VPWR VPWR pp_row36_6 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_56_1 s$3027 s$3029 s$3031 VGND VGND VPWR VPWR c$3622 s$3623 sky130_fd_sc_hd__fa_1
XFILLER_86_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0415_ clknet_leaf_155_clk booth_b18_m59 VGND VGND VPWR VPWR pp_row77_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_68_844 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1395_ clknet_leaf_181_clk net159 VGND VGND VPWR VPWR pp_row127_2 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_49_0 c$2978 c$2980 c$2982 VGND VGND VPWR VPWR c$3592 s$3593 sky130_fd_sc_hd__fa_1
XFILLER_67_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0346_ clknet_leaf_203_clk booth_b64_m10 VGND VGND VPWR VPWR pp_row74_28 sky130_fd_sc_hd__dfxtp_1
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_2_23_0 pp_row23_0 pp_row23_1 VGND VGND VPWR VPWR c$1052 s$1053 sky130_fd_sc_hd__ha_1
XU$$3970_1800 VGND VGND VPWR VPWR U$$3970_1800/HI net1800 sky130_fd_sc_hd__conb_1
XFILLER_95_696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0277_ clknet_leaf_124_clk booth_b58_m55 VGND VGND VPWR VPWR pp_row113_5 sky130_fd_sc_hd__dfxtp_1
X_2016_ clknet_leaf_135_clk booth_b58_m50 VGND VGND VPWR VPWR pp_row108_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_35_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_102_1 pp_row102_3 pp_row102_4 pp_row102_5 VGND VGND VPWR VPWR c$1944 s$1945
+ sky130_fd_sc_hd__fa_1
XFILLER_168_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1080 t$4956 net1188 VGND VGND VPWR VPWR booth_b14_m57 sky130_fd_sc_hd__xor2_1
XU$$1091 net1535 net391 net1527 net657 VGND VGND VPWR VPWR t$4962 sky130_fd_sc_hd__a22o_1
XFILLER_50_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_123_0 pp_row123_0 pp_row123_1 pp_row123_2 VGND VGND VPWR VPWR c$3888 s$3889
+ sky130_fd_sc_hd__fa_1
Xclkbuf_leaf_30_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_177_996 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4437_1839 VGND VGND VPWR VPWR U$$4437_1839/HI net1839 sky130_fd_sc_hd__conb_1
XFILLER_2_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_81_2 pp_row81_6 pp_row81_7 pp_row81_8 VGND VGND VPWR VPWR c$910 s$911
+ sky130_fd_sc_hd__fa_1
Xfanout610 net612 VGND VGND VPWR VPWR net610 sky130_fd_sc_hd__buf_4
Xfanout1608 net1610 VGND VGND VPWR VPWR net1608 sky130_fd_sc_hd__buf_4
Xfanout621 net622 VGND VGND VPWR VPWR net621 sky130_fd_sc_hd__buf_4
Xfanout1619 net115 VGND VGND VPWR VPWR net1619 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_74_1 pp_row74_11 pp_row74_12 pp_row74_13 VGND VGND VPWR VPWR c$782 s$783
+ sky130_fd_sc_hd__fa_1
Xfanout632 net634 VGND VGND VPWR VPWR net632 sky130_fd_sc_hd__buf_4
XFILLER_77_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout643 net644 VGND VGND VPWR VPWR net643 sky130_fd_sc_hd__buf_4
XFILLER_59_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout654 net655 VGND VGND VPWR VPWR net654 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_4_51_0 s$1349 c$2238 c$2240 VGND VGND VPWR VPWR c$2996 s$2997 sky130_fd_sc_hd__fa_1
Xclkbuf_leaf_97_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_97_clk sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_1_67_0 pp_row67_18 pp_row67_19 pp_row67_20 VGND VGND VPWR VPWR c$654 s$655
+ sky130_fd_sc_hd__fa_1
Xfanout665 net666 VGND VGND VPWR VPWR net665 sky130_fd_sc_hd__clkbuf_8
Xfanout676 net678 VGND VGND VPWR VPWR net676 sky130_fd_sc_hd__buf_4
Xfanout687 net692 VGND VGND VPWR VPWR net687 sky130_fd_sc_hd__buf_4
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout698 net699 VGND VGND VPWR VPWR net698 sky130_fd_sc_hd__clkbuf_4
XTAP_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2709 net1681 net546 net1656 net819 VGND VGND VPWR VPWR t$5789 sky130_fd_sc_hd__a22o_1
XTAP_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_21_clk clknet_5_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_6_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_96_2 c$1876 s$1879 s$1881 VGND VGND VPWR VPWR c$2610 s$2611 sky130_fd_sc_hd__fa_1
XFILLER_136_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_1131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_89_1 c$1786 c$1788 c$1790 VGND VGND VPWR VPWR c$2552 s$2553 sky130_fd_sc_hd__fa_2
XFILLER_151_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_66_0 c$3656 c$3658 s$3661 VGND VGND VPWR VPWR c$4028 s$4029 sky130_fd_sc_hd__fa_1
XFILLER_150_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_749 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_88_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_88_clk sky130_fd_sc_hd__clkbuf_16
X_0200_ clknet_leaf_180_clk booth_b64_m48 VGND VGND VPWR VPWR pp_row112_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_65_803 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1180_ clknet_leaf_49_clk booth_b14_m6 VGND VGND VPWR VPWR pp_row20_7 sky130_fd_sc_hd__dfxtp_1
XU$$3900 net1052 net463 net1044 net736 VGND VGND VPWR VPWR t$6398 sky130_fd_sc_hd__a22o_1
XFILLER_77_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3911 t$6403 net1297 VGND VGND VPWR VPWR booth_b56_m34 sky130_fd_sc_hd__xor2_1
XTAP_4260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_118_1 pp_row118_3 pp_row118_4 pp_row118_5 VGND VGND VPWR VPWR c$3400 s$3401
+ sky130_fd_sc_hd__fa_1
XTAP_4271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3922 net945 net464 net929 net737 VGND VGND VPWR VPWR t$6409 sky130_fd_sc_hd__a22o_1
XU$$3933 t$6414 net1298 VGND VGND VPWR VPWR booth_b56_m45 sky130_fd_sc_hd__xor2_1
XU$$3696_1796 VGND VGND VPWR VPWR U$$3696_1796/HI net1796 sky130_fd_sc_hd__conb_1
XTAP_4282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3944 net1659 net462 net1651 net735 VGND VGND VPWR VPWR t$6420 sky130_fd_sc_hd__a22o_1
XTAP_4293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3955 t$6425 net1297 VGND VGND VPWR VPWR booth_b56_m56 sky130_fd_sc_hd__xor2_1
XU$$3966 net1549 net462 net1541 net735 VGND VGND VPWR VPWR t$6431 sky130_fd_sc_hd__a22o_1
XTAP_3570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3977 notblock$6435\[2\] net54 net1292 t$6436 notblock$6435\[0\] VGND VGND VPWR
+ VPWR sel_0$6437 sky130_fd_sc_hd__a32o_1
XU$$3988 t$6443 net1283 VGND VGND VPWR VPWR booth_b58_m4 sky130_fd_sc_hd__xor2_1
XU$$160 t$4487 net1389 VGND VGND VPWR VPWR booth_b2_m8 sky130_fd_sc_hd__xor2_1
XU$$3999 net1502 net455 net66 net728 VGND VGND VPWR VPWR t$6449 sky130_fd_sc_hd__a22o_1
XTAP_3592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$171 net1194 net620 net1175 net893 VGND VGND VPWR VPWR t$4493 sky130_fd_sc_hd__a22o_1
XU$$182 t$4498 net1389 VGND VGND VPWR VPWR booth_b2_m19 sky130_fd_sc_hd__xor2_1
XU$$193 net1080 net619 net1071 net892 VGND VGND VPWR VPWR t$4504 sky130_fd_sc_hd__a22o_1
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0964_ clknet_leaf_116_clk booth_b40_m59 VGND VGND VPWR VPWR pp_row99_3 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_12_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_174_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0895_ clknet_leaf_100_clk booth_b56_m39 VGND VGND VPWR VPWR pp_row95_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_91_1 pp_row91_12 pp_row91_13 pp_row91_14 VGND VGND VPWR VPWR c$1820 s$1821
+ sky130_fd_sc_hd__fa_1
Xdadda_fa_2_84_0 pp_row84_20 pp_row84_21 pp_row84_22 VGND VGND VPWR VPWR c$1734 s$1735
+ sky130_fd_sc_hd__fa_1
Xoutput257 net257 VGND VGND VPWR VPWR o[0] sky130_fd_sc_hd__buf_2
Xoutput268 net268 VGND VGND VPWR VPWR o[10] sky130_fd_sc_hd__buf_2
X_1516_ clknet_leaf_17_clk booth_b24_m14 VGND VGND VPWR VPWR pp_row38_12 sky130_fd_sc_hd__dfxtp_1
Xoutput279 net279 VGND VGND VPWR VPWR o[11] sky130_fd_sc_hd__buf_2
X_2496_ clknet_leaf_141_clk booth_b32_m37 VGND VGND VPWR VPWR pp_row69_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_142_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1447_ clknet_leaf_64_clk booth_b20_m15 VGND VGND VPWR VPWR pp_row35_10 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_79_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_79_clk sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_1_60_7 c$36 c$38 s$41 VGND VGND VPWR VPWR c$542 s$543 sky130_fd_sc_hd__fa_1
XFILLER_56_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1378_ clknet_leaf_43_clk booth_b12_m20 VGND VGND VPWR VPWR pp_row32_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_28_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_53_6 pp_row53_20 pp_row53_21 pp_row53_22 VGND VGND VPWR VPWR c$414 s$415
+ sky130_fd_sc_hd__fa_1
XFILLER_83_633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0329_ clknet_leaf_201_clk booth_b34_m40 VGND VGND VPWR VPWR pp_row74_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_95_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_46_5 pp_row46_15 pp_row46_16 pp_row46_17 VGND VGND VPWR VPWR c$298 s$299
+ sky130_fd_sc_hd__fa_1
XFILLER_167_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_7_5_0 s$3419 c$3904 s$3907 VGND VGND VPWR VPWR c$4162 s$4163 sky130_fd_sc_hd__fa_1
XFILLER_82_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_83_0 s$3731 c$4060 s$4063 VGND VGND VPWR VPWR c$4318 s$4319 sky130_fd_sc_hd__fa_2
XFILLER_87_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_99_0 s$1923 c$2622 c$2624 VGND VGND VPWR VPWR c$3284 s$3285 sky130_fd_sc_hd__fa_1
XFILLER_99_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1405 net1407 VGND VGND VPWR VPWR net1405 sky130_fd_sc_hd__buf_6
Xfanout1416 net3 VGND VGND VPWR VPWR net1416 sky130_fd_sc_hd__buf_6
XFILLER_132_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1427 net1429 VGND VGND VPWR VPWR net1427 sky130_fd_sc_hd__buf_6
Xfanout440 net441 VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__buf_4
Xfanout1438 net27 VGND VGND VPWR VPWR net1438 sky130_fd_sc_hd__buf_8
Xfanout1449 net1450 VGND VGND VPWR VPWR net1449 sky130_fd_sc_hd__buf_4
Xfanout451 net459 VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__buf_4
Xfanout462 net463 VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__buf_4
Xfanout473 net475 VGND VGND VPWR VPWR net473 sky130_fd_sc_hd__buf_4
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout484 net487 VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__buf_4
XFILLER_171_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout495 net496 VGND VGND VPWR VPWR net495 sky130_fd_sc_hd__clkbuf_8
XU$$3207 net1086 net502 net1076 net775 VGND VGND VPWR VPWR t$6044 sky130_fd_sc_hd__a22o_1
XU$$3218 t$6049 net1351 VGND VGND VPWR VPWR booth_b46_m30 sky130_fd_sc_hd__xor2_1
XFILLER_24_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3229 net975 net503 net966 net776 VGND VGND VPWR VPWR t$6055 sky130_fd_sc_hd__a22o_1
XU$$2506 net1162 net554 net1150 net827 VGND VGND VPWR VPWR t$5686 sky130_fd_sc_hd__a22o_1
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2517 t$5691 net1404 VGND VGND VPWR VPWR booth_b36_m22 sky130_fd_sc_hd__xor2_1
XFILLER_104_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2528 net1058 net554 net1050 net827 VGND VGND VPWR VPWR t$5697 sky130_fd_sc_hd__a22o_1
XU$$2539 t$5702 net1410 VGND VGND VPWR VPWR booth_b36_m33 sky130_fd_sc_hd__xor2_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1805 net1509 net597 net1500 net870 VGND VGND VPWR VPWR t$5328 sky130_fd_sc_hd__a22o_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1816 t$5333 net1458 VGND VGND VPWR VPWR booth_b26_m14 sky130_fd_sc_hd__xor2_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1827 net1132 net594 net1116 net867 VGND VGND VPWR VPWR t$5339 sky130_fd_sc_hd__a22o_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1838 t$5344 net1461 VGND VGND VPWR VPWR booth_b26_m25 sky130_fd_sc_hd__xor2_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1849 net1025 net596 net1017 net869 VGND VGND VPWR VPWR t$5350 sky130_fd_sc_hd__a22o_1
XFILLER_9_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4459_1850 VGND VGND VPWR VPWR U$$4459_1850/HI net1850 sky130_fd_sc_hd__conb_1
XFILLER_128_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0680_ clknet_leaf_180_clk booth_b42_m44 VGND VGND VPWR VPWR pp_row86_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2350_ clknet_leaf_77_clk booth_b30_m35 VGND VGND VPWR VPWR pp_row65_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_69_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1301_ clknet_leaf_250_clk booth_b8_m20 VGND VGND VPWR VPWR pp_row28_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_123_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2281_ clknet_leaf_153_clk booth_b40_m23 VGND VGND VPWR VPWR pp_row63_20 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_63_5 s$593 s$595 s$597 VGND VGND VPWR VPWR c$1492 s$1493 sky130_fd_sc_hd__fa_2
X_1232_ clknet_leaf_12_clk booth_b4_m20 VGND VGND VPWR VPWR pp_row24_2 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_1_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_56_4 s$461 s$463 s$465 VGND VGND VPWR VPWR c$1406 s$1407 sky130_fd_sc_hd__fa_1
XU$$4420 net1177 sel_0$6647 net1168 net694 VGND VGND VPWR VPWR t$6664 sky130_fd_sc_hd__a22o_1
XU$$4431 t$6669 net1836 VGND VGND VPWR VPWR booth_b64_m20 sky130_fd_sc_hd__xor2_1
XFILLER_77_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4442 net1078 sel_0$6647 net1070 net698 VGND VGND VPWR VPWR t$6675 sky130_fd_sc_hd__a22o_1
XU$$4453 t$6680 net1847 VGND VGND VPWR VPWR booth_b64_m31 sky130_fd_sc_hd__xor2_1
X_1163_ clknet_leaf_50_clk booth_b6_m13 VGND VGND VPWR VPWR pp_row19_3 sky130_fd_sc_hd__dfxtp_1
XU$$4464 net971 sel_0$6647 net963 net699 VGND VGND VPWR VPWR t$6686 sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_49_3 c$328 c$330 s$333 VGND VGND VPWR VPWR c$1320 s$1321 sky130_fd_sc_hd__fa_1
XU$$3730 t$6311 net1304 VGND VGND VPWR VPWR booth_b54_m12 sky130_fd_sc_hd__xor2_1
XU$$4475 t$6691 net1858 VGND VGND VPWR VPWR booth_b64_m42 sky130_fd_sc_hd__xor2_1
XTAP_4090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4486 net1696 sel_0$6647 net1688 net693 VGND VGND VPWR VPWR t$6697 sky130_fd_sc_hd__a22o_1
XU$$3741 net1151 net468 net1141 net741 VGND VGND VPWR VPWR t$6317 sky130_fd_sc_hd__a22o_1
XU$$3752 t$6322 net1301 VGND VGND VPWR VPWR booth_b54_m23 sky130_fd_sc_hd__xor2_1
XU$$4497 t$6702 net1869 VGND VGND VPWR VPWR booth_b64_m53 sky130_fd_sc_hd__xor2_1
X_1094_ clknet_leaf_121_clk booth_b54_m48 VGND VGND VPWR VPWR pp_row102_9 sky130_fd_sc_hd__dfxtp_1
XU$$3763 net1052 net469 net1044 net742 VGND VGND VPWR VPWR t$6328 sky130_fd_sc_hd__a22o_1
XFILLER_64_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3774 t$6333 net1301 VGND VGND VPWR VPWR booth_b54_m34 sky130_fd_sc_hd__xor2_1
XU$$3785 net946 net472 net930 net745 VGND VGND VPWR VPWR t$6339 sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_19_1 s$2805 s$2807 s$2809 VGND VGND VPWR VPWR c$3474 s$3475 sky130_fd_sc_hd__fa_1
XU$$3796 t$6344 net1307 VGND VGND VPWR VPWR booth_b54_m45 sky130_fd_sc_hd__xor2_1
XFILLER_100_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1996_ clknet_leaf_69_clk booth_b28_m27 VGND VGND VPWR VPWR pp_row55_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_193_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0947_ clknet_leaf_113_clk booth_b42_m56 VGND VGND VPWR VPWR pp_row98_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_162_903 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0878_ clknet_leaf_93_clk booth_b62_m32 VGND VGND VPWR VPWR pp_row94_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_133_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2479_ clknet_leaf_198_clk net221 VGND VGND VPWR VPWR pp_row68_32 sky130_fd_sc_hd__dfxtp_2
Xdadda_fa_1_51_3 pp_row51_9 pp_row51_10 pp_row51_11 VGND VGND VPWR VPWR c$372 s$373
+ sky130_fd_sc_hd__fa_1
XFILLER_84_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$907 t$4868 net1314 VGND VGND VPWR VPWR booth_b12_m39 sky130_fd_sc_hd__xor2_1
XU$$918 net1724 net398 net1715 net664 VGND VGND VPWR VPWR t$4874 sky130_fd_sc_hd__a22o_1
XU$$929 t$4879 net1317 VGND VGND VPWR VPWR booth_b12_m50 sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_44_2 pp_row44_6 pp_row44_7 pp_row44_8 VGND VGND VPWR VPWR c$268 s$269
+ sky130_fd_sc_hd__fa_1
XFILLER_141_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_21_1 c$2002 c$2004 s$2007 VGND VGND VPWR VPWR c$2818 s$2819 sky130_fd_sc_hd__fa_1
XFILLER_58_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_14_0 pp_row14_2 pp_row14_3 pp_row14_4 VGND VGND VPWR VPWR c$2774 s$2775
+ sky130_fd_sc_hd__fa_1
XFILLER_145_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_29__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_5_29__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_79_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1202 net1209 VGND VGND VPWR VPWR net1202 sky130_fd_sc_hd__buf_4
XFILLER_67_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1213 net1215 VGND VGND VPWR VPWR net1213 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_3_66_3 s$1523 s$1525 s$1527 VGND VGND VPWR VPWR c$2372 s$2373 sky130_fd_sc_hd__fa_1
XFILLER_182_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1224 net1226 VGND VGND VPWR VPWR net1224 sky130_fd_sc_hd__buf_4
Xfanout1235 net64 VGND VGND VPWR VPWR net1235 sky130_fd_sc_hd__buf_6
Xfanout1246 net1247 VGND VGND VPWR VPWR net1246 sky130_fd_sc_hd__buf_4
XFILLER_121_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_59_2 c$1432 s$1435 s$1437 VGND VGND VPWR VPWR c$2314 s$2315 sky130_fd_sc_hd__fa_1
XFILLER_120_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1257 net1258 VGND VGND VPWR VPWR net1257 sky130_fd_sc_hd__buf_4
XU$$4489_1865 VGND VGND VPWR VPWR U$$4489_1865/HI net1865 sky130_fd_sc_hd__conb_1
Xfanout1268 net58 VGND VGND VPWR VPWR net1268 sky130_fd_sc_hd__buf_4
Xfanout1279 net1281 VGND VGND VPWR VPWR net1279 sky130_fd_sc_hd__buf_6
XFILLER_120_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3004 t$5939 net1374 VGND VGND VPWR VPWR booth_b42_m60 sky130_fd_sc_hd__xor2_1
XU$$3015 net39 VGND VGND VPWR VPWR notblock$5945\[1\] sky130_fd_sc_hd__inv_1
XFILLER_75_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_29_0 c$3508 c$3510 s$3513 VGND VGND VPWR VPWR c$3954 s$3955 sky130_fd_sc_hd__fa_1
XU$$3026 net1034 net510 net935 net783 VGND VGND VPWR VPWR t$5952 sky130_fd_sc_hd__a22o_1
XU$$3037 t$5957 net1362 VGND VGND VPWR VPWR booth_b44_m8 sky130_fd_sc_hd__xor2_1
XU$$2303 t$5581 net1435 VGND VGND VPWR VPWR booth_b32_m52 sky130_fd_sc_hd__xor2_1
XFILLER_75_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3048 net1196 net511 net1178 net784 VGND VGND VPWR VPWR t$5963 sky130_fd_sc_hd__a22o_1
XU$$3059 t$5968 net1360 VGND VGND VPWR VPWR booth_b44_m19 sky130_fd_sc_hd__xor2_1
XU$$2314 net1596 net573 net1587 net846 VGND VGND VPWR VPWR t$5587 sky130_fd_sc_hd__a22o_1
XU$$2325 t$5592 net1437 VGND VGND VPWR VPWR booth_b32_m63 sky130_fd_sc_hd__xor2_1
XU$$2336 t$5599 net1423 VGND VGND VPWR VPWR booth_b34_m0 sky130_fd_sc_hd__xor2_1
XU$$2347 net1561 net561 net1521 net834 VGND VGND VPWR VPWR t$5605 sky130_fd_sc_hd__a22o_1
XU$$1602 t$5223 net1480 VGND VGND VPWR VPWR booth_b22_m44 sky130_fd_sc_hd__xor2_1
XFILLER_34_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1613 net1681 net616 net1654 net889 VGND VGND VPWR VPWR t$5229 sky130_fd_sc_hd__a22o_1
XU$$2358 t$5610 net1420 VGND VGND VPWR VPWR booth_b34_m11 sky130_fd_sc_hd__xor2_1
XFILLER_188_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2369 net1162 net563 net1150 net836 VGND VGND VPWR VPWR t$5616 sky130_fd_sc_hd__a22o_1
XU$$1624 t$5234 net1483 VGND VGND VPWR VPWR booth_b22_m55 sky130_fd_sc_hd__xor2_1
XU$$1635 net1553 net617 net1544 net890 VGND VGND VPWR VPWR t$5240 sky130_fd_sc_hd__a22o_1
XU$$1646 net1471 VGND VGND VPWR VPWR notblock$5245\[2\] sky130_fd_sc_hd__inv_1
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1657 t$5252 net1466 VGND VGND VPWR VPWR booth_b24_m3 sky130_fd_sc_hd__xor2_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1668 net1509 net605 net1499 net878 VGND VGND VPWR VPWR t$5258 sky130_fd_sc_hd__a22o_1
XFILLER_43_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1679 t$5263 net1469 VGND VGND VPWR VPWR booth_b24_m14 sky130_fd_sc_hd__xor2_1
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1850_ clknet_leaf_135_clk booth_b52_m55 VGND VGND VPWR VPWR pp_row107_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_147_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0801_ clknet_leaf_139_clk booth_b42_m49 VGND VGND VPWR VPWR pp_row91_8 sky130_fd_sc_hd__dfxtp_1
X_1781_ clknet_leaf_222_clk booth_b32_m16 VGND VGND VPWR VPWR pp_row48_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_128_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0732_ clknet_leaf_163_clk booth_b46_m42 VGND VGND VPWR VPWR pp_row88_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_116_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0663_ clknet_leaf_172_clk booth_b58_m27 VGND VGND VPWR VPWR pp_row85_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_115_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2402_ clknet_leaf_99_clk booth_b58_m8 VGND VGND VPWR VPWR pp_row66_29 sky130_fd_sc_hd__dfxtp_1
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0594_ clknet_leaf_193_clk booth_b30_m53 VGND VGND VPWR VPWR pp_row83_6 sky130_fd_sc_hd__dfxtp_1
X_2333_ clknet_leaf_198_clk net217 VGND VGND VPWR VPWR pp_row64_33 sky130_fd_sc_hd__dfxtp_1
XFILLER_97_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_61_2 c$538 c$540 c$542 VGND VGND VPWR VPWR c$1462 s$1463 sky130_fd_sc_hd__fa_1
XFILLER_112_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2264_ clknet_leaf_230_clk booth_b8_m55 VGND VGND VPWR VPWR pp_row63_4 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$309 final_adder.p_new$308 final_adder.g_new$311 final_adder.g_new$309
+ VGND VGND VPWR VPWR final_adder.g_new$437 sky130_fd_sc_hd__a21o_1
XFILLER_112_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_54_1 c$406 c$408 c$410 VGND VGND VPWR VPWR c$1376 s$1377 sky130_fd_sc_hd__fa_1
X_1215_ clknet_leaf_47_clk booth_b0_m23 VGND VGND VPWR VPWR pp_row23_0 sky130_fd_sc_hd__dfxtp_1
X_2195_ clknet_leaf_223_clk booth_b14_m47 VGND VGND VPWR VPWR pp_row61_7 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_31_0 c$2870 c$2872 c$2874 VGND VGND VPWR VPWR c$3520 s$3521 sky130_fd_sc_hd__fa_1
Xdadda_fa_2_47_0 pp_row47_20 pp_row47_21 pp_row47_22 VGND VGND VPWR VPWR c$1290 s$1291
+ sky130_fd_sc_hd__fa_1
XU$$4250 net1256 notblock$6575\[1\] VGND VGND VPWR VPWR t$6576 sky130_fd_sc_hd__and2_1
XU$$4261 net939 net422 net1678 net704 VGND VGND VPWR VPWR t$6583 sky130_fd_sc_hd__a22o_1
XFILLER_93_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4272 t$6588 net1258 VGND VGND VPWR VPWR booth_b62_m9 sky130_fd_sc_hd__xor2_1
XU$$4283 net1178 net421 net1169 net703 VGND VGND VPWR VPWR t$6594 sky130_fd_sc_hd__a22o_1
X_1146_ clknet_leaf_15_clk booth_b0_m18 VGND VGND VPWR VPWR pp_row18_0 sky130_fd_sc_hd__dfxtp_1
XU$$4294 t$6599 net1255 VGND VGND VPWR VPWR booth_b62_m20 sky130_fd_sc_hd__xor2_1
XFILLER_37_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3560 t$6223 net1336 VGND VGND VPWR VPWR booth_b50_m64 sky130_fd_sc_hd__xor2_1
XU$$3571 t$6230 net1324 VGND VGND VPWR VPWR booth_b52_m1 sky130_fd_sc_hd__xor2_1
XU$$3582 net1522 net476 net1514 net749 VGND VGND VPWR VPWR t$6236 sky130_fd_sc_hd__a22o_1
XFILLER_129_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3593 t$6241 net1324 VGND VGND VPWR VPWR booth_b52_m12 sky130_fd_sc_hd__xor2_1
X_1077_ clknet_leaf_52_clk booth_b2_m9 VGND VGND VPWR VPWR pp_row11_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_179_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2870 net1550 net540 net1542 net813 VGND VGND VPWR VPWR t$5871 sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_8_1 pp_row8_5 pp_row8_6 s$2751 VGND VGND VPWR VPWR c$3430 s$3431 sky130_fd_sc_hd__fa_1
XU$$2881 notblock$5875\[2\] net37 net1379 t$5876 notblock$5875\[0\] VGND VGND VPWR
+ VPWR sel_0$5877 sky130_fd_sc_hd__a32o_4
XU$$2892 t$5883 net1368 VGND VGND VPWR VPWR booth_b42_m4 sky130_fd_sc_hd__xor2_1
XFILLER_178_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1979_ clknet_leaf_235_clk net206 VGND VGND VPWR VPWR pp_row54_29 sky130_fd_sc_hd__dfxtp_4
XFILLER_162_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_916 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_76_2 s$2449 s$2451 s$2453 VGND VGND VPWR VPWR c$3150 s$3151 sky130_fd_sc_hd__fa_1
XFILLER_88_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_69_1 c$2386 c$2388 s$2391 VGND VGND VPWR VPWR c$3106 s$3107 sky130_fd_sc_hd__fa_1
Xdadda_fa_7_46_0 s$3583 c$3986 s$3989 VGND VGND VPWR VPWR c$4244 s$4245 sky130_fd_sc_hd__fa_2
XFILLER_29_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$821 final_adder.p_new$836 final_adder.g_new$749 final_adder.g_new$837
+ VGND VGND VPWR VPWR final_adder.g_new$949 sky130_fd_sc_hd__a21o_2
XFILLER_75_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$843 final_adder.p_new$874 final_adder.g_new$939 final_adder.g_new$875
+ VGND VGND VPWR VPWR final_adder.g_new$971 sky130_fd_sc_hd__a21o_2
Xfinal_adder.U$$865 final_adder.p_new$896 final_adder.g_new$961 final_adder.g_new$897
+ VGND VGND VPWR VPWR final_adder.g_new$993 sky130_fd_sc_hd__a21o_1
XU$$704 t$4765 net1412 VGND VGND VPWR VPWR booth_b10_m6 sky130_fd_sc_hd__xor2_1
XU$$715 net1211 net406 net1204 net672 VGND VGND VPWR VPWR t$4771 sky130_fd_sc_hd__a22o_1
XFILLER_56_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$726 t$4776 net1412 VGND VGND VPWR VPWR booth_b10_m17 sky130_fd_sc_hd__xor2_1
XFILLER_16_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$887 final_adder.p_new$918 final_adder.g_new$751 final_adder.g_new$919
+ VGND VGND VPWR VPWR final_adder.g_new$1015 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$898 final_adder.$signal$1216 final_adder.g_new$965 final_adder.$signal$254
+ VGND VGND VPWR VPWR final_adder.g_new$1026 sky130_fd_sc_hd__a21o_1
XU$$737 net1100 net404 net1091 net670 VGND VGND VPWR VPWR t$4782 sky130_fd_sc_hd__a22o_1
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$748 t$4787 net1415 VGND VGND VPWR VPWR booth_b10_m28 sky130_fd_sc_hd__xor2_1
XU$$759 net990 net402 net982 net668 VGND VGND VPWR VPWR t$4793 sky130_fd_sc_hd__a22o_1
XFILLER_25_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_9 final_adder.g_new$967 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_71_1 c$1570 c$1572 c$1574 VGND VGND VPWR VPWR c$2408 s$2409 sky130_fd_sc_hd__fa_1
XFILLER_106_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1010 net1011 VGND VGND VPWR VPWR net1010 sky130_fd_sc_hd__buf_6
Xdadda_fa_3_64_0 s$617 c$1482 c$1484 VGND VGND VPWR VPWR c$2350 s$2351 sky130_fd_sc_hd__fa_1
XFILLER_117_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1021 net1022 VGND VGND VPWR VPWR net1021 sky130_fd_sc_hd__buf_6
XFILLER_6_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1032 net1033 VGND VGND VPWR VPWR net1032 sky130_fd_sc_hd__buf_4
Xfanout1043 net1045 VGND VGND VPWR VPWR net1043 sky130_fd_sc_hd__buf_4
XFILLER_121_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1054 net85 VGND VGND VPWR VPWR net1054 sky130_fd_sc_hd__buf_6
Xfanout1065 net83 VGND VGND VPWR VPWR net1065 sky130_fd_sc_hd__buf_2
Xfanout1076 net1078 VGND VGND VPWR VPWR net1076 sky130_fd_sc_hd__buf_4
Xfanout1087 net81 VGND VGND VPWR VPWR net1087 sky130_fd_sc_hd__buf_4
XFILLER_47_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1098 net1099 VGND VGND VPWR VPWR net1098 sky130_fd_sc_hd__clkbuf_8
X_1000_ clknet_leaf_119_clk booth_b40_m61 VGND VGND VPWR VPWR pp_row101_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_74_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2100 t$5478 net1440 VGND VGND VPWR VPWR booth_b30_m19 sky130_fd_sc_hd__xor2_1
XU$$2111 net1084 net580 net1074 net853 VGND VGND VPWR VPWR t$5484 sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_100_1 c$2634 c$2636 s$2639 VGND VGND VPWR VPWR c$3292 s$3293 sky130_fd_sc_hd__fa_1
XU$$2122 t$5489 net1440 VGND VGND VPWR VPWR booth_b30_m30 sky130_fd_sc_hd__xor2_1
XU$$2133 net978 net580 net972 net853 VGND VGND VPWR VPWR t$5495 sky130_fd_sc_hd__a22o_1
XU$$2144 t$5500 net1445 VGND VGND VPWR VPWR booth_b30_m41 sky130_fd_sc_hd__xor2_1
XU$$1410 net1157 net629 net1147 net902 VGND VGND VPWR VPWR t$5126 sky130_fd_sc_hd__a22o_1
XU$$2155 net1705 net579 net1697 net852 VGND VGND VPWR VPWR t$5506 sky130_fd_sc_hd__a22o_1
XU$$2166 t$5511 net1445 VGND VGND VPWR VPWR booth_b30_m52 sky130_fd_sc_hd__xor2_1
XU$$1421 t$5131 net1486 VGND VGND VPWR VPWR booth_b20_m22 sky130_fd_sc_hd__xor2_1
XFILLER_62_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1432 net1056 net628 net1048 net901 VGND VGND VPWR VPWR t$5137 sky130_fd_sc_hd__a22o_1
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2177 net1598 net582 net1589 net855 VGND VGND VPWR VPWR t$5517 sky130_fd_sc_hd__a22o_1
XU$$2188 t$5522 net1447 VGND VGND VPWR VPWR booth_b30_m63 sky130_fd_sc_hd__xor2_1
XU$$1443 t$5142 net1488 VGND VGND VPWR VPWR booth_b20_m33 sky130_fd_sc_hd__xor2_1
XU$$1454 net949 net632 net941 net905 VGND VGND VPWR VPWR t$5148 sky130_fd_sc_hd__a22o_1
XFILLER_62_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2199 t$5529 net1432 VGND VGND VPWR VPWR booth_b32_m0 sky130_fd_sc_hd__xor2_1
XU$$1465 t$5153 net1493 VGND VGND VPWR VPWR booth_b20_m44 sky130_fd_sc_hd__xor2_1
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1476 net1683 net634 net1657 net907 VGND VGND VPWR VPWR t$5159 sky130_fd_sc_hd__a22o_1
X_1902_ clknet_leaf_71_clk booth_b34_m18 VGND VGND VPWR VPWR pp_row52_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_163_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1487 t$5164 net1492 VGND VGND VPWR VPWR booth_b20_m55 sky130_fd_sc_hd__xor2_1
Xdadda_fa_7_121_0 s$3883 c$4136 s$4139 VGND VGND VPWR VPWR c$4394 s$4395 sky130_fd_sc_hd__fa_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1498 net1553 net633 net1544 net906 VGND VGND VPWR VPWR t$5170 sky130_fd_sc_hd__a22o_1
XFILLER_124_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1833_ clknet_leaf_18_clk booth_b20_m30 VGND VGND VPWR VPWR pp_row50_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_191_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1764_ clknet_leaf_235_clk booth_b0_m48 VGND VGND VPWR VPWR pp_row48_0 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_86_1 s$3207 s$3209 s$3211 VGND VGND VPWR VPWR c$3742 s$3743 sky130_fd_sc_hd__fa_1
X_0715_ clknet_leaf_165_clk booth_b60_m27 VGND VGND VPWR VPWR pp_row87_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_144_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1695_ clknet_leaf_18_clk booth_b26_m19 VGND VGND VPWR VPWR pp_row45_13 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_79_0 c$3158 c$3160 c$3162 VGND VGND VPWR VPWR c$3712 s$3713 sky130_fd_sc_hd__fa_1
XFILLER_144_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0646_ clknet_leaf_182_clk booth_b26_m59 VGND VGND VPWR VPWR pp_row85_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_135_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_12__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_5_12__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_135_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_78_8 pp_row78_26 pp_row78_27 c$200 VGND VGND VPWR VPWR c$868 s$869 sky130_fd_sc_hd__fa_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0577_ clknet_leaf_120_clk booth_b60_m56 VGND VGND VPWR VPWR pp_row116_5 sky130_fd_sc_hd__dfxtp_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2316_ clknet_leaf_184_clk net141 VGND VGND VPWR VPWR pp_row110_11 sky130_fd_sc_hd__dfxtp_2
XFILLER_85_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$106 c$4362 s$4365 VGND VGND VPWR VPWR final_adder.$signal$214 final_adder.$signal$1196
+ sky130_fd_sc_hd__ha_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$117 c$4384 s$4387 VGND VGND VPWR VPWR final_adder.$signal$236 final_adder.$signal$1207
+ sky130_fd_sc_hd__ha_1
XFILLER_39_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$139 final_adder.$signal$1207 final_adder.$signal$234 final_adder.$signal$236
+ VGND VGND VPWR VPWR final_adder.g_new$267 sky130_fd_sc_hd__a21o_1
XFILLER_85_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2247_ clknet_leaf_213_clk booth_b46_m16 VGND VGND VPWR VPWR pp_row62_23 sky130_fd_sc_hd__dfxtp_1
XFILLER_100_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2178_ clknet_leaf_224_clk booth_b50_m10 VGND VGND VPWR VPWR pp_row60_25 sky130_fd_sc_hd__dfxtp_1
XFILLER_122_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4080 t$6489 net1285 VGND VGND VPWR VPWR booth_b58_m50 sky130_fd_sc_hd__xor2_1
XU$$3422_1792 VGND VGND VPWR VPWR U$$3422_1792/HI net1792 sky130_fd_sc_hd__conb_1
XU$$4091 net1617 net456 net1610 net729 VGND VGND VPWR VPWR t$6495 sky130_fd_sc_hd__a22o_1
X_1129_ clknet_leaf_13_clk booth_b10_m6 VGND VGND VPWR VPWR pp_row16_5 sky130_fd_sc_hd__dfxtp_1
XU$$3390 net1700 net498 net1693 net771 VGND VGND VPWR VPWR t$6137 sky130_fd_sc_hd__a22o_1
XFILLER_40_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_81_0 s$1709 c$2478 c$2480 VGND VGND VPWR VPWR c$3176 s$3177 sky130_fd_sc_hd__fa_1
XFILLER_190_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_102_3 s$1943 s$1945 s$1947 VGND VGND VPWR VPWR c$2660 s$2661 sky130_fd_sc_hd__fa_1
XFILLER_134_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_746 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput102 b[43] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_4
XFILLER_103_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput113 b[53] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__buf_2
XFILLER_89_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput124 b[63] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__buf_4
XFILLER_103_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput135 c[105] VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_1
Xinput146 c[115] VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_1
Xinput157 c[125] VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_1
Xinput168 c[1] VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$640 final_adder.p_new$664 final_adder.p_new$648 VGND VGND VPWR VPWR
+ final_adder.p_new$768 sky130_fd_sc_hd__and2_1
Xinput179 c[2] VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_1
XTAP_3922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$651 final_adder.p_new$658 final_adder.g_new$675 final_adder.g_new$659
+ VGND VGND VPWR VPWR final_adder.g_new$779 sky130_fd_sc_hd__a21o_1
XTAP_3933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$501 net1745 net426 net1737 net708 VGND VGND VPWR VPWR t$4661 sky130_fd_sc_hd__a22o_1
XFILLER_99_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_109_0 c$3828 c$3830 s$3833 VGND VGND VPWR VPWR c$4114 s$4115 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$662 final_adder.p_new$686 final_adder.p_new$670 VGND VGND VPWR VPWR
+ final_adder.p_new$790 sky130_fd_sc_hd__and2_1
XTAP_3944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$673 final_adder.p_new$680 final_adder.g_new$697 final_adder.g_new$681
+ VGND VGND VPWR VPWR final_adder.g_new$801 sky130_fd_sc_hd__a21o_1
XU$$512 t$4666 net1250 VGND VGND VPWR VPWR booth_b6_m47 sky130_fd_sc_hd__xor2_1
XTAP_3955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$523 net1638 net428 net1629 net710 VGND VGND VPWR VPWR t$4672 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$684 final_adder.p_new$708 final_adder.p_new$692 VGND VGND VPWR VPWR
+ final_adder.p_new$812 sky130_fd_sc_hd__and2_1
XTAP_3966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$534 t$4677 net1246 VGND VGND VPWR VPWR booth_b6_m58 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$695 final_adder.p_new$702 final_adder.g_new$719 final_adder.g_new$703
+ VGND VGND VPWR VPWR final_adder.g_new$823 sky130_fd_sc_hd__a21o_1
XFILLER_186_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$545 net1531 net432 net1881 net714 VGND VGND VPWR VPWR t$4683 sky130_fd_sc_hd__a22o_1
XTAP_3988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$556 net1231 net413 net1127 net679 VGND VGND VPWR VPWR t$4690 sky130_fd_sc_hd__a22o_1
XTAP_3999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_29_3 s$1083 s$1085 s$1087 VGND VGND VPWR VPWR c$2076 s$2077 sky130_fd_sc_hd__fa_1
XFILLER_72_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$567 t$4695 net1241 VGND VGND VPWR VPWR booth_b8_m6 sky130_fd_sc_hd__xor2_1
XU$$578 net1216 net413 net1206 net679 VGND VGND VPWR VPWR t$4701 sky130_fd_sc_hd__a22o_1
XFILLER_147_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$589 t$4706 net1236 VGND VGND VPWR VPWR booth_b8_m17 sky130_fd_sc_hd__xor2_1
XFILLER_189_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_6_96_0 c$3776 c$3778 s$3781 VGND VGND VPWR VPWR c$4088 s$4089 sky130_fd_sc_hd__fa_1
XFILLER_184_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0500_ clknet_leaf_179_clk booth_b62_m64 VGND VGND VPWR VPWR pp_row126_1 sky130_fd_sc_hd__dfxtp_1
X_1480_ clknet_leaf_241_clk booth_b0_m37 VGND VGND VPWR VPWR pp_row37_0 sky130_fd_sc_hd__dfxtp_1
X_0431_ clknet_leaf_154_clk booth_b48_m29 VGND VGND VPWR VPWR pp_row77_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0362_ clknet_leaf_192_clk booth_b36_m39 VGND VGND VPWR VPWR pp_row75_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_94_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_2_32_5 pp_row32_15 pp_row32_16 VGND VGND VPWR VPWR c$1120 s$1121 sky130_fd_sc_hd__ha_2
X_2101_ clknet_leaf_32_clk booth_b38_m20 VGND VGND VPWR VPWR pp_row58_19 sky130_fd_sc_hd__dfxtp_1
X_0293_ clknet_leaf_199_clk booth_b26_m47 VGND VGND VPWR VPWR pp_row73_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_55_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2032_ clknet_leaf_72_clk booth_b36_m20 VGND VGND VPWR VPWR pp_row56_18 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_31_3 pp_row31_9 pp_row31_10 pp_row31_11 VGND VGND VPWR VPWR c$1106 s$1107
+ sky130_fd_sc_hd__fa_1
XFILLER_47_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1240 t$5039 net1664 VGND VGND VPWR VPWR booth_b18_m0 sky130_fd_sc_hd__xor2_1
XU$$1251 net1561 net635 net1521 net908 VGND VGND VPWR VPWR t$5045 sky130_fd_sc_hd__a22o_1
XU$$1262 t$5050 net1662 VGND VGND VPWR VPWR booth_b18_m11 sky130_fd_sc_hd__xor2_1
XU$$1273 net1161 net637 net1149 net910 VGND VGND VPWR VPWR t$5056 sky130_fd_sc_hd__a22o_1
XFILLER_50_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1284 t$5061 net1667 VGND VGND VPWR VPWR booth_b18_m22 sky130_fd_sc_hd__xor2_1
XU$$1295 net1056 net639 net1048 net912 VGND VGND VPWR VPWR t$5067 sky130_fd_sc_hd__a22o_1
X_1816_ clknet_leaf_141_clk booth_b46_m61 VGND VGND VPWR VPWR pp_row107_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_163_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1747_ clknet_leaf_238_clk booth_b20_m27 VGND VGND VPWR VPWR pp_row47_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_117_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1678_ clknet_leaf_239_clk net1357 VGND VGND VPWR VPWR pp_row44_23 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_83_6 pp_row83_18 pp_row83_19 pp_row83_20 VGND VGND VPWR VPWR c$950 s$951
+ sky130_fd_sc_hd__fa_1
Xfanout803 sel_1$4548 VGND VGND VPWR VPWR net803 sky130_fd_sc_hd__buf_6
XFILLER_132_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout814 net815 VGND VGND VPWR VPWR net814 sky130_fd_sc_hd__clkbuf_4
X_0629_ clknet_leaf_177_clk booth_b44_m40 VGND VGND VPWR VPWR pp_row84_13 sky130_fd_sc_hd__dfxtp_1
Xfanout825 net826 VGND VGND VPWR VPWR net825 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_1_76_5 pp_row76_20 pp_row76_21 pp_row76_22 VGND VGND VPWR VPWR c$826 s$827
+ sky130_fd_sc_hd__fa_1
Xfanout836 net837 VGND VGND VPWR VPWR net836 sky130_fd_sc_hd__buf_4
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout847 net848 VGND VGND VPWR VPWR net847 sky130_fd_sc_hd__buf_4
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout858 net859 VGND VGND VPWR VPWR net858 sky130_fd_sc_hd__clkbuf_4
XFILLER_140_780 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_69_4 pp_row69_27 pp_row69_28 pp_row69_29 VGND VGND VPWR VPWR c$698 s$699
+ sky130_fd_sc_hd__fa_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout869 net870 VGND VGND VPWR VPWR net869 sky130_fd_sc_hd__buf_4
XFILLER_133_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_39_2 s$2153 s$2155 s$2157 VGND VGND VPWR VPWR c$2928 s$2929 sky130_fd_sc_hd__fa_1
XFILLER_85_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_207 net1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_218 net1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_229 net1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_817 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_100_0 pp_row100_14 pp_row100_15 pp_row100_16 VGND VGND VPWR VPWR c$2638
+ s$2639 sky130_fd_sc_hd__fa_1
XFILLER_135_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_0_64_3 pp_row64_9 pp_row64_10 pp_row64_11 VGND VGND VPWR VPWR c$90 s$91
+ sky130_fd_sc_hd__fa_1
XFILLER_190_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_41_2 c$1216 s$1219 s$1221 VGND VGND VPWR VPWR c$2170 s$2171 sky130_fd_sc_hd__fa_1
XFILLER_188_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$470 final_adder.p_new$476 final_adder.p_new$472 VGND VGND VPWR VPWR
+ final_adder.p_new$598 sky130_fd_sc_hd__and2_1
XTAP_3752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$320 net1131 net528 net1115 net801 VGND VGND VPWR VPWR t$4569 sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_34_1 c$1126 c$1128 c$1130 VGND VGND VPWR VPWR c$2112 s$2113 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$481 final_adder.p_new$482 final_adder.g_new$487 final_adder.g_new$483
+ VGND VGND VPWR VPWR final_adder.g_new$609 sky130_fd_sc_hd__a21o_1
XTAP_3763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$492 final_adder.p_new$498 final_adder.p_new$494 VGND VGND VPWR VPWR
+ final_adder.p_new$620 sky130_fd_sc_hd__and2_1
XU$$331 t$4574 net1273 VGND VGND VPWR VPWR booth_b4_m25 sky130_fd_sc_hd__xor2_1
XTAP_3774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$342 net1026 net534 net1018 net807 VGND VGND VPWR VPWR t$4580 sky130_fd_sc_hd__a22o_1
XTAP_3785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$353 t$4585 net1273 VGND VGND VPWR VPWR booth_b4_m36 sky130_fd_sc_hd__xor2_1
XFILLER_91_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_11_0 c$3436 c$3438 s$3441 VGND VGND VPWR VPWR c$3918 s$3919 sky130_fd_sc_hd__fa_1
Xdadda_fa_3_27_0 pp_row27_8 pp_row27_9 pp_row27_10 VGND VGND VPWR VPWR c$2054 s$2055
+ sky130_fd_sc_hd__fa_1
XFILLER_60_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$364 net1745 net529 net1737 net802 VGND VGND VPWR VPWR t$4591 sky130_fd_sc_hd__a22o_1
XU$$375 t$4596 net1278 VGND VGND VPWR VPWR booth_b4_m47 sky130_fd_sc_hd__xor2_1
XFILLER_45_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$386 net1641 net533 net1633 net806 VGND VGND VPWR VPWR t$4602 sky130_fd_sc_hd__a22o_1
XU$$397 t$4607 net1275 VGND VGND VPWR VPWR booth_b4_m58 sky130_fd_sc_hd__xor2_1
XFILLER_189_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0980_ clknet_leaf_114_clk booth_b36_m64 VGND VGND VPWR VPWR pp_row100_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_13_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1601_ clknet_leaf_243_clk booth_b2_m40 VGND VGND VPWR VPWR pp_row42_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_8_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_93_5 c$1034 c$1036 s$1039 VGND VGND VPWR VPWR c$1852 s$1853 sky130_fd_sc_hd__fa_1
Xclkbuf_leaf_247_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_247_clk
+ sky130_fd_sc_hd__clkbuf_16
X_1532_ clknet_leaf_44_clk booth_b8_m31 VGND VGND VPWR VPWR pp_row39_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_99_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_86_4 c$976 s$979 s$981 VGND VGND VPWR VPWR c$1766 s$1767 sky130_fd_sc_hd__fa_1
XFILLER_10_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_79_3 c$868 s$871 s$873 VGND VGND VPWR VPWR c$1680 s$1681 sky130_fd_sc_hd__fa_2
X_1463_ clknet_leaf_40_clk booth_b10_m26 VGND VGND VPWR VPWR pp_row36_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_45_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0414_ clknet_leaf_193_clk booth_b16_m61 VGND VGND VPWR VPWR pp_row77_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_79_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1394_ clknet_leaf_164_clk notsign$6504 VGND VGND VPWR VPWR pp_row123_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_68_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_49_1 s$2985 s$2987 s$2989 VGND VGND VPWR VPWR c$3594 s$3595 sky130_fd_sc_hd__fa_1
X_0345_ clknet_leaf_203_clk booth_b62_m12 VGND VGND VPWR VPWR pp_row74_27 sky130_fd_sc_hd__dfxtp_1
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0276_ clknet_leaf_202_clk booth_b58_m14 VGND VGND VPWR VPWR pp_row72_26 sky130_fd_sc_hd__dfxtp_1
XFILLER_82_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2015_ clknet_leaf_81_clk booth_b6_m50 VGND VGND VPWR VPWR pp_row56_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_51_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_102_2 pp_row102_6 pp_row102_7 pp_row102_8 VGND VGND VPWR VPWR c$1946 s$1947
+ sky130_fd_sc_hd__fa_1
XFILLER_169_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1070 t$4951 net1191 VGND VGND VPWR VPWR booth_b14_m52 sky130_fd_sc_hd__xor2_1
XFILLER_177_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1081 net1596 net390 net1587 net656 VGND VGND VPWR VPWR t$4957 sky130_fd_sc_hd__a22o_1
XU$$1092 t$4962 net1188 VGND VGND VPWR VPWR booth_b14_m63 sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_123_1 pp_row123_3 pp_row123_4 c$3414 VGND VGND VPWR VPWR c$3890 s$3891
+ sky130_fd_sc_hd__fa_1
XFILLER_12_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_116_0 c$3380 c$3382 c$3384 VGND VGND VPWR VPWR c$3860 s$3861 sky130_fd_sc_hd__fa_1
XFILLER_163_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_238_clk clknet_5_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_238_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_2_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_81_3 pp_row81_9 pp_row81_10 pp_row81_11 VGND VGND VPWR VPWR c$912 s$913
+ sky130_fd_sc_hd__fa_1
XFILLER_132_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout600 net601 VGND VGND VPWR VPWR net600 sky130_fd_sc_hd__buf_6
Xfanout1609 net1610 VGND VGND VPWR VPWR net1609 sky130_fd_sc_hd__buf_4
Xfanout611 net612 VGND VGND VPWR VPWR net611 sky130_fd_sc_hd__buf_2
Xfanout622 sel_0$4477 VGND VGND VPWR VPWR net622 sky130_fd_sc_hd__clkbuf_8
Xdadda_fa_1_74_2 pp_row74_14 pp_row74_15 pp_row74_16 VGND VGND VPWR VPWR c$784 s$785
+ sky130_fd_sc_hd__fa_1
Xfanout633 net634 VGND VGND VPWR VPWR net633 sky130_fd_sc_hd__clkbuf_4
Xfanout644 net647 VGND VGND VPWR VPWR net644 sky130_fd_sc_hd__buf_6
Xdadda_fa_4_51_1 c$2242 c$2244 s$2247 VGND VGND VPWR VPWR c$2998 s$2999 sky130_fd_sc_hd__fa_1
Xfanout655 net658 VGND VGND VPWR VPWR net655 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_1_67_1 pp_row67_21 pp_row67_22 pp_row67_23 VGND VGND VPWR VPWR c$656 s$657
+ sky130_fd_sc_hd__fa_1
Xfanout666 sel_1$4828 VGND VGND VPWR VPWR net666 sky130_fd_sc_hd__buf_6
Xfanout677 net678 VGND VGND VPWR VPWR net677 sky130_fd_sc_hd__buf_4
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout688 net689 VGND VGND VPWR VPWR net688 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_4_44_0 s$1265 c$2182 c$2184 VGND VGND VPWR VPWR c$2954 s$2955 sky130_fd_sc_hd__fa_1
Xfanout699 sel_1$6648 VGND VGND VPWR VPWR net699 sky130_fd_sc_hd__clkbuf_8
XTAP_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_96_3 s$1883 s$1885 s$1887 VGND VGND VPWR VPWR c$2612 s$2613 sky130_fd_sc_hd__fa_1
XFILLER_6_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_229_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_229_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_89_2 c$1792 s$1795 s$1797 VGND VGND VPWR VPWR c$2554 s$2555 sky130_fd_sc_hd__fa_1
Xdadda_fa_2_100_0_1904 VGND VGND VPWR VPWR net1904 dadda_fa_2_100_0_1904/LO sky130_fd_sc_hd__conb_1
XFILLER_135_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_59_0 c$3628 c$3630 s$3633 VGND VGND VPWR VPWR c$4014 s$4015 sky130_fd_sc_hd__fa_1
XFILLER_151_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_0_62_0 pp_row62_0 pp_row62_1 pp_row62_2 VGND VGND VPWR VPWR c$60 s$61 sky130_fd_sc_hd__fa_1
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_815 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3901 t$6398 net1294 VGND VGND VPWR VPWR booth_b56_m29 sky130_fd_sc_hd__xor2_1
XFILLER_77_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3912 net988 net464 net979 net737 VGND VGND VPWR VPWR t$6404 sky130_fd_sc_hd__a22o_1
XFILLER_65_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3923 t$6409 net1299 VGND VGND VPWR VPWR booth_b56_m40 sky130_fd_sc_hd__xor2_1
XTAP_4272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3934 net1718 net466 net1709 net739 VGND VGND VPWR VPWR t$6415 sky130_fd_sc_hd__a22o_1
XFILLER_92_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3945 t$6420 net1293 VGND VGND VPWR VPWR booth_b56_m51 sky130_fd_sc_hd__xor2_1
XFILLER_18_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3956 net1608 net465 net1600 net738 VGND VGND VPWR VPWR t$6426 sky130_fd_sc_hd__a22o_1
XTAP_3560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3967 t$6431 net1293 VGND VGND VPWR VPWR booth_b56_m62 sky130_fd_sc_hd__xor2_1
XTAP_3571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3978 net54 net1292 VGND VGND VPWR VPWR sel_1$6438 sky130_fd_sc_hd__xor2_1
XU$$150 t$4482 net1390 VGND VGND VPWR VPWR booth_b2_m3 sky130_fd_sc_hd__xor2_1
XTAP_3582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3989 net1674 net451 net1563 net724 VGND VGND VPWR VPWR t$6444 sky130_fd_sc_hd__a22o_1
XTAP_3593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$161 net1508 net624 net1499 net897 VGND VGND VPWR VPWR t$4488 sky130_fd_sc_hd__a22o_1
XFILLER_17_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$172 t$4493 net1386 VGND VGND VPWR VPWR booth_b2_m14 sky130_fd_sc_hd__xor2_1
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$183 net1133 net623 net1117 net896 VGND VGND VPWR VPWR t$4499 sky130_fd_sc_hd__a22o_1
XU$$194 t$4504 net1385 VGND VGND VPWR VPWR booth_b2_m25 sky130_fd_sc_hd__xor2_1
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0963_ clknet_leaf_114_clk booth_b38_m61 VGND VGND VPWR VPWR pp_row99_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_186_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0894_ clknet_leaf_100_clk booth_b54_m41 VGND VGND VPWR VPWR pp_row95_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_185_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_91_2 pp_row91_15 pp_row91_16 pp_row91_17 VGND VGND VPWR VPWR c$1822 s$1823
+ sky130_fd_sc_hd__fa_2
Xdadda_fa_2_84_1 pp_row84_23 pp_row84_24 c$938 VGND VGND VPWR VPWR c$1736 s$1737 sky130_fd_sc_hd__fa_1
XFILLER_114_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput258 net258 VGND VGND VPWR VPWR o[100] sky130_fd_sc_hd__buf_2
X_1515_ clknet_leaf_17_clk booth_b22_m16 VGND VGND VPWR VPWR pp_row38_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_142_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput269 net269 VGND VGND VPWR VPWR o[110] sky130_fd_sc_hd__buf_2
Xdadda_fa_5_61_0 c$3050 c$3052 c$3054 VGND VGND VPWR VPWR c$3640 s$3641 sky130_fd_sc_hd__fa_1
X_2495_ clknet_leaf_142_clk booth_b30_m39 VGND VGND VPWR VPWR pp_row69_13 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_77_0 s$201 c$816 c$818 VGND VGND VPWR VPWR c$1650 s$1651 sky130_fd_sc_hd__fa_1
XFILLER_141_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1446_ clknet_leaf_64_clk booth_b18_m17 VGND VGND VPWR VPWR pp_row35_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_60_8 s$43 s$45 s$47 VGND VGND VPWR VPWR c$544 s$545 sky130_fd_sc_hd__fa_1
X_1377_ clknet_leaf_7_clk booth_b10_m22 VGND VGND VPWR VPWR pp_row32_5 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_53_7 pp_row53_23 pp_row53_24 pp_row53_25 VGND VGND VPWR VPWR c$416 s$417
+ sky130_fd_sc_hd__fa_1
XFILLER_56_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0328_ clknet_leaf_227_clk booth_b32_m42 VGND VGND VPWR VPWR pp_row74_12 sky130_fd_sc_hd__dfxtp_1
X_0259_ clknet_leaf_211_clk booth_b26_m46 VGND VGND VPWR VPWR pp_row72_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_1135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_99_1 c$2626 c$2628 s$2631 VGND VGND VPWR VPWR c$3286 s$3287 sky130_fd_sc_hd__fa_1
XFILLER_164_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_76_0 s$3703 c$4046 s$4049 VGND VGND VPWR VPWR c$4304 s$4305 sky130_fd_sc_hd__fa_2
XFILLER_136_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1406 net1407 VGND VGND VPWR VPWR net1406 sky130_fd_sc_hd__buf_6
XFILLER_48_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1417 net1418 VGND VGND VPWR VPWR net1417 sky130_fd_sc_hd__buf_4
XFILLER_28_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1428 net1429 VGND VGND VPWR VPWR net1428 sky130_fd_sc_hd__buf_6
Xfanout430 net431 VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__buf_4
XFILLER_132_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1439 net1440 VGND VGND VPWR VPWR net1439 sky130_fd_sc_hd__buf_6
Xfanout441 sel_0$6507 VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__clkbuf_4
Xfanout452 net459 VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__buf_2
Xfanout463 sel_0$6367 VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__clkbuf_8
XFILLER_48_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout474 net475 VGND VGND VPWR VPWR net474 sky130_fd_sc_hd__buf_4
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout485 net487 VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__buf_4
Xfanout496 sel_0$6087 VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__buf_4
XFILLER_111_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3208 t$6044 net1349 VGND VGND VPWR VPWR booth_b46_m25 sky130_fd_sc_hd__xor2_1
XFILLER_0_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3219 net1027 net502 net1019 net775 VGND VGND VPWR VPWR t$6050 sky130_fd_sc_hd__a22o_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2507 t$5686 net1406 VGND VGND VPWR VPWR booth_b36_m17 sky130_fd_sc_hd__xor2_1
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2518 net1098 net552 net1090 net825 VGND VGND VPWR VPWR t$5692 sky130_fd_sc_hd__a22o_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2529 t$5697 net1406 VGND VGND VPWR VPWR booth_b36_m28 sky130_fd_sc_hd__xor2_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1806 t$5328 net1460 VGND VGND VPWR VPWR booth_b26_m9 sky130_fd_sc_hd__xor2_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1817 net1173 net593 net1164 net866 VGND VGND VPWR VPWR t$5334 sky130_fd_sc_hd__a22o_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1828 t$5339 net1458 VGND VGND VPWR VPWR booth_b26_m20 sky130_fd_sc_hd__xor2_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1839 net1074 net596 net1066 net869 VGND VGND VPWR VPWR t$5345 sky130_fd_sc_hd__a22o_1
XFILLER_15_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_94_0 s$1045 c$1842 c$1844 VGND VGND VPWR VPWR c$2590 s$2591 sky130_fd_sc_hd__fa_1
XFILLER_143_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1300_ clknet_leaf_250_clk booth_b6_m22 VGND VGND VPWR VPWR pp_row28_3 sky130_fd_sc_hd__dfxtp_1
X_2280_ clknet_leaf_212_clk booth_b38_m25 VGND VGND VPWR VPWR pp_row63_19 sky130_fd_sc_hd__dfxtp_1
X_1231_ clknet_leaf_12_clk booth_b2_m22 VGND VGND VPWR VPWR pp_row24_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_96_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4410 net1502 sel_0$6647 net1222 net694 VGND VGND VPWR VPWR t$6659 sky130_fd_sc_hd__a22o_1
XU$$4421 t$6664 net1831 VGND VGND VPWR VPWR booth_b64_m15 sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_56_5 s$467 s$469 s$471 VGND VGND VPWR VPWR c$1408 s$1409 sky130_fd_sc_hd__fa_2
XU$$4432 net1119 sel_0$6647 net1112 net693 VGND VGND VPWR VPWR t$6670 sky130_fd_sc_hd__a22o_1
XU$$4443 t$6675 net1842 VGND VGND VPWR VPWR booth_b64_m26 sky130_fd_sc_hd__xor2_1
XFILLER_49_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1162_ clknet_leaf_46_clk booth_b4_m15 VGND VGND VPWR VPWR pp_row19_2 sky130_fd_sc_hd__dfxtp_1
XU$$4454 net1022 sel_0$6647 net1005 net699 VGND VGND VPWR VPWR t$6681 sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_49_4 s$335 s$337 s$339 VGND VGND VPWR VPWR c$1322 s$1323 sky130_fd_sc_hd__fa_1
XU$$4465 t$6686 net1853 VGND VGND VPWR VPWR booth_b64_m37 sky130_fd_sc_hd__xor2_1
XU$$3720 t$6306 net1300 VGND VGND VPWR VPWR booth_b54_m7 sky130_fd_sc_hd__xor2_1
XU$$3731 net1208 net472 net1200 net745 VGND VGND VPWR VPWR t$6312 sky130_fd_sc_hd__a22o_1
XFILLER_53_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4476 net1743 sel_0$6647 net1735 net696 VGND VGND VPWR VPWR t$6692 sky130_fd_sc_hd__a22o_1
XTAP_4080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4487 t$6697 net1864 VGND VGND VPWR VPWR booth_b64_m48 sky130_fd_sc_hd__xor2_1
XU$$3742 t$6317 net1300 VGND VGND VPWR VPWR booth_b54_m18 sky130_fd_sc_hd__xor2_1
XTAP_4091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1093_ clknet_leaf_59_clk booth_b0_m13 VGND VGND VPWR VPWR pp_row13_0 sky130_fd_sc_hd__dfxtp_1
XU$$3753 net1094 net468 net1086 net741 VGND VGND VPWR VPWR t$6323 sky130_fd_sc_hd__a22o_1
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4498 net1636 sel_0$6647 net1625 net696 VGND VGND VPWR VPWR t$6703 sky130_fd_sc_hd__a22o_1
XU$$3764 t$6328 net1303 VGND VGND VPWR VPWR booth_b54_m29 sky130_fd_sc_hd__xor2_1
XFILLER_46_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3775 net985 net470 net976 net743 VGND VGND VPWR VPWR t$6334 sky130_fd_sc_hd__a22o_1
XFILLER_64_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3786 t$6339 net1305 VGND VGND VPWR VPWR booth_b54_m40 sky130_fd_sc_hd__xor2_1
XU$$3797 net1718 net474 net1709 net747 VGND VGND VPWR VPWR t$6345 sky130_fd_sc_hd__a22o_1
XTAP_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4507_1874 VGND VGND VPWR VPWR U$$4507_1874/HI net1874 sky130_fd_sc_hd__conb_1
XANTENNA_390 net1518 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1995_ clknet_leaf_67_clk booth_b26_m29 VGND VGND VPWR VPWR pp_row55_13 sky130_fd_sc_hd__dfxtp_1
X_0946_ clknet_leaf_113_clk booth_b40_m58 VGND VGND VPWR VPWR pp_row98_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_118_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_978 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0877_ clknet_leaf_133_clk booth_b58_m62 VGND VGND VPWR VPWR pp_row120_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_109_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_1_45_5 pp_row45_15 pp_row45_16 VGND VGND VPWR VPWR c$286 s$287 sky130_fd_sc_hd__ha_1
XFILLER_87_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2478_ clknet_leaf_99_clk booth_b64_m4 VGND VGND VPWR VPWR pp_row68_31 sky130_fd_sc_hd__dfxtp_1
XFILLER_130_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1429_ clknet_leaf_64_clk booth_b26_m8 VGND VGND VPWR VPWR pp_row34_13 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_51_4 pp_row51_12 pp_row51_13 pp_row51_14 VGND VGND VPWR VPWR c$374 s$375
+ sky130_fd_sc_hd__fa_1
XFILLER_28_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$908 net944 net397 net928 net663 VGND VGND VPWR VPWR t$4869 sky130_fd_sc_hd__a22o_1
XU$$919 t$4874 net1315 VGND VGND VPWR VPWR booth_b12_m45 sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_44_3 pp_row44_9 pp_row44_10 pp_row44_11 VGND VGND VPWR VPWR c$270 s$271
+ sky130_fd_sc_hd__fa_1
Xdadda_fa_4_21_2 s$2009 s$2011 s$2013 VGND VGND VPWR VPWR c$2820 s$2821 sky130_fd_sc_hd__fa_1
XFILLER_37_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_14_1 pp_row14_5 pp_row14_6 pp_row14_7 VGND VGND VPWR VPWR c$2776 s$2777
+ sky130_fd_sc_hd__fa_1
XFILLER_110_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1203 net1204 VGND VGND VPWR VPWR net1203 sky130_fd_sc_hd__buf_4
XFILLER_160_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1214 net1215 VGND VGND VPWR VPWR net1214 sky130_fd_sc_hd__buf_6
Xfanout1225 net1226 VGND VGND VPWR VPWR net1225 sky130_fd_sc_hd__buf_2
XFILLER_182_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1236 net64 VGND VGND VPWR VPWR net1236 sky130_fd_sc_hd__clkbuf_8
Xfanout1247 net1253 VGND VGND VPWR VPWR net1247 sky130_fd_sc_hd__buf_4
Xfanout1258 net60 VGND VGND VPWR VPWR net1258 sky130_fd_sc_hd__buf_4
Xdadda_fa_3_59_3 s$1439 s$1441 s$1443 VGND VGND VPWR VPWR c$2316 s$2317 sky130_fd_sc_hd__fa_1
Xfanout1269 net1272 VGND VGND VPWR VPWR net1269 sky130_fd_sc_hd__buf_6
XFILLER_8_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3005 net1556 net525 net1548 net798 VGND VGND VPWR VPWR t$5940 sky130_fd_sc_hd__a22o_1
XU$$3016 net1359 VGND VGND VPWR VPWR notblock$5945\[2\] sky130_fd_sc_hd__inv_1
XFILLER_86_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3027 t$5952 net1357 VGND VGND VPWR VPWR booth_b44_m3 sky130_fd_sc_hd__xor2_1
XU$$3038 net1509 net514 net1500 net787 VGND VGND VPWR VPWR t$5958 sky130_fd_sc_hd__a22o_1
XFILLER_35_818 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2304 net1639 net574 net1631 net847 VGND VGND VPWR VPWR t$5582 sky130_fd_sc_hd__a22o_1
XU$$3049 t$5963 net1358 VGND VGND VPWR VPWR booth_b44_m14 sky130_fd_sc_hd__xor2_1
XFILLER_75_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2315 t$5587 net1436 VGND VGND VPWR VPWR booth_b32_m58 sky130_fd_sc_hd__xor2_1
XU$$2326 net124 net575 net1774 net848 VGND VGND VPWR VPWR t$5593 sky130_fd_sc_hd__a22o_1
XFILLER_46_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2337 net1232 net563 net1126 net836 VGND VGND VPWR VPWR t$5600 sky130_fd_sc_hd__a22o_1
XU$$2348 t$5605 net1421 VGND VGND VPWR VPWR booth_b34_m6 sky130_fd_sc_hd__xor2_1
XU$$1603 net1727 net618 net1719 net891 VGND VGND VPWR VPWR t$5224 sky130_fd_sc_hd__a22o_1
XU$$1614 t$5229 net1483 VGND VGND VPWR VPWR booth_b22_m50 sky130_fd_sc_hd__xor2_1
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2359 net1213 net560 net1202 net833 VGND VGND VPWR VPWR t$5611 sky130_fd_sc_hd__a22o_1
XU$$1625 net1614 net616 net1606 net889 VGND VGND VPWR VPWR t$5235 sky130_fd_sc_hd__a22o_1
XFILLER_90_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1636 t$5240 net1481 VGND VGND VPWR VPWR booth_b22_m61 sky130_fd_sc_hd__xor2_1
XU$$1647 net1471 notblock$5245\[1\] VGND VGND VPWR VPWR t$5246 sky130_fd_sc_hd__and2_1
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1658 net932 net602 net1671 net875 VGND VGND VPWR VPWR t$5253 sky130_fd_sc_hd__a22o_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1669 t$5258 net1469 VGND VGND VPWR VPWR booth_b24_m9 sky130_fd_sc_hd__xor2_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0800_ clknet_leaf_123_clk booth_b40_m51 VGND VGND VPWR VPWR pp_row91_7 sky130_fd_sc_hd__dfxtp_1
X_1780_ clknet_leaf_222_clk booth_b30_m18 VGND VGND VPWR VPWR pp_row48_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_11_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0731_ clknet_leaf_135_clk booth_b44_m44 VGND VGND VPWR VPWR pp_row88_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_183_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0662_ clknet_leaf_172_clk booth_b56_m29 VGND VGND VPWR VPWR pp_row85_18 sky130_fd_sc_hd__dfxtp_1
X_2401_ clknet_leaf_74_clk booth_b56_m10 VGND VGND VPWR VPWR pp_row66_28 sky130_fd_sc_hd__dfxtp_1
X_0593_ clknet_leaf_186_clk booth_b28_m55 VGND VGND VPWR VPWR pp_row83_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_130_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2332_ clknet_leaf_100_clk booth_b64_m0 VGND VGND VPWR VPWR pp_row64_32 sky130_fd_sc_hd__dfxtp_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_61_3 c$544 s$547 s$549 VGND VGND VPWR VPWR c$1464 s$1465 sky130_fd_sc_hd__fa_1
X_2263_ clknet_leaf_230_clk booth_b6_m57 VGND VGND VPWR VPWR pp_row63_3 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_54_2 c$412 c$414 c$416 VGND VGND VPWR VPWR c$1378 s$1379 sky130_fd_sc_hd__fa_1
X_1214_ clknet_leaf_245_clk net171 VGND VGND VPWR VPWR pp_row22_13 sky130_fd_sc_hd__dfxtp_2
Xdadda_fa_5_31_1 s$2877 s$2879 s$2881 VGND VGND VPWR VPWR c$3522 s$3523 sky130_fd_sc_hd__fa_1
X_2194_ clknet_leaf_184_clk net139 VGND VGND VPWR VPWR pp_row109_11 sky130_fd_sc_hd__dfxtp_2
XU$$4240 net1549 net439 net1541 net721 VGND VGND VPWR VPWR t$6571 sky130_fd_sc_hd__a22o_1
XU$$4251 notblock$6575\[2\] net59 net1266 t$6576 notblock$6575\[0\] VGND VGND VPWR
+ VPWR sel_0$6577 sky130_fd_sc_hd__a32o_1
XU$$4262 t$6583 net1259 VGND VGND VPWR VPWR booth_b62_m4 sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_47_1 pp_row47_23 pp_row47_24 c$288 VGND VGND VPWR VPWR c$1292 s$1293 sky130_fd_sc_hd__fa_1
XFILLER_66_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4273 net1502 net418 net1222 net700 VGND VGND VPWR VPWR t$6589 sky130_fd_sc_hd__a22o_1
X_1145_ clknet_leaf_245_clk net165 VGND VGND VPWR VPWR pp_row17_9 sky130_fd_sc_hd__dfxtp_2
XFILLER_25_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4284 t$6594 net1258 VGND VGND VPWR VPWR booth_b62_m15 sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_24_0 c$2828 c$2830 c$2832 VGND VGND VPWR VPWR c$3492 s$3493 sky130_fd_sc_hd__fa_1
XU$$4295 net1119 net419 net1112 net701 VGND VGND VPWR VPWR t$6600 sky130_fd_sc_hd__a22o_1
XU$$3550 t$6218 net1334 VGND VGND VPWR VPWR booth_b50_m59 sky130_fd_sc_hd__xor2_1
XU$$3561 net1330 VGND VGND VPWR VPWR notsign$6224 sky130_fd_sc_hd__inv_1
XU$$3572 net1129 net480 net1037 net753 VGND VGND VPWR VPWR t$6231 sky130_fd_sc_hd__a22o_1
XFILLER_37_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3583 t$6236 net1319 VGND VGND VPWR VPWR booth_b52_m7 sky130_fd_sc_hd__xor2_1
X_1076_ clknet_leaf_52_clk booth_b0_m11 VGND VGND VPWR VPWR pp_row11_0 sky130_fd_sc_hd__dfxtp_1
XU$$3594 net1208 net480 net1200 net753 VGND VGND VPWR VPWR t$6242 sky130_fd_sc_hd__a22o_1
XU$$2860 net1609 net540 net1602 net813 VGND VGND VPWR VPWR t$5866 sky130_fd_sc_hd__a22o_1
XU$$2871 t$5871 net1383 VGND VGND VPWR VPWR booth_b40_m62 sky130_fd_sc_hd__xor2_1
XFILLER_179_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2882 net37 net1379 VGND VGND VPWR VPWR sel_1$5878 sky130_fd_sc_hd__xor2_4
XU$$2893 net1673 net519 net1562 net792 VGND VGND VPWR VPWR t$5884 sky130_fd_sc_hd__a22o_1
XFILLER_179_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1978_ clknet_leaf_72_clk net1304 VGND VGND VPWR VPWR pp_row54_28 sky130_fd_sc_hd__dfxtp_1
XFILLER_193_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_1053 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0929_ clknet_leaf_112_clk booth_b46_m51 VGND VGND VPWR VPWR pp_row97_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_107_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_69_2 s$2393 s$2395 s$2397 VGND VGND VPWR VPWR c$3108 s$3109 sky130_fd_sc_hd__fa_1
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$800 final_adder.p_new$848 final_adder.p_new$816 VGND VGND VPWR VPWR
+ final_adder.p_new$928 sky130_fd_sc_hd__and2_1
Xdadda_ha_1_36_1 pp_row36_3 pp_row36_4 VGND VGND VPWR VPWR c$210 s$211 sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$811 final_adder.p_new$826 final_adder.g_new$859 final_adder.g_new$827
+ VGND VGND VPWR VPWR final_adder.g_new$939 sky130_fd_sc_hd__a21o_1
XFILLER_69_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_39_0 s$3555 c$3972 s$3975 VGND VGND VPWR VPWR c$4230 s$4231 sky130_fd_sc_hd__fa_1
XFILLER_69_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$833 final_adder.p_new$848 final_adder.g_new$383 final_adder.g_new$849
+ VGND VGND VPWR VPWR final_adder.g_new$961 sky130_fd_sc_hd__a21o_2
Xfinal_adder.U$$855 final_adder.p_new$886 final_adder.g_new$951 final_adder.g_new$887
+ VGND VGND VPWR VPWR final_adder.g_new$983 sky130_fd_sc_hd__a21o_2
XFILLER_29_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$705 net1519 net402 net1513 net668 VGND VGND VPWR VPWR t$4766 sky130_fd_sc_hd__a22o_1
XFILLER_72_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$716 t$4771 net1415 VGND VGND VPWR VPWR booth_b10_m12 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$877 final_adder.p_new$908 final_adder.g_new$861 final_adder.g_new$909
+ VGND VGND VPWR VPWR final_adder.g_new$1005 sky130_fd_sc_hd__a21o_1
XU$$727 net1146 net401 net1138 net667 VGND VGND VPWR VPWR t$4777 sky130_fd_sc_hd__a22o_1
Xdadda_fa_1_42_0 pp_row42_0 pp_row42_1 pp_row42_2 VGND VGND VPWR VPWR c$244 s$245
+ sky130_fd_sc_hd__fa_1
XFILLER_16_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$738 t$4782 net1414 VGND VGND VPWR VPWR booth_b10_m23 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$899 final_adder.$signal$1214 final_adder.g_new$967 final_adder.$signal$250
+ VGND VGND VPWR VPWR final_adder.g_new$1027 sky130_fd_sc_hd__a21o_1
XU$$749 net1049 net406 net1041 net672 VGND VGND VPWR VPWR t$4788 sky130_fd_sc_hd__a22o_1
XFILLER_189_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_804 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_71_2 c$1576 s$1579 s$1581 VGND VGND VPWR VPWR c$2410 s$2411 sky130_fd_sc_hd__fa_1
Xfanout1000 net1001 VGND VGND VPWR VPWR net1000 sky130_fd_sc_hd__buf_4
XFILLER_156_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1011 net9 VGND VGND VPWR VPWR net1011 sky130_fd_sc_hd__buf_6
Xdadda_fa_3_64_1 c$1486 c$1488 c$1490 VGND VGND VPWR VPWR c$2352 s$2353 sky130_fd_sc_hd__fa_1
Xfanout1022 net89 VGND VGND VPWR VPWR net1022 sky130_fd_sc_hd__buf_8
Xfanout1033 net1034 VGND VGND VPWR VPWR net1033 sky130_fd_sc_hd__buf_2
XFILLER_0_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_41_0 c$3556 c$3558 s$3561 VGND VGND VPWR VPWR c$3978 s$3979 sky130_fd_sc_hd__fa_1
Xfanout1044 net1045 VGND VGND VPWR VPWR net1044 sky130_fd_sc_hd__buf_2
Xfanout1055 net1056 VGND VGND VPWR VPWR net1055 sky130_fd_sc_hd__buf_4
Xdadda_fa_3_57_0 s$491 c$1398 c$1400 VGND VGND VPWR VPWR c$2294 s$2295 sky130_fd_sc_hd__fa_1
Xfanout1066 net1067 VGND VGND VPWR VPWR net1066 sky130_fd_sc_hd__buf_4
Xfanout1077 net1078 VGND VGND VPWR VPWR net1077 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1088 net1093 VGND VGND VPWR VPWR net1088 sky130_fd_sc_hd__buf_4
XFILLER_19_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1099 net79 VGND VGND VPWR VPWR net1099 sky130_fd_sc_hd__buf_4
XFILLER_63_913 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2101 net1134 net580 net1117 net853 VGND VGND VPWR VPWR t$5479 sky130_fd_sc_hd__a22o_1
XFILLER_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2112 t$5484 net1442 VGND VGND VPWR VPWR booth_b30_m25 sky130_fd_sc_hd__xor2_1
XFILLER_47_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_100_2 s$2641 s$2643 s$2645 VGND VGND VPWR VPWR c$3294 s$3295 sky130_fd_sc_hd__fa_1
XFILLER_35_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2123 net1026 net582 net1018 net855 VGND VGND VPWR VPWR t$5490 sky130_fd_sc_hd__a22o_1
XU$$2134 t$5495 net1443 VGND VGND VPWR VPWR booth_b30_m36 sky130_fd_sc_hd__xor2_1
XU$$2145 net1746 net579 net1738 net852 VGND VGND VPWR VPWR t$5501 sky130_fd_sc_hd__a22o_1
XU$$1400 net1212 net629 net1203 net902 VGND VGND VPWR VPWR t$5121 sky130_fd_sc_hd__a22o_1
XU$$2156 t$5506 net1445 VGND VGND VPWR VPWR booth_b30_m47 sky130_fd_sc_hd__xor2_1
XU$$1411 t$5126 net1487 VGND VGND VPWR VPWR booth_b20_m17 sky130_fd_sc_hd__xor2_1
XU$$1422 net1097 net631 net1088 net904 VGND VGND VPWR VPWR t$5132 sky130_fd_sc_hd__a22o_1
XU$$2167 net1639 net578 net1631 net851 VGND VGND VPWR VPWR t$5512 sky130_fd_sc_hd__a22o_1
XU$$1433 t$5137 net1486 VGND VGND VPWR VPWR booth_b20_m28 sky130_fd_sc_hd__xor2_1
XFILLER_16_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2178 t$5517 net1446 VGND VGND VPWR VPWR booth_b30_m58 sky130_fd_sc_hd__xor2_1
XU$$2189 net1531 net582 net1772 net855 VGND VGND VPWR VPWR t$5523 sky130_fd_sc_hd__a22o_1
XU$$1444 net993 net630 net987 net903 VGND VGND VPWR VPWR t$5143 sky130_fd_sc_hd__a22o_1
XU$$1455 t$5148 net1490 VGND VGND VPWR VPWR booth_b20_m39 sky130_fd_sc_hd__xor2_1
XU$$1466 net1724 net634 net1715 net907 VGND VGND VPWR VPWR t$5154 sky130_fd_sc_hd__a22o_1
X_1901_ clknet_leaf_63_clk booth_b32_m20 VGND VGND VPWR VPWR pp_row52_16 sky130_fd_sc_hd__dfxtp_1
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1477 t$5159 net1493 VGND VGND VPWR VPWR booth_b20_m50 sky130_fd_sc_hd__xor2_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1488 net1612 net633 net1604 net906 VGND VGND VPWR VPWR t$5165 sky130_fd_sc_hd__a22o_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1499 t$5170 net1493 VGND VGND VPWR VPWR booth_b20_m61 sky130_fd_sc_hd__xor2_1
XFILLER_124_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1832_ clknet_leaf_18_clk booth_b18_m32 VGND VGND VPWR VPWR pp_row50_9 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_7_114_0 s$3855 c$4122 s$4125 VGND VGND VPWR VPWR c$4380 s$4381 sky130_fd_sc_hd__fa_1
X_1763_ clknet_leaf_235_clk net198 VGND VGND VPWR VPWR pp_row47_24 sky130_fd_sc_hd__dfxtp_1
XFILLER_129_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0714_ clknet_leaf_165_clk booth_b58_m29 VGND VGND VPWR VPWR pp_row87_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_183_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1694_ clknet_leaf_123_clk booth_b50_m56 VGND VGND VPWR VPWR pp_row106_5 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_79_1 s$3165 s$3167 s$3169 VGND VGND VPWR VPWR c$3714 s$3715 sky130_fd_sc_hd__fa_1
X_0645_ clknet_leaf_183_clk booth_b24_m61 VGND VGND VPWR VPWR pp_row85_2 sky130_fd_sc_hd__dfxtp_1
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0576_ clknet_leaf_189_clk booth_b48_m34 VGND VGND VPWR VPWR pp_row82_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2315_ clknet_leaf_30_clk booth_b34_m30 VGND VGND VPWR VPWR pp_row64_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_100_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$107 c$4364 s$4367 VGND VGND VPWR VPWR final_adder.$signal$216 final_adder.$signal$1197
+ sky130_fd_sc_hd__ha_1
XFILLER_111_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$118 c$4386 s$4389 VGND VGND VPWR VPWR final_adder.$signal$238 final_adder.$signal$1208
+ sky130_fd_sc_hd__ha_1
XFILLER_170_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2246_ clknet_leaf_30_clk booth_b44_m18 VGND VGND VPWR VPWR pp_row62_22 sky130_fd_sc_hd__dfxtp_1
XFILLER_39_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4070 t$6484 net1289 VGND VGND VPWR VPWR booth_b58_m45 sky130_fd_sc_hd__xor2_1
X_2177_ clknet_leaf_224_clk booth_b48_m12 VGND VGND VPWR VPWR pp_row60_24 sky130_fd_sc_hd__dfxtp_1
XFILLER_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4081 net1659 net453 net1651 net726 VGND VGND VPWR VPWR t$6490 sky130_fd_sc_hd__a22o_1
XU$$4092 t$6495 net1288 VGND VGND VPWR VPWR booth_b58_m56 sky130_fd_sc_hd__xor2_1
XFILLER_0_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1128_ clknet_leaf_12_clk booth_b8_m8 VGND VGND VPWR VPWR pp_row16_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_53_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3380 net1742 net498 net1734 net771 VGND VGND VPWR VPWR t$6132 sky130_fd_sc_hd__a22o_1
XFILLER_0_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3391 t$6137 net1344 VGND VGND VPWR VPWR booth_b48_m48 sky130_fd_sc_hd__xor2_1
XFILLER_20_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1059_ clknet_leaf_51_clk booth_b0_m9 VGND VGND VPWR VPWR pp_row9_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_179_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2690 t$5779 net1397 VGND VGND VPWR VPWR booth_b38_m40 sky130_fd_sc_hd__xor2_1
XFILLER_55_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_81_1 c$2482 c$2484 s$2487 VGND VGND VPWR VPWR c$3178 s$3179 sky130_fd_sc_hd__fa_1
XFILLER_162_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_74_0 s$1625 c$2422 c$2424 VGND VGND VPWR VPWR c$3134 s$3135 sky130_fd_sc_hd__fa_1
XFILLER_116_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput103 b[44] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__buf_2
XFILLER_163_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput114 b[54] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput125 b[6] VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__buf_4
XFILLER_0_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput136 c[106] VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput147 c[116] VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_1
XFILLER_56_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput158 c[126] VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput169 c[20] VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_1
XFILLER_186_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$630 final_adder.p_new$654 final_adder.p_new$638 VGND VGND VPWR VPWR
+ final_adder.p_new$758 sky130_fd_sc_hd__and2_1
XTAP_3912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$641 final_adder.p_new$648 final_adder.g_new$665 final_adder.g_new$649
+ VGND VGND VPWR VPWR final_adder.g_new$769 sky130_fd_sc_hd__a21o_1
XTAP_3923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$652 final_adder.p_new$676 final_adder.p_new$660 VGND VGND VPWR VPWR
+ final_adder.p_new$780 sky130_fd_sc_hd__and2_1
XTAP_3934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$502 t$4661 net1245 VGND VGND VPWR VPWR booth_b6_m42 sky130_fd_sc_hd__xor2_1
XFILLER_5_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$663 final_adder.p_new$670 final_adder.g_new$687 final_adder.g_new$671
+ VGND VGND VPWR VPWR final_adder.g_new$791 sky130_fd_sc_hd__a21o_1
XTAP_3945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$513 net1699 net430 net1691 net712 VGND VGND VPWR VPWR t$4667 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$674 final_adder.p_new$698 final_adder.p_new$682 VGND VGND VPWR VPWR
+ final_adder.p_new$802 sky130_fd_sc_hd__and2_1
XTAP_3956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$524 t$4672 net1247 VGND VGND VPWR VPWR booth_b6_m53 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$685 final_adder.p_new$692 final_adder.g_new$709 final_adder.g_new$693
+ VGND VGND VPWR VPWR final_adder.g_new$813 sky130_fd_sc_hd__a21o_1
XTAP_3967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$696 final_adder.p_new$720 final_adder.p_new$704 VGND VGND VPWR VPWR
+ final_adder.p_new$824 sky130_fd_sc_hd__and2_1
XU$$535 net1590 net432 net1582 net714 VGND VGND VPWR VPWR t$4678 sky130_fd_sc_hd__a22o_1
XTAP_3978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$546 t$4683 net1251 VGND VGND VPWR VPWR booth_b6_m64 sky130_fd_sc_hd__xor2_1
XTAP_3989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$557 t$4690 net1239 VGND VGND VPWR VPWR booth_b8_m1 sky130_fd_sc_hd__xor2_1
XFILLER_189_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$568 net1521 net415 net1513 net681 VGND VGND VPWR VPWR t$4696 sky130_fd_sc_hd__a22o_1
XU$$579 t$4701 net1239 VGND VGND VPWR VPWR booth_b8_m12 sky130_fd_sc_hd__xor2_1
XFILLER_32_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_798 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_89_0 c$3748 c$3750 s$3753 VGND VGND VPWR VPWR c$4074 s$4075 sky130_fd_sc_hd__fa_2
XFILLER_193_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0430_ clknet_leaf_207_clk booth_b46_m31 VGND VGND VPWR VPWR pp_row77_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_140_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0361_ clknet_leaf_204_clk booth_b34_m41 VGND VGND VPWR VPWR pp_row75_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_121_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2100_ clknet_leaf_32_clk booth_b36_m22 VGND VGND VPWR VPWR pp_row58_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_94_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0292_ clknet_leaf_199_clk booth_b24_m49 VGND VGND VPWR VPWR pp_row73_8 sky130_fd_sc_hd__dfxtp_1
X_2031_ clknet_leaf_72_clk booth_b34_m22 VGND VGND VPWR VPWR pp_row56_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_47_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_551 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1230 net1527 net649 net1756 net922 VGND VGND VPWR VPWR t$5033 sky130_fd_sc_hd__a22o_1
XFILLER_189_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1241 net1230 net637 net1123 net910 VGND VGND VPWR VPWR t$5040 sky130_fd_sc_hd__a22o_1
XU$$1252 t$5045 net1662 VGND VGND VPWR VPWR booth_b18_m6 sky130_fd_sc_hd__xor2_1
XU$$1263 net1210 net635 net1201 net908 VGND VGND VPWR VPWR t$5051 sky130_fd_sc_hd__a22o_1
XU$$1274 t$5056 net1665 VGND VGND VPWR VPWR booth_b18_m17 sky130_fd_sc_hd__xor2_1
XFILLER_149_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1285 net1097 net635 net1088 net908 VGND VGND VPWR VPWR t$5062 sky130_fd_sc_hd__a22o_1
XFILLER_149_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1296 t$5067 net1663 VGND VGND VPWR VPWR booth_b18_m28 sky130_fd_sc_hd__xor2_1
XFILLER_149_848 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1815_ clknet_leaf_25_clk booth_b40_m9 VGND VGND VPWR VPWR pp_row49_20 sky130_fd_sc_hd__dfxtp_1
XFILLER_191_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_91_0 c$3230 c$3232 c$3234 VGND VGND VPWR VPWR c$3760 s$3761 sky130_fd_sc_hd__fa_1
XFILLER_163_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1746_ clknet_leaf_234_clk booth_b18_m29 VGND VGND VPWR VPWR pp_row47_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_117_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_929 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1677_ clknet_leaf_22_clk booth_b44_m0 VGND VGND VPWR VPWR pp_row44_22 sky130_fd_sc_hd__dfxtp_1
XFILLER_117_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0628_ clknet_leaf_179_clk booth_b42_m42 VGND VGND VPWR VPWR pp_row84_12 sky130_fd_sc_hd__dfxtp_1
Xfanout804 net805 VGND VGND VPWR VPWR net804 sky130_fd_sc_hd__buf_4
Xfanout815 sel_1$5808 VGND VGND VPWR VPWR net815 sky130_fd_sc_hd__buf_8
Xdadda_fa_1_76_6 pp_row76_23 pp_row76_24 pp_row76_25 VGND VGND VPWR VPWR c$828 s$829
+ sky130_fd_sc_hd__fa_1
Xfanout826 net832 VGND VGND VPWR VPWR net826 sky130_fd_sc_hd__buf_4
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout837 net841 VGND VGND VPWR VPWR net837 sky130_fd_sc_hd__buf_4
Xfanout848 sel_1$5528 VGND VGND VPWR VPWR net848 sky130_fd_sc_hd__buf_6
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0559_ clknet_leaf_195_clk net236 VGND VGND VPWR VPWR pp_row81_25 sky130_fd_sc_hd__dfxtp_2
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout859 net865 VGND VGND VPWR VPWR net859 sky130_fd_sc_hd__buf_4
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_69_5 pp_row69_30 pp_row69_31 c$132 VGND VGND VPWR VPWR c$700 s$701 sky130_fd_sc_hd__fa_1
XFILLER_140_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2229_ clknet_leaf_229_clk booth_b12_m50 VGND VGND VPWR VPWR pp_row62_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_85_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_208 net1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_219 net1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_1_96_0 net1916 pp_row96_1 VGND VGND VPWR VPWR c$1048 s$1049 sky130_fd_sc_hd__ha_1
XFILLER_107_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_100_1 c$1914 c$1916 c$1918 VGND VGND VPWR VPWR c$2640 s$2641 sky130_fd_sc_hd__fa_1
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1060 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_121_0 c$3876 c$3878 s$3881 VGND VGND VPWR VPWR c$4138 s$4139 sky130_fd_sc_hd__fa_1
XFILLER_27_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_0_64_4 pp_row64_12 pp_row64_13 pp_row64_14 VGND VGND VPWR VPWR c$92 s$93
+ sky130_fd_sc_hd__fa_1
XFILLER_67_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_41_3 s$1223 s$1225 s$1227 VGND VGND VPWR VPWR c$2172 s$2173 sky130_fd_sc_hd__fa_1
XTAP_3720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$460 final_adder.p_new$466 final_adder.p_new$462 VGND VGND VPWR VPWR
+ final_adder.p_new$588 sky130_fd_sc_hd__and2_1
XTAP_3742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$310 net1179 net532 net1166 net805 VGND VGND VPWR VPWR t$4564 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$471 final_adder.p_new$472 final_adder.g_new$477 final_adder.g_new$473
+ VGND VGND VPWR VPWR final_adder.g_new$599 sky130_fd_sc_hd__a21o_1
XTAP_3753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$321 t$4569 net1274 VGND VGND VPWR VPWR booth_b4_m20 sky130_fd_sc_hd__xor2_1
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_34_2 c$1132 s$1135 s$1137 VGND VGND VPWR VPWR c$2114 s$2115 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$482 final_adder.p_new$488 final_adder.p_new$484 VGND VGND VPWR VPWR
+ final_adder.p_new$610 sky130_fd_sc_hd__and2_1
XFILLER_45_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$332 net1071 net527 net1063 net800 VGND VGND VPWR VPWR t$4575 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$493 final_adder.p_new$494 final_adder.g_new$499 final_adder.g_new$495
+ VGND VGND VPWR VPWR final_adder.g_new$621 sky130_fd_sc_hd__a21o_1
XTAP_3775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$343 t$4580 net1278 VGND VGND VPWR VPWR booth_b4_m31 sky130_fd_sc_hd__xor2_1
XTAP_3786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$354 net964 net527 net956 net800 VGND VGND VPWR VPWR t$4586 sky130_fd_sc_hd__a22o_1
XTAP_3797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_916 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$365 t$4591 net1274 VGND VGND VPWR VPWR booth_b4_m42 sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_27_1 pp_row27_11 pp_row27_12 pp_row27_13 VGND VGND VPWR VPWR c$2056 s$2057
+ sky130_fd_sc_hd__fa_1
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$376 net1699 net533 net1690 net806 VGND VGND VPWR VPWR t$4597 sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_192_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_192_clk
+ sky130_fd_sc_hd__clkbuf_16
XU$$387 t$4602 net1280 VGND VGND VPWR VPWR booth_b4_m53 sky130_fd_sc_hd__xor2_1
XU$$398 net1586 net529 net1578 net802 VGND VGND VPWR VPWR t$4608 sky130_fd_sc_hd__a22o_1
XFILLER_38_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1600_ clknet_leaf_237_clk booth_b0_m42 VGND VGND VPWR VPWR pp_row42_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_126_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1531_ clknet_leaf_44_clk booth_b6_m33 VGND VGND VPWR VPWR pp_row39_3 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_86_5 s$983 s$985 s$987 VGND VGND VPWR VPWR c$1768 s$1769 sky130_fd_sc_hd__fa_2
X_1462_ clknet_leaf_41_clk booth_b8_m28 VGND VGND VPWR VPWR pp_row36_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_141_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_79_4 s$875 s$877 s$879 VGND VGND VPWR VPWR c$1682 s$1683 sky130_fd_sc_hd__fa_1
X_0413_ clknet_leaf_192_clk booth_b14_m63 VGND VGND VPWR VPWR pp_row77_1 sky130_fd_sc_hd__dfxtp_1
X_1393_ clknet_leaf_110_clk booth_b50_m54 VGND VGND VPWR VPWR pp_row104_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_122_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0344_ clknet_leaf_129_clk booth_b52_m62 VGND VGND VPWR VPWR pp_row114_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_110_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0275_ clknet_leaf_217_clk booth_b56_m16 VGND VGND VPWR VPWR pp_row72_25 sky130_fd_sc_hd__dfxtp_1
X_2014_ clknet_leaf_81_clk booth_b4_m52 VGND VGND VPWR VPWR pp_row56_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_24_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_183_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_183_clk
+ sky130_fd_sc_hd__clkbuf_16
XU$$1060 t$4946 net1190 VGND VGND VPWR VPWR booth_b14_m47 sky130_fd_sc_hd__xor2_1
XU$$1071 net1641 net392 net1633 net658 VGND VGND VPWR VPWR t$4952 sky130_fd_sc_hd__a22o_1
XFILLER_10_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1082 t$4957 net1189 VGND VGND VPWR VPWR booth_b14_m58 sky130_fd_sc_hd__xor2_1
XU$$1093 net1530 net390 net1754 net656 VGND VGND VPWR VPWR t$4963 sky130_fd_sc_hd__a22o_1
XU$$3157_1789 VGND VGND VPWR VPWR U$$3157_1789/HI net1789 sky130_fd_sc_hd__conb_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_116_1 s$3387 s$3389 s$3391 VGND VGND VPWR VPWR c$3862 s$3863 sky130_fd_sc_hd__fa_1
XFILLER_192_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_109_0 c$3338 c$3340 c$3342 VGND VGND VPWR VPWR c$3832 s$3833 sky130_fd_sc_hd__fa_1
XFILLER_3_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1729_ clknet_leaf_21_clk booth_b38_m8 VGND VGND VPWR VPWR pp_row46_19 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_81_4 pp_row81_12 pp_row81_13 pp_row81_14 VGND VGND VPWR VPWR c$914 s$915
+ sky130_fd_sc_hd__fa_1
XFILLER_137_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout601 sel_0$5317 VGND VGND VPWR VPWR net601 sky130_fd_sc_hd__buf_6
Xfanout612 sel_0$5177 VGND VGND VPWR VPWR net612 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_74_3 pp_row74_17 pp_row74_18 pp_row74_19 VGND VGND VPWR VPWR c$786 s$787
+ sky130_fd_sc_hd__fa_1
Xfanout623 net625 VGND VGND VPWR VPWR net623 sky130_fd_sc_hd__clkbuf_4
Xfanout634 sel_0$5107 VGND VGND VPWR VPWR net634 sky130_fd_sc_hd__buf_6
XFILLER_86_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout645 net646 VGND VGND VPWR VPWR net645 sky130_fd_sc_hd__clkbuf_8
Xfanout656 net657 VGND VGND VPWR VPWR net656 sky130_fd_sc_hd__clkbuf_8
Xdadda_fa_4_51_2 s$2249 s$2251 s$2253 VGND VGND VPWR VPWR c$3000 s$3001 sky130_fd_sc_hd__fa_1
Xfanout667 net668 VGND VGND VPWR VPWR net667 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_67_2 pp_row67_24 pp_row67_25 pp_row67_26 VGND VGND VPWR VPWR c$658 s$659
+ sky130_fd_sc_hd__fa_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout678 net683 VGND VGND VPWR VPWR net678 sky130_fd_sc_hd__buf_4
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout689 net691 VGND VGND VPWR VPWR net689 sky130_fd_sc_hd__buf_2
Xdadda_fa_4_44_1 c$2186 c$2188 s$2191 VGND VGND VPWR VPWR c$2956 s$2957 sky130_fd_sc_hd__fa_1
XTAP_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_21_0 s$3483 c$3936 s$3939 VGND VGND VPWR VPWR c$4194 s$4195 sky130_fd_sc_hd__fa_1
XTAP_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_37_0 s$1181 c$2126 c$2128 VGND VGND VPWR VPWR c$2912 s$2913 sky130_fd_sc_hd__fa_1
XTAP_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_174_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_174_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1078 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_0_70_4 pp_row70_12 pp_row70_13 VGND VGND VPWR VPWR c$162 s$163 sky130_fd_sc_hd__ha_1
Xdadda_fa_3_89_3 s$1799 s$1801 s$1803 VGND VGND VPWR VPWR c$2556 s$2557 sky130_fd_sc_hd__fa_1
XFILLER_108_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_0_56_2 pp_row56_6 pp_row56_7 VGND VGND VPWR VPWR c$16 s$17 sky130_fd_sc_hd__ha_1
XFILLER_190_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_0_62_1 pp_row62_3 pp_row62_4 pp_row62_5 VGND VGND VPWR VPWR c$62 s$63 sky130_fd_sc_hd__fa_1
XFILLER_49_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3902 net1044 net463 net1028 net736 VGND VGND VPWR VPWR t$6399 sky130_fd_sc_hd__a22o_1
XFILLER_65_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3913 t$6404 net1299 VGND VGND VPWR VPWR booth_b56_m35 sky130_fd_sc_hd__xor2_1
Xdadda_fa_0_55_0 pp_row55_0 pp_row55_1 pp_row55_2 VGND VGND VPWR VPWR c$8 s$9 sky130_fd_sc_hd__fa_1
XU$$3924 net929 net465 net1750 net738 VGND VGND VPWR VPWR t$6410 sky130_fd_sc_hd__a22o_1
XTAP_4273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3935 t$6415 net1298 VGND VGND VPWR VPWR booth_b56_m46 sky130_fd_sc_hd__xor2_1
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3946 net1651 net462 net1643 net735 VGND VGND VPWR VPWR t$6421 sky130_fd_sc_hd__a22o_1
XTAP_4295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3957 t$6426 net1297 VGND VGND VPWR VPWR booth_b56_m57 sky130_fd_sc_hd__xor2_1
XTAP_3561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$290 final_adder.p_new$292 final_adder.p_new$290 VGND VGND VPWR VPWR
+ final_adder.p_new$418 sky130_fd_sc_hd__and2_1
XTAP_3572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$140 net1387 notblock$4475\[1\] VGND VGND VPWR VPWR t$4476 sky130_fd_sc_hd__and2_1
XFILLER_91_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3968 net1541 net463 net1533 net736 VGND VGND VPWR VPWR t$6432 sky130_fd_sc_hd__a22o_1
XU$$151 net937 net624 net1675 net897 VGND VGND VPWR VPWR t$4483 sky130_fd_sc_hd__a22o_1
XU$$3979 net1801 net455 net1233 net728 VGND VGND VPWR VPWR t$6439 sky130_fd_sc_hd__a22o_1
XTAP_3583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_165_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_165_clk
+ sky130_fd_sc_hd__clkbuf_16
XU$$162 t$4488 net1390 VGND VGND VPWR VPWR booth_b2_m9 sky130_fd_sc_hd__xor2_1
XU$$173 net1175 net620 net1166 net893 VGND VGND VPWR VPWR t$4494 sky130_fd_sc_hd__a22o_1
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$184 t$4499 net1389 VGND VGND VPWR VPWR booth_b2_m20 sky130_fd_sc_hd__xor2_1
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$195 net1071 net619 net1063 net892 VGND VGND VPWR VPWR t$4505 sky130_fd_sc_hd__a22o_1
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0962_ clknet_leaf_114_clk booth_b36_m63 VGND VGND VPWR VPWR pp_row99_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_192_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0893_ clknet_leaf_101_clk booth_b52_m43 VGND VGND VPWR VPWR pp_row95_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_146_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_91_3 pp_row91_18 pp_row91_19 pp_row91_20 VGND VGND VPWR VPWR c$1824 s$1825
+ sky130_fd_sc_hd__fa_1
XFILLER_160_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_84_2 c$940 c$942 c$944 VGND VGND VPWR VPWR c$1738 s$1739 sky130_fd_sc_hd__fa_1
X_1514_ clknet_leaf_17_clk booth_b20_m18 VGND VGND VPWR VPWR pp_row38_10 sky130_fd_sc_hd__dfxtp_1
Xoutput259 net259 VGND VGND VPWR VPWR o[101] sky130_fd_sc_hd__buf_2
XFILLER_99_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2494_ clknet_leaf_142_clk booth_b28_m41 VGND VGND VPWR VPWR pp_row69_12 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_61_1 s$3057 s$3059 s$3061 VGND VGND VPWR VPWR c$3642 s$3643 sky130_fd_sc_hd__fa_1
Xdadda_fa_2_77_1 c$820 c$822 c$824 VGND VGND VPWR VPWR c$1652 s$1653 sky130_fd_sc_hd__fa_1
X_1445_ clknet_leaf_65_clk booth_b16_m19 VGND VGND VPWR VPWR pp_row35_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_114_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_54_0 c$3008 c$3010 c$3012 VGND VGND VPWR VPWR c$3612 s$3613 sky130_fd_sc_hd__fa_1
XFILLER_68_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1376_ clknet_leaf_7_clk booth_b8_m24 VGND VGND VPWR VPWR pp_row32_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_114_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_53_8 pp_row53_26 pp_row53_27 c$1 VGND VGND VPWR VPWR c$418 s$419 sky130_fd_sc_hd__fa_1
X_0327_ clknet_leaf_227_clk booth_b30_m44 VGND VGND VPWR VPWR pp_row74_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_55_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0258_ clknet_leaf_211_clk booth_b24_m48 VGND VGND VPWR VPWR pp_row72_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_36_551 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_156_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_156_clk
+ sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_2_100_0 net1904 pp_row100_1 pp_row100_2 VGND VGND VPWR VPWR c$1924 s$1925
+ sky130_fd_sc_hd__fa_1
X_0189_ clknet_leaf_180_clk booth_b62_m50 VGND VGND VPWR VPWR pp_row112_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_24_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_913 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_99_2 s$2633 s$2635 s$2637 VGND VGND VPWR VPWR c$3288 s$3289 sky130_fd_sc_hd__fa_1
XFILLER_178_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_810 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_69_0 s$3675 c$4032 s$4035 VGND VGND VPWR VPWR c$4290 s$4291 sky130_fd_sc_hd__fa_1
Xfanout1407 net31 VGND VGND VPWR VPWR net1407 sky130_fd_sc_hd__clkbuf_4
XFILLER_160_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1418 net1419 VGND VGND VPWR VPWR net1418 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_72_0 pp_row72_11 pp_row72_12 pp_row72_13 VGND VGND VPWR VPWR c$744 s$745
+ sky130_fd_sc_hd__fa_1
Xfanout420 net421 VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__buf_4
Xfanout431 net433 VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__buf_4
Xfanout1429 net29 VGND VGND VPWR VPWR net1429 sky130_fd_sc_hd__buf_8
XFILLER_87_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout442 net450 VGND VGND VPWR VPWR net442 sky130_fd_sc_hd__buf_4
XFILLER_63_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout453 net454 VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__buf_4
XFILLER_115_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_559 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout464 net467 VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__clkbuf_8
XFILLER_87_974 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout475 sel_0$6297 VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__buf_6
XFILLER_150_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout486 net487 VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__clkbuf_4
XFILLER_171_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout497 net500 VGND VGND VPWR VPWR net497 sky130_fd_sc_hd__buf_4
XFILLER_46_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3209 net1073 net501 net1065 net774 VGND VGND VPWR VPWR t$6045 sky130_fd_sc_hd__a22o_1
XFILLER_74_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2508 net1149 net554 net1144 net827 VGND VGND VPWR VPWR t$5687 sky130_fd_sc_hd__a22o_1
XFILLER_74_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2519 t$5692 net1404 VGND VGND VPWR VPWR booth_b36_m23 sky130_fd_sc_hd__xor2_1
XFILLER_61_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1807 net1499 net596 net1224 net869 VGND VGND VPWR VPWR t$5329 sky130_fd_sc_hd__a22o_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_147_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_147_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1818 t$5334 net1457 VGND VGND VPWR VPWR booth_b26_m15 sky130_fd_sc_hd__xor2_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1829 net1116 net595 net1107 net868 VGND VGND VPWR VPWR t$5340 sky130_fd_sc_hd__a22o_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_94_1 c$1846 c$1848 c$1850 VGND VGND VPWR VPWR c$2592 s$2593 sky130_fd_sc_hd__fa_2
XFILLER_7_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_71_0 c$3676 c$3678 s$3681 VGND VGND VPWR VPWR c$4038 s$4039 sky130_fd_sc_hd__fa_1
XFILLER_170_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_87_0 s$999 c$1758 c$1760 VGND VGND VPWR VPWR c$2534 s$2535 sky130_fd_sc_hd__fa_1
XFILLER_151_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1230_ clknet_leaf_12_clk booth_b0_m24 VGND VGND VPWR VPWR pp_row24_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_111_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4400 net1677 sel_0$6647 net1566 net696 VGND VGND VPWR VPWR t$6654 sky130_fd_sc_hd__a22o_1
XU$$4411 t$6659 net1826 VGND VGND VPWR VPWR booth_b64_m10 sky130_fd_sc_hd__xor2_1
XU$$4422 net1169 sel_0$6647 net1160 net695 VGND VGND VPWR VPWR t$6665 sky130_fd_sc_hd__a22o_1
XFILLER_77_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4433 t$6670 net1837 VGND VGND VPWR VPWR booth_b64_m21 sky130_fd_sc_hd__xor2_1
XFILLER_65_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1161_ clknet_leaf_46_clk booth_b2_m17 VGND VGND VPWR VPWR pp_row19_1 sky130_fd_sc_hd__dfxtp_1
XU$$4444 net1070 sel_0$6647 net1062 net698 VGND VGND VPWR VPWR t$6676 sky130_fd_sc_hd__a22o_1
XFILLER_37_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4455 t$6681 net1848 VGND VGND VPWR VPWR booth_b64_m32 sky130_fd_sc_hd__xor2_1
XFILLER_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3710 t$6301 net1305 VGND VGND VPWR VPWR booth_b54_m2 sky130_fd_sc_hd__xor2_1
XU$$4466 net963 sel_0$6647 net953 net697 VGND VGND VPWR VPWR t$6687 sky130_fd_sc_hd__a22o_1
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_49_5 s$341 s$343 s$345 VGND VGND VPWR VPWR c$1324 s$1325 sky130_fd_sc_hd__fa_1
XU$$3721 net1514 net471 net1507 net744 VGND VGND VPWR VPWR t$6307 sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_116_0 pp_row116_2 pp_row116_3 pp_row116_4 VGND VGND VPWR VPWR c$3386 s$3387
+ sky130_fd_sc_hd__fa_1
XTAP_4070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3732 t$6312 net1304 VGND VGND VPWR VPWR booth_b54_m13 sky130_fd_sc_hd__xor2_1
XFILLER_92_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4477 t$6692 net1859 VGND VGND VPWR VPWR booth_b64_m43 sky130_fd_sc_hd__xor2_1
X_1092_ clknet_leaf_248_clk net160 VGND VGND VPWR VPWR pp_row12_8 sky130_fd_sc_hd__dfxtp_2
XU$$3743 net1141 net468 net1136 net741 VGND VGND VPWR VPWR t$6318 sky130_fd_sc_hd__a22o_1
XU$$4488 net1694 sel_0$6647 net1685 net696 VGND VGND VPWR VPWR t$6698 sky130_fd_sc_hd__a22o_1
XTAP_4092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3754 t$6323 net1300 VGND VGND VPWR VPWR booth_b54_m24 sky130_fd_sc_hd__xor2_1
XU$$4499 t$6703 net1870 VGND VGND VPWR VPWR booth_b64_m54 sky130_fd_sc_hd__xor2_1
XU$$3765 net1044 net469 net1028 net742 VGND VGND VPWR VPWR t$6329 sky130_fd_sc_hd__a22o_1
XU$$3776 t$6334 net1301 VGND VGND VPWR VPWR booth_b54_m35 sky130_fd_sc_hd__xor2_1
XFILLER_46_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_138_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_138_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3787 net928 net472 net1749 net745 VGND VGND VPWR VPWR t$6340 sky130_fd_sc_hd__a22o_1
XTAP_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3798 t$6345 net1307 VGND VGND VPWR VPWR booth_b54_m46 sky130_fd_sc_hd__xor2_1
XFILLER_178_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_380 net1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_391 net1530 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1994_ clknet_leaf_143_clk booth_b54_m54 VGND VGND VPWR VPWR pp_row108_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_193_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_913 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0945_ clknet_leaf_113_clk booth_b38_m60 VGND VGND VPWR VPWR pp_row98_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_186_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0876_ clknet_leaf_93_clk booth_b60_m34 VGND VGND VPWR VPWR pp_row94_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_146_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2477_ clknet_leaf_99_clk booth_b62_m6 VGND VGND VPWR VPWR pp_row68_30 sky130_fd_sc_hd__dfxtp_1
XFILLER_88_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1428_ clknet_leaf_121_clk booth_b56_m48 VGND VGND VPWR VPWR pp_row104_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_68_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_ha_4_122_0_1919 VGND VGND VPWR VPWR net1919 dadda_ha_4_122_0_1919/LO sky130_fd_sc_hd__conb_1
Xdadda_fa_1_51_5 pp_row51_15 pp_row51_16 pp_row51_17 VGND VGND VPWR VPWR c$376 s$377
+ sky130_fd_sc_hd__fa_1
X_1359_ clknet_leaf_10_clk booth_b12_m19 VGND VGND VPWR VPWR pp_row31_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_18_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$909 t$4869 net1314 VGND VGND VPWR VPWR booth_b12_m40 sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_44_4 pp_row44_12 pp_row44_13 pp_row44_14 VGND VGND VPWR VPWR c$272 s$273
+ sky130_fd_sc_hd__fa_1
XFILLER_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_129_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_129_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_70_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_14_2 pp_row14_8 pp_row14_9 s$1975 VGND VGND VPWR VPWR c$2778 s$2779 sky130_fd_sc_hd__fa_1
XFILLER_52_896 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1204 net1209 VGND VGND VPWR VPWR net1204 sky130_fd_sc_hd__clkbuf_4
Xfanout1215 net67 VGND VGND VPWR VPWR net1215 sky130_fd_sc_hd__clkbuf_4
Xfanout1226 net66 VGND VGND VPWR VPWR net1226 sky130_fd_sc_hd__buf_6
Xfanout1237 net1238 VGND VGND VPWR VPWR net1237 sky130_fd_sc_hd__buf_6
XFILLER_94_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1248 net1249 VGND VGND VPWR VPWR net1248 sky130_fd_sc_hd__buf_4
Xfanout1259 net1262 VGND VGND VPWR VPWR net1259 sky130_fd_sc_hd__buf_6
XFILLER_8_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3006 t$5940 net1374 VGND VGND VPWR VPWR booth_b42_m61 sky130_fd_sc_hd__xor2_1
XU$$3017 net1359 notblock$5945\[1\] VGND VGND VPWR VPWR t$5946 sky130_fd_sc_hd__and2_1
XFILLER_75_966 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4385_1810 VGND VGND VPWR VPWR U$$4385_1810/HI net1810 sky130_fd_sc_hd__conb_1
XU$$3028 net935 net510 net1673 net783 VGND VGND VPWR VPWR t$5953 sky130_fd_sc_hd__a22o_1
XU$$3039 t$5958 net1362 VGND VGND VPWR VPWR booth_b44_m9 sky130_fd_sc_hd__xor2_1
XFILLER_19_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_903 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2305 t$5582 net1436 VGND VGND VPWR VPWR booth_b32_m53 sky130_fd_sc_hd__xor2_1
XFILLER_62_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2316 net1590 net575 net1582 net848 VGND VGND VPWR VPWR t$5588 sky130_fd_sc_hd__a22o_1
XFILLER_90_936 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2327 t$5593 net1437 VGND VGND VPWR VPWR booth_b32_m64 sky130_fd_sc_hd__xor2_1
XU$$2338 t$5600 net1423 VGND VGND VPWR VPWR booth_b34_m1 sky130_fd_sc_hd__xor2_1
XU$$2349 net1519 net560 net1511 net833 VGND VGND VPWR VPWR t$5606 sky130_fd_sc_hd__a22o_1
XU$$1604 t$5224 net1484 VGND VGND VPWR VPWR booth_b22_m45 sky130_fd_sc_hd__xor2_1
XU$$1615 net1654 net616 net1646 net889 VGND VGND VPWR VPWR t$5230 sky130_fd_sc_hd__a22o_1
XU$$1626 t$5235 net1483 VGND VGND VPWR VPWR booth_b22_m56 sky130_fd_sc_hd__xor2_1
XFILLER_188_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1637 net1544 net617 net1536 net890 VGND VGND VPWR VPWR t$5241 sky130_fd_sc_hd__a22o_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1648 notblock$5245\[2\] net17 net1482 t$5246 notblock$5245\[0\] VGND VGND VPWR
+ VPWR sel_0$5247 sky130_fd_sc_hd__a32o_4
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1659 t$5253 net1466 VGND VGND VPWR VPWR booth_b24_m4 sky130_fd_sc_hd__xor2_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_913 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0730_ clknet_leaf_135_clk booth_b42_m46 VGND VGND VPWR VPWR pp_row88_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_155_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0661_ clknet_leaf_176_clk booth_b54_m31 VGND VGND VPWR VPWR pp_row85_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_7_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1028 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2400_ clknet_leaf_74_clk booth_b54_m12 VGND VGND VPWR VPWR pp_row66_27 sky130_fd_sc_hd__dfxtp_1
X_0592_ clknet_leaf_186_clk booth_b26_m57 VGND VGND VPWR VPWR pp_row83_4 sky130_fd_sc_hd__dfxtp_1
X_2331_ clknet_leaf_99_clk booth_b62_m2 VGND VGND VPWR VPWR pp_row64_31 sky130_fd_sc_hd__dfxtp_1
XFILLER_69_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2262_ clknet_leaf_230_clk booth_b4_m59 VGND VGND VPWR VPWR pp_row63_2 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_61_4 s$551 s$553 s$555 VGND VGND VPWR VPWR c$1466 s$1467 sky130_fd_sc_hd__fa_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_900 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1213_ clknet_leaf_49_clk net1478 VGND VGND VPWR VPWR pp_row22_12 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_54_3 c$418 s$421 s$423 VGND VGND VPWR VPWR c$1380 s$1381 sky130_fd_sc_hd__fa_1
X_2193_ clknet_leaf_227_clk booth_b12_m49 VGND VGND VPWR VPWR pp_row61_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_38_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4230 net1606 net435 net1598 net717 VGND VGND VPWR VPWR t$6566 sky130_fd_sc_hd__a22o_1
XU$$4241 t$6571 net1271 VGND VGND VPWR VPWR booth_b60_m62 sky130_fd_sc_hd__xor2_1
XU$$4252 net59 net1266 VGND VGND VPWR VPWR sel_1$6578 sky130_fd_sc_hd__xor2_2
XFILLER_168_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4263 net1678 net422 net1567 net704 VGND VGND VPWR VPWR t$6584 sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_47_2 c$290 c$292 c$294 VGND VGND VPWR VPWR c$1294 s$1295 sky130_fd_sc_hd__fa_1
X_1144_ clknet_leaf_11_clk booth_b16_m1 VGND VGND VPWR VPWR pp_row17_8 sky130_fd_sc_hd__dfxtp_1
XU$$4274 t$6589 net1254 VGND VGND VPWR VPWR booth_b62_m10 sky130_fd_sc_hd__xor2_1
XU$$3540 t$6213 net1335 VGND VGND VPWR VPWR booth_b50_m54 sky130_fd_sc_hd__xor2_1
XFILLER_19_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4285 net1169 net418 net1160 net700 VGND VGND VPWR VPWR t$6595 sky130_fd_sc_hd__a22o_1
XFILLER_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_24_1 s$2835 s$2837 s$2839 VGND VGND VPWR VPWR c$3494 s$3495 sky130_fd_sc_hd__fa_1
XU$$3551 net1583 net489 net1556 net762 VGND VGND VPWR VPWR t$6219 sky130_fd_sc_hd__a22o_1
XU$$4296 t$6600 net1255 VGND VGND VPWR VPWR booth_b62_m21 sky130_fd_sc_hd__xor2_1
XFILLER_168_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3562 net1330 VGND VGND VPWR VPWR notblock$6225\[0\] sky130_fd_sc_hd__inv_1
XU$$3573 t$6231 net1324 VGND VGND VPWR VPWR booth_b52_m2 sky130_fd_sc_hd__xor2_1
X_1075_ clknet_leaf_248_clk net140 VGND VGND VPWR VPWR pp_row10_7 sky130_fd_sc_hd__dfxtp_2
XU$$3584 net1514 net476 net1507 net749 VGND VGND VPWR VPWR t$6237 sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_17_0 c$2786 c$2788 c$2790 VGND VGND VPWR VPWR c$3464 s$3465 sky130_fd_sc_hd__fa_1
XU$$3595 t$6242 net1324 VGND VGND VPWR VPWR booth_b52_m13 sky130_fd_sc_hd__xor2_1
XU$$2850 net1652 net540 net1642 net813 VGND VGND VPWR VPWR t$5861 sky130_fd_sc_hd__a22o_1
XU$$2861 t$5866 net1382 VGND VGND VPWR VPWR booth_b40_m57 sky130_fd_sc_hd__xor2_1
XFILLER_178_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2872 net1540 net541 net1532 net814 VGND VGND VPWR VPWR t$5872 sky130_fd_sc_hd__a22o_1
XU$$2883 net1785 net519 net1227 net792 VGND VGND VPWR VPWR t$5879 sky130_fd_sc_hd__a22o_1
XU$$2894 t$5884 net1367 VGND VGND VPWR VPWR booth_b42_m5 sky130_fd_sc_hd__xor2_1
XFILLER_61_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1977_ clknet_leaf_72_clk booth_b54_m0 VGND VGND VPWR VPWR pp_row54_27 sky130_fd_sc_hd__dfxtp_1
XFILLER_159_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0928_ clknet_leaf_112_clk booth_b44_m53 VGND VGND VPWR VPWR pp_row97_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0859_ clknet_leaf_194_clk net249 VGND VGND VPWR VPWR pp_row93_19 sky130_fd_sc_hd__dfxtp_2
XFILLER_146_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$801 final_adder.p_new$816 final_adder.g_new$849 final_adder.g_new$817
+ VGND VGND VPWR VPWR final_adder.g_new$929 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$823 final_adder.p_new$838 final_adder.g_new$751 final_adder.g_new$839
+ VGND VGND VPWR VPWR final_adder.g_new$951 sky130_fd_sc_hd__a21o_2
XFILLER_21_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$845 final_adder.p_new$876 final_adder.g_new$941 final_adder.g_new$877
+ VGND VGND VPWR VPWR final_adder.g_new$973 sky130_fd_sc_hd__a21o_2
XU$$706 t$4766 net1412 VGND VGND VPWR VPWR booth_b10_m7 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$867 final_adder.p_new$898 final_adder.g_new$851 final_adder.g_new$899
+ VGND VGND VPWR VPWR final_adder.g_new$995 sky130_fd_sc_hd__a21o_2
XU$$717 net1204 net406 net1194 net672 VGND VGND VPWR VPWR t$4772 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$889 final_adder.p_new$920 final_adder.g_new$753 final_adder.g_new$921
+ VGND VGND VPWR VPWR final_adder.g_new$1017 sky130_fd_sc_hd__a21o_1
Xdadda_fa_1_42_1 pp_row42_3 pp_row42_4 pp_row42_5 VGND VGND VPWR VPWR c$246 s$247
+ sky130_fd_sc_hd__fa_1
XU$$728 t$4777 net1412 VGND VGND VPWR VPWR booth_b10_m18 sky130_fd_sc_hd__xor2_1
XU$$739 net1091 net405 net1083 net671 VGND VGND VPWR VPWR t$4783 sky130_fd_sc_hd__a22o_1
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_816 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_90_0_1901 VGND VGND VPWR VPWR net1901 dadda_fa_1_90_0_1901/LO sky130_fd_sc_hd__conb_1
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1050 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_71_3 s$1583 s$1585 s$1587 VGND VGND VPWR VPWR c$2412 s$2413 sky130_fd_sc_hd__fa_1
XFILLER_134_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1001 net1005 VGND VGND VPWR VPWR net1001 sky130_fd_sc_hd__buf_4
Xfanout1012 net1014 VGND VGND VPWR VPWR net1012 sky130_fd_sc_hd__buf_6
XFILLER_67_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_64_2 c$1492 s$1495 s$1497 VGND VGND VPWR VPWR c$2354 s$2355 sky130_fd_sc_hd__fa_1
XFILLER_0_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1023 net1024 VGND VGND VPWR VPWR net1023 sky130_fd_sc_hd__buf_4
Xfanout1034 net87 VGND VGND VPWR VPWR net1034 sky130_fd_sc_hd__buf_6
Xfanout1045 net1046 VGND VGND VPWR VPWR net1045 sky130_fd_sc_hd__buf_6
Xdadda_fa_3_57_1 c$1402 c$1404 c$1406 VGND VGND VPWR VPWR c$2296 s$2297 sky130_fd_sc_hd__fa_1
XFILLER_0_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1056 net1059 VGND VGND VPWR VPWR net1056 sky130_fd_sc_hd__buf_6
Xfanout1067 net83 VGND VGND VPWR VPWR net1067 sky130_fd_sc_hd__buf_4
XFILLER_86_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1078 net1079 VGND VGND VPWR VPWR net1078 sky130_fd_sc_hd__buf_6
Xfanout1089 net1093 VGND VGND VPWR VPWR net1089 sky130_fd_sc_hd__buf_2
Xdadda_fa_6_34_0 c$3528 c$3530 s$3533 VGND VGND VPWR VPWR c$3964 s$3965 sky130_fd_sc_hd__fa_1
XFILLER_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_988 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2102 t$5479 net1441 VGND VGND VPWR VPWR booth_b30_m20 sky130_fd_sc_hd__xor2_1
XU$$2113 net1075 net581 net1067 net854 VGND VGND VPWR VPWR t$5485 sky130_fd_sc_hd__a22o_1
XFILLER_74_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2124 t$5490 net1442 VGND VGND VPWR VPWR booth_b30_m31 sky130_fd_sc_hd__xor2_1
XU$$2135 net972 net582 net963 net855 VGND VGND VPWR VPWR t$5496 sky130_fd_sc_hd__a22o_1
XFILLER_63_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1401 t$5121 net1487 VGND VGND VPWR VPWR booth_b20_m12 sky130_fd_sc_hd__xor2_1
XU$$2146 t$5501 net1445 VGND VGND VPWR VPWR booth_b30_m42 sky130_fd_sc_hd__xor2_1
XU$$2157 net1696 net579 net1688 net852 VGND VGND VPWR VPWR t$5507 sky130_fd_sc_hd__a22o_1
XU$$1412 net1146 net629 net1139 net902 VGND VGND VPWR VPWR t$5127 sky130_fd_sc_hd__a22o_1
XU$$1423 t$5132 net1485 VGND VGND VPWR VPWR booth_b20_m23 sky130_fd_sc_hd__xor2_1
XU$$2168 t$5512 net1445 VGND VGND VPWR VPWR booth_b30_m53 sky130_fd_sc_hd__xor2_1
XFILLER_16_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1434 net1048 net628 net1040 net901 VGND VGND VPWR VPWR t$5138 sky130_fd_sc_hd__a22o_1
XU$$2179 net1589 net579 net1580 net852 VGND VGND VPWR VPWR t$5518 sky130_fd_sc_hd__a22o_1
XU$$1445 t$5143 net1489 VGND VGND VPWR VPWR booth_b20_m34 sky130_fd_sc_hd__xor2_1
XFILLER_43_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1456 net941 net632 net925 net905 VGND VGND VPWR VPWR t$5149 sky130_fd_sc_hd__a22o_1
XFILLER_188_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1900_ clknet_leaf_63_clk booth_b30_m22 VGND VGND VPWR VPWR pp_row52_15 sky130_fd_sc_hd__dfxtp_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1467 t$5154 net1493 VGND VGND VPWR VPWR booth_b20_m45 sky130_fd_sc_hd__xor2_1
XU$$1478 net1654 net632 net1646 net905 VGND VGND VPWR VPWR t$5160 sky130_fd_sc_hd__a22o_1
XFILLER_163_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1489 t$5165 net1492 VGND VGND VPWR VPWR booth_b20_m56 sky130_fd_sc_hd__xor2_1
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1831_ clknet_leaf_25_clk booth_b16_m34 VGND VGND VPWR VPWR pp_row50_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1762_ clknet_leaf_220_clk booth_b46_m1 VGND VGND VPWR VPWR pp_row47_23 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_107_0 s$3827 c$4108 s$4111 VGND VGND VPWR VPWR c$4366 s$4367 sky130_fd_sc_hd__fa_1
XFILLER_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0713_ clknet_leaf_165_clk booth_b56_m31 VGND VGND VPWR VPWR pp_row87_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_128_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1693_ clknet_leaf_18_clk booth_b24_m21 VGND VGND VPWR VPWR pp_row45_12 sky130_fd_sc_hd__dfxtp_1
X_0644_ clknet_leaf_164_clk booth_b56_m61 VGND VGND VPWR VPWR pp_row117_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_98_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0575_ clknet_leaf_189_clk booth_b46_m36 VGND VGND VPWR VPWR pp_row82_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_112_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2314_ clknet_leaf_30_clk booth_b32_m32 VGND VGND VPWR VPWR pp_row64_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_98_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$108 c$4366 s$4369 VGND VGND VPWR VPWR final_adder.$signal$218 final_adder.$signal$1198
+ sky130_fd_sc_hd__ha_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2245_ clknet_leaf_29_clk booth_b42_m20 VGND VGND VPWR VPWR pp_row62_21 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$119 c$4388 s$4391 VGND VGND VPWR VPWR final_adder.$signal$240 final_adder.$signal$1209
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_2_52_0 s c$366 c$368 VGND VGND VPWR VPWR c$1350 s$1351 sky130_fd_sc_hd__fa_1
XFILLER_85_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1590 net1593 VGND VGND VPWR VPWR net1590 sky130_fd_sc_hd__buf_6
XFILLER_54_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2176_ clknet_leaf_223_clk booth_b46_m14 VGND VGND VPWR VPWR pp_row60_23 sky130_fd_sc_hd__dfxtp_1
XFILLER_122_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4060 t$6479 net1289 VGND VGND VPWR VPWR booth_b58_m40 sky130_fd_sc_hd__xor2_1
XU$$4071 net1718 net457 net1709 net730 VGND VGND VPWR VPWR t$6485 sky130_fd_sc_hd__a22o_1
XU$$4082 t$6490 net1285 VGND VGND VPWR VPWR booth_b58_m51 sky130_fd_sc_hd__xor2_1
X_1127_ clknet_leaf_119_clk booth_b60_m42 VGND VGND VPWR VPWR pp_row102_12 sky130_fd_sc_hd__dfxtp_1
XU$$4093 net1610 net456 net1601 net729 VGND VGND VPWR VPWR t$6496 sky130_fd_sc_hd__a22o_1
XU$$3370 net959 net494 net950 net767 VGND VGND VPWR VPWR t$6127 sky130_fd_sc_hd__a22o_1
XU$$3381 t$6132 net1344 VGND VGND VPWR VPWR booth_b48_m43 sky130_fd_sc_hd__xor2_1
XU$$3392 net1693 net498 net1684 net771 VGND VGND VPWR VPWR t$6138 sky130_fd_sc_hd__a22o_1
XFILLER_94_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1058_ clknet_leaf_248_clk net245 VGND VGND VPWR VPWR pp_row8_6 sky130_fd_sc_hd__dfxtp_2
XFILLER_15_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_6_0 pp_row6_0 pp_row6_1 pp_row6_2 VGND VGND VPWR VPWR c$3420 s$3421 sky130_fd_sc_hd__fa_1
XFILLER_22_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2680 t$5774 net1394 VGND VGND VPWR VPWR booth_b38_m35 sky130_fd_sc_hd__xor2_1
XU$$2691 net926 net545 net1747 net818 VGND VGND VPWR VPWR t$5780 sky130_fd_sc_hd__a22o_1
XFILLER_179_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_60_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_60_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_21_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1990 net1001 net591 net996 net864 VGND VGND VPWR VPWR t$5422 sky130_fd_sc_hd__a22o_1
XFILLER_22_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_81_2 s$2489 s$2491 s$2493 VGND VGND VPWR VPWR c$3180 s$3181 sky130_fd_sc_hd__fa_1
XFILLER_162_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_74_1 c$2426 c$2428 s$2431 VGND VGND VPWR VPWR c$3136 s$3137 sky130_fd_sc_hd__fa_1
XFILLER_134_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_7_51_0 s$3603 c$3996 s$3999 VGND VGND VPWR VPWR c$4254 s$4255 sky130_fd_sc_hd__fa_2
Xdadda_fa_4_67_0 s$1541 c$2366 c$2368 VGND VGND VPWR VPWR c$3092 s$3093 sky130_fd_sc_hd__fa_1
Xinput104 b[45] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__buf_6
Xinput115 b[55] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__buf_2
XFILLER_163_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput126 b[7] VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_2
Xinput137 c[107] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_1
Xinput148 c[117] VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_1
Xinput159 c[127] VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_1
XFILLER_130_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$631 final_adder.p_new$638 final_adder.g_new$655 final_adder.g_new$639
+ VGND VGND VPWR VPWR final_adder.g_new$759 sky130_fd_sc_hd__a21o_1
XTAP_3913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$642 final_adder.p_new$666 final_adder.p_new$650 VGND VGND VPWR VPWR
+ final_adder.p_new$770 sky130_fd_sc_hd__and2_1
XTAP_3924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$653 final_adder.p_new$660 final_adder.g_new$677 final_adder.g_new$661
+ VGND VGND VPWR VPWR final_adder.g_new$781 sky130_fd_sc_hd__a21o_1
XTAP_3935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$664 final_adder.p_new$688 final_adder.p_new$672 VGND VGND VPWR VPWR
+ final_adder.p_new$792 sky130_fd_sc_hd__and2_1
XU$$503 net1738 net428 net1730 net710 VGND VGND VPWR VPWR t$4662 sky130_fd_sc_hd__a22o_1
XTAP_3946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$514 t$4667 net1250 VGND VGND VPWR VPWR booth_b6_m48 sky130_fd_sc_hd__xor2_1
XFILLER_57_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$675 final_adder.p_new$682 final_adder.g_new$699 final_adder.g_new$683
+ VGND VGND VPWR VPWR final_adder.g_new$803 sky130_fd_sc_hd__a21o_1
XFILLER_179_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$525 net1630 net428 net1621 net710 VGND VGND VPWR VPWR t$4673 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$686 final_adder.p_new$710 final_adder.p_new$694 VGND VGND VPWR VPWR
+ final_adder.p_new$814 sky130_fd_sc_hd__and2_1
XFILLER_29_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$697 final_adder.p_new$704 final_adder.g_new$721 final_adder.g_new$705
+ VGND VGND VPWR VPWR final_adder.g_new$825 sky130_fd_sc_hd__a21o_1
XU$$536 t$4678 net1251 VGND VGND VPWR VPWR booth_b6_m59 sky130_fd_sc_hd__xor2_1
XTAP_3979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$547 net1246 VGND VGND VPWR VPWR notsign$4684 sky130_fd_sc_hd__inv_1
XFILLER_147_1016 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$558 net1126 net414 net1036 net680 VGND VGND VPWR VPWR t$4691 sky130_fd_sc_hd__a22o_1
XU$$569 t$4696 net1241 VGND VGND VPWR VPWR booth_b8_m7 sky130_fd_sc_hd__xor2_1
XFILLER_189_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4423_1832 VGND VGND VPWR VPWR U$$4423_1832/HI net1832 sky130_fd_sc_hd__conb_1
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_51_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_51_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_13_866 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0360_ clknet_leaf_192_clk booth_b32_m43 VGND VGND VPWR VPWR pp_row75_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0291_ clknet_leaf_199_clk booth_b22_m51 VGND VGND VPWR VPWR pp_row73_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2030_ clknet_leaf_76_clk booth_b32_m24 VGND VGND VPWR VPWR pp_row56_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_82_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1220 net1586 net649 net1578 net922 VGND VGND VPWR VPWR t$5028 sky130_fd_sc_hd__a22o_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1231 t$5033 net1013 VGND VGND VPWR VPWR booth_b16_m64 sky130_fd_sc_hd__xor2_1
XFILLER_22_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1242 t$5040 net1664 VGND VGND VPWR VPWR booth_b18_m1 sky130_fd_sc_hd__xor2_1
XU$$1253 net1519 net636 net1513 net909 VGND VGND VPWR VPWR t$5046 sky130_fd_sc_hd__a22o_1
XU$$1264 t$5051 net1662 VGND VGND VPWR VPWR booth_b18_m12 sky130_fd_sc_hd__xor2_1
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_42_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_16
XU$$1275 net1150 net637 net1143 net910 VGND VGND VPWR VPWR t$5057 sky130_fd_sc_hd__a22o_1
XFILLER_176_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1286 t$5062 net1662 VGND VGND VPWR VPWR booth_b18_m23 sky130_fd_sc_hd__xor2_1
XU$$1297 net1048 net636 net1040 net909 VGND VGND VPWR VPWR t$5068 sky130_fd_sc_hd__a22o_1
X_1814_ clknet_leaf_26_clk booth_b38_m11 VGND VGND VPWR VPWR pp_row49_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_91_1 s$3237 s$3239 s$3241 VGND VGND VPWR VPWR c$3762 s$3763 sky130_fd_sc_hd__fa_1
XFILLER_8_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1745_ clknet_leaf_237_clk booth_b16_m31 VGND VGND VPWR VPWR pp_row47_8 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_84_0 c$3188 c$3190 c$3192 VGND VGND VPWR VPWR c$3732 s$3733 sky130_fd_sc_hd__fa_1
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1080 final_adder.$signal$1209 final_adder.g_new$1030 VGND VGND VPWR
+ VPWR net278 sky130_fd_sc_hd__xor2_2
XFILLER_144_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1676_ clknet_leaf_22_clk booth_b42_m2 VGND VGND VPWR VPWR pp_row44_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_116_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0627_ clknet_leaf_177_clk booth_b40_m44 VGND VGND VPWR VPWR pp_row84_11 sky130_fd_sc_hd__dfxtp_1
Xfanout805 net807 VGND VGND VPWR VPWR net805 sky130_fd_sc_hd__buf_4
Xfanout816 net817 VGND VGND VPWR VPWR net816 sky130_fd_sc_hd__buf_4
Xfanout827 net832 VGND VGND VPWR VPWR net827 sky130_fd_sc_hd__buf_4
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_76_7 pp_row76_26 pp_row76_27 pp_row76_28 VGND VGND VPWR VPWR c$830 s$831
+ sky130_fd_sc_hd__fa_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0558_ clknet_leaf_157_clk booth_b64_m17 VGND VGND VPWR VPWR pp_row81_24 sky130_fd_sc_hd__dfxtp_1
XFILLER_58_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout838 net841 VGND VGND VPWR VPWR net838 sky130_fd_sc_hd__clkbuf_8
Xfanout849 net856 VGND VGND VPWR VPWR net849 sky130_fd_sc_hd__buf_4
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_69_6 c$134 c$136 c$138 VGND VGND VPWR VPWR c$702 s$703 sky130_fd_sc_hd__fa_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0489_ clknet_leaf_159_clk booth_b44_m35 VGND VGND VPWR VPWR pp_row79_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_85_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2228_ clknet_leaf_227_clk booth_b10_m52 VGND VGND VPWR VPWR pp_row62_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_209 net1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2159_ clknet_leaf_214_clk booth_b18_m42 VGND VGND VPWR VPWR pp_row60_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_38_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_33_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_107_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_99_0 s$3795 c$4092 s$4095 VGND VGND VPWR VPWR c$4350 s$4351 sky130_fd_sc_hd__fa_1
XFILLER_167_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_100_2 c$1920 c$1922 s$1925 VGND VGND VPWR VPWR c$2642 s$2643 sky130_fd_sc_hd__fa_1
XFILLER_123_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4453_1847 VGND VGND VPWR VPWR U$$4453_1847/HI net1847 sky130_fd_sc_hd__conb_1
XFILLER_27_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_0_64_5 pp_row64_15 pp_row64_16 pp_row64_17 VGND VGND VPWR VPWR c$94 s$95
+ sky130_fd_sc_hd__fa_1
Xdadda_fa_6_114_0 c$3848 c$3850 s$3853 VGND VGND VPWR VPWR c$4124 s$4125 sky130_fd_sc_hd__fa_1
XTAP_3710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$450 final_adder.p_new$456 final_adder.p_new$452 VGND VGND VPWR VPWR
+ final_adder.p_new$578 sky130_fd_sc_hd__and2_1
XFILLER_188_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$300 net1496 net532 net1221 net805 VGND VGND VPWR VPWR t$4559 sky130_fd_sc_hd__a22o_1
XTAP_3732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$461 final_adder.p_new$462 final_adder.g_new$467 final_adder.g_new$463
+ VGND VGND VPWR VPWR final_adder.g_new$589 sky130_fd_sc_hd__a21o_1
XTAP_3743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$311 t$4564 net1279 VGND VGND VPWR VPWR booth_b4_m15 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$472 final_adder.p_new$478 final_adder.p_new$474 VGND VGND VPWR VPWR
+ final_adder.p_new$600 sky130_fd_sc_hd__and2_1
XTAP_3754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$322 net1114 net528 net1105 net801 VGND VGND VPWR VPWR t$4570 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$483 final_adder.p_new$484 final_adder.g_new$489 final_adder.g_new$485
+ VGND VGND VPWR VPWR final_adder.g_new$611 sky130_fd_sc_hd__a21o_1
Xdadda_fa_3_34_3 s$1139 s$1141 s$1143 VGND VGND VPWR VPWR c$2116 s$2117 sky130_fd_sc_hd__fa_1
XTAP_3765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$333 t$4575 net1273 VGND VGND VPWR VPWR booth_b4_m26 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$494 final_adder.p_new$500 final_adder.p_new$496 VGND VGND VPWR VPWR
+ final_adder.p_new$622 sky130_fd_sc_hd__and2_1
XTAP_3776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$344 net1017 net532 net1000 net805 VGND VGND VPWR VPWR t$4581 sky130_fd_sc_hd__a22o_1
XTAP_3787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_27_2 pp_row27_14 c$1062 c$1064 VGND VGND VPWR VPWR c$2058 s$2059 sky130_fd_sc_hd__fa_1
XU$$355 t$4586 net1273 VGND VGND VPWR VPWR booth_b4_m37 sky130_fd_sc_hd__xor2_1
XTAP_3798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$366 net1737 net529 net1729 net802 VGND VGND VPWR VPWR t$4592 sky130_fd_sc_hd__a22o_1
XU$$377 t$4597 net1278 VGND VGND VPWR VPWR booth_b4_m48 sky130_fd_sc_hd__xor2_1
XFILLER_189_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$388 net1633 net533 net1623 net806 VGND VGND VPWR VPWR t$4603 sky130_fd_sc_hd__a22o_1
XU$$399 t$4608 net1275 VGND VGND VPWR VPWR booth_b4_m59 sky130_fd_sc_hd__xor2_1
Xclkbuf_2_3_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_3_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_38_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_24_clk clknet_5_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_73_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1530_ clknet_leaf_17_clk booth_b4_m35 VGND VGND VPWR VPWR pp_row39_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_154_885 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1461_ clknet_leaf_110_clk booth_b62_m42 VGND VGND VPWR VPWR pp_row104_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_79_5 s$881 s$883 s$885 VGND VGND VPWR VPWR c$1684 s$1685 sky130_fd_sc_hd__fa_2
X_0412_ clknet_leaf_192_clk notsign$4894 VGND VGND VPWR VPWR pp_row77_0 sky130_fd_sc_hd__dfxtp_1
X_1392_ clknet_leaf_54_clk booth_b0_m33 VGND VGND VPWR VPWR pp_row33_0 sky130_fd_sc_hd__dfxtp_1
Xdadda_ha_2_30_4 pp_row30_12 pp_row30_13 VGND VGND VPWR VPWR c$1098 s$1099 sky130_fd_sc_hd__ha_1
XU$$1924_1769 VGND VGND VPWR VPWR U$$1924_1769/HI net1769 sky130_fd_sc_hd__conb_1
XFILLER_45_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0343_ clknet_leaf_203_clk booth_b60_m14 VGND VGND VPWR VPWR pp_row74_26 sky130_fd_sc_hd__dfxtp_1
XFILLER_94_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0274_ clknet_leaf_217_clk booth_b54_m18 VGND VGND VPWR VPWR pp_row72_24 sky130_fd_sc_hd__dfxtp_1
Xdadda_ha_7_0_0 pp_row0_0 pp_row0_1 VGND VGND VPWR VPWR c$4152 s$4153 sky130_fd_sc_hd__ha_1
X_2013_ clknet_leaf_83_clk booth_b2_m54 VGND VGND VPWR VPWR pp_row56_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_36_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_991 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_15_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_16
XU$$1050 t$4941 net1187 VGND VGND VPWR VPWR booth_b14_m42 sky130_fd_sc_hd__xor2_1
XU$$1061 net1695 net390 net1687 net656 VGND VGND VPWR VPWR t$4947 sky130_fd_sc_hd__a22o_1
XU$$1072 t$4952 net1191 VGND VGND VPWR VPWR booth_b14_m53 sky130_fd_sc_hd__xor2_1
XFILLER_149_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1083 net1586 net390 net1578 net656 VGND VGND VPWR VPWR t$4958 sky130_fd_sc_hd__a22o_1
XFILLER_176_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1094 t$4963 net1189 VGND VGND VPWR VPWR booth_b14_m64 sky130_fd_sc_hd__xor2_1
XFILLER_177_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_1_82_7 pp_row82_21 pp_row82_22 VGND VGND VPWR VPWR c$936 s$937 sky130_fd_sc_hd__ha_1
XFILLER_176_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_109_1 s$3345 s$3347 s$3349 VGND VGND VPWR VPWR c$3834 s$3835 sky130_fd_sc_hd__fa_1
X_1728_ clknet_leaf_164_clk booth_b64_m59 VGND VGND VPWR VPWR pp_row123_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_81_5 pp_row81_15 pp_row81_16 pp_row81_17 VGND VGND VPWR VPWR c$916 s$917
+ sky130_fd_sc_hd__fa_1
X_1659_ clknet_leaf_21_clk booth_b12_m32 VGND VGND VPWR VPWR pp_row44_6 sky130_fd_sc_hd__dfxtp_1
Xfanout602 net604 VGND VGND VPWR VPWR net602 sky130_fd_sc_hd__buf_4
Xfanout613 net615 VGND VGND VPWR VPWR net613 sky130_fd_sc_hd__buf_4
Xfanout624 net625 VGND VGND VPWR VPWR net624 sky130_fd_sc_hd__clkbuf_4
Xfanout635 net636 VGND VGND VPWR VPWR net635 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_74_4 pp_row74_20 pp_row74_21 pp_row74_22 VGND VGND VPWR VPWR c$788 s$789
+ sky130_fd_sc_hd__fa_1
XFILLER_98_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout646 net647 VGND VGND VPWR VPWR net646 sky130_fd_sc_hd__buf_6
Xfanout657 net658 VGND VGND VPWR VPWR net657 sky130_fd_sc_hd__buf_6
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_67_3 pp_row67_27 pp_row67_28 pp_row67_29 VGND VGND VPWR VPWR c$660 s$661
+ sky130_fd_sc_hd__fa_1
Xfanout668 net674 VGND VGND VPWR VPWR net668 sky130_fd_sc_hd__buf_4
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout679 net680 VGND VGND VPWR VPWR net679 sky130_fd_sc_hd__buf_4
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_44_2 s$2193 s$2195 s$2197 VGND VGND VPWR VPWR c$2958 s$2959 sky130_fd_sc_hd__fa_1
XFILLER_86_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_37_1 c$2130 c$2132 s$2135 VGND VGND VPWR VPWR c$2914 s$2915 sky130_fd_sc_hd__fa_1
XTAP_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_14_0 s$3455 c$3922 s$3925 VGND VGND VPWR VPWR c$4180 s$4181 sky130_fd_sc_hd__fa_1
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_0_62_2 pp_row62_6 pp_row62_7 pp_row62_8 VGND VGND VPWR VPWR c$64 s$65 sky130_fd_sc_hd__fa_1
XFILLER_49_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3903 t$6399 net1294 VGND VGND VPWR VPWR booth_b56_m30 sky130_fd_sc_hd__xor2_1
XFILLER_65_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3914 net979 net465 net970 net738 VGND VGND VPWR VPWR t$6405 sky130_fd_sc_hd__a22o_1
XTAP_4263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3925 t$6410 net1297 VGND VGND VPWR VPWR booth_b56_m41 sky130_fd_sc_hd__xor2_1
XTAP_4274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3936 net1709 net466 net1701 net739 VGND VGND VPWR VPWR t$6416 sky130_fd_sc_hd__a22o_1
XTAP_3540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_32_0 pp_row32_17 pp_row32_18 c$1100 VGND VGND VPWR VPWR c$2094 s$2095
+ sky130_fd_sc_hd__fa_2
XU$$3947 t$6421 net1293 VGND VGND VPWR VPWR booth_b56_m52 sky130_fd_sc_hd__xor2_1
XTAP_4296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$280 final_adder.p_new$282 final_adder.p_new$280 VGND VGND VPWR VPWR
+ final_adder.p_new$408 sky130_fd_sc_hd__and2_1
XFILLER_45_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3958 net1601 net465 net1591 net738 VGND VGND VPWR VPWR t$6427 sky130_fd_sc_hd__a22o_1
XTAP_3562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$130 net1543 net444 net1535 net686 VGND VGND VPWR VPWR t$4472 sky130_fd_sc_hd__a22o_1
XU$$3969 t$6432 net1293 VGND VGND VPWR VPWR booth_b56_m63 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$291 final_adder.p_new$290 final_adder.g_new$293 final_adder.g_new$291
+ VGND VGND VPWR VPWR final_adder.g_new$419 sky130_fd_sc_hd__a21o_1
XTAP_3573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$141 notblock$4475\[2\] net23 net1571 t$4476 notblock$4475\[0\] VGND VGND VPWR
+ VPWR sel_0$4477 sky130_fd_sc_hd__a32o_4
XU$$152 t$4483 net1390 VGND VGND VPWR VPWR booth_b2_m4 sky130_fd_sc_hd__xor2_1
XTAP_3584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$163 net1499 net624 net1224 net897 VGND VGND VPWR VPWR t$4489 sky130_fd_sc_hd__a22o_1
XFILLER_72_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$174 t$4494 net1386 VGND VGND VPWR VPWR booth_b2_m15 sky130_fd_sc_hd__xor2_1
XU$$185 net1117 net623 net1108 net896 VGND VGND VPWR VPWR t$4500 sky130_fd_sc_hd__a22o_1
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$196 t$4505 net1385 VGND VGND VPWR VPWR booth_b2_m26 sky130_fd_sc_hd__xor2_1
XFILLER_60_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0961_ clknet_leaf_114_clk notsign$5664 VGND VGND VPWR VPWR pp_row99_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_174_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0892_ clknet_leaf_100_clk booth_b50_m45 VGND VGND VPWR VPWR pp_row95_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_185_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_91_4 c$1018 c$1020 c$1022 VGND VGND VPWR VPWR c$1826 s$1827 sky130_fd_sc_hd__fa_1
XFILLER_142_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_84_3 c$946 c$948 c$950 VGND VGND VPWR VPWR c$1740 s$1741 sky130_fd_sc_hd__fa_1
X_1513_ clknet_leaf_44_clk booth_b18_m20 VGND VGND VPWR VPWR pp_row38_9 sky130_fd_sc_hd__dfxtp_1
X_2493_ clknet_leaf_90_clk booth_b26_m43 VGND VGND VPWR VPWR pp_row69_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_99_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_77_2 c$826 c$828 c$830 VGND VGND VPWR VPWR c$1654 s$1655 sky130_fd_sc_hd__fa_1
XFILLER_102_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_4_clk clknet_5_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_16
X_1444_ clknet_leaf_54_clk booth_b14_m21 VGND VGND VPWR VPWR pp_row35_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_96_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_54_1 s$3015 s$3017 s$3019 VGND VGND VPWR VPWR c$3614 s$3615 sky130_fd_sc_hd__fa_1
X_1375_ clknet_leaf_7_clk booth_b6_m26 VGND VGND VPWR VPWR pp_row32_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_67_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_47_0 c$2966 c$2968 c$2970 VGND VGND VPWR VPWR c$3584 s$3585 sky130_fd_sc_hd__fa_1
X_0326_ clknet_leaf_201_clk booth_b28_m46 VGND VGND VPWR VPWR pp_row74_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_83_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0257_ clknet_leaf_209_clk booth_b22_m50 VGND VGND VPWR VPWR pp_row72_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_55_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0188_ clknet_leaf_148_clk booth_b20_m50 VGND VGND VPWR VPWR pp_row70_8 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_100_1 pp_row100_3 pp_row100_4 pp_row100_5 VGND VGND VPWR VPWR c$1926 s$1927
+ sky130_fd_sc_hd__fa_1
XFILLER_169_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3020_1787 VGND VGND VPWR VPWR U$$3020_1787/HI net1787 sky130_fd_sc_hd__conb_1
Xdadda_fa_5_121_0 pp_row121_3 pp_row121_4 pp_row121_5 VGND VGND VPWR VPWR c$3880 s$3881
+ sky130_fd_sc_hd__fa_2
Xclkbuf_5_18__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_5_18__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_176_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout410 net412 VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__buf_4
Xfanout1408 net1411 VGND VGND VPWR VPWR net1408 sky130_fd_sc_hd__clkbuf_8
Xfanout1419 net3 VGND VGND VPWR VPWR net1419 sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_1_72_1 pp_row72_14 pp_row72_15 pp_row72_16 VGND VGND VPWR VPWR c$746 s$747
+ sky130_fd_sc_hd__fa_1
Xfanout421 sel_0$6577 VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__buf_6
Xfanout432 net433 VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__buf_6
XFILLER_48_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout443 net450 VGND VGND VPWR VPWR net443 sky130_fd_sc_hd__buf_2
XFILLER_115_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout454 net459 VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__buf_4
XFILLER_63_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_65_0 pp_row65_18 pp_row65_19 pp_row65_20 VGND VGND VPWR VPWR c$618 s$619
+ sky130_fd_sc_hd__fa_2
Xfanout465 net467 VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__clkbuf_8
XFILLER_24_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout476 net479 VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__buf_6
XFILLER_86_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout487 sel_0$6157 VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__clkbuf_8
Xfanout498 net499 VGND VGND VPWR VPWR net498 sky130_fd_sc_hd__buf_4
XFILLER_58_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1029 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2509 t$5687 net1406 VGND VGND VPWR VPWR booth_b36_m18 sky130_fd_sc_hd__xor2_1
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1808 t$5329 net1460 VGND VGND VPWR VPWR booth_b26_m10 sky130_fd_sc_hd__xor2_1
XU$$1819 net1165 net593 net1155 net866 VGND VGND VPWR VPWR t$5335 sky130_fd_sc_hd__a22o_1
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_936 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_94_2 c$1852 s$1855 s$1857 VGND VGND VPWR VPWR c$2594 s$2595 sky130_fd_sc_hd__fa_1
XFILLER_182_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_87_1 c$1762 c$1764 c$1766 VGND VGND VPWR VPWR c$2536 s$2537 sky130_fd_sc_hd__fa_1
XFILLER_123_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_6_64_0 c$3648 c$3650 s$3653 VGND VGND VPWR VPWR c$4024 s$4025 sky130_fd_sc_hd__fa_1
XFILLER_89_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4401 t$6654 net1821 VGND VGND VPWR VPWR booth_b64_m5 sky130_fd_sc_hd__xor2_1
XU$$4412 net1222 sel_0$6647 net1214 net694 VGND VGND VPWR VPWR t$6660 sky130_fd_sc_hd__a22o_1
XFILLER_49_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1160_ clknet_leaf_182_clk net132 VGND VGND VPWR VPWR pp_row102_15 sky130_fd_sc_hd__dfxtp_4
XU$$4423 t$6665 net1832 VGND VGND VPWR VPWR booth_b64_m16 sky130_fd_sc_hd__xor2_1
XU$$4434 net1112 sel_0$6647 net1103 net695 VGND VGND VPWR VPWR t$6671 sky130_fd_sc_hd__a22o_1
XU$$3700 net50 VGND VGND VPWR VPWR notblock$6295\[1\] sky130_fd_sc_hd__inv_1
XU$$4445 t$6676 net1843 VGND VGND VPWR VPWR booth_b64_m27 sky130_fd_sc_hd__xor2_1
XU$$4456 net1005 sel_0$6647 net997 net697 VGND VGND VPWR VPWR t$6682 sky130_fd_sc_hd__a22o_1
XFILLER_65_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3711 net1037 net472 net938 net745 VGND VGND VPWR VPWR t$6302 sky130_fd_sc_hd__a22o_1
XTAP_4060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4467 t$6687 net1854 VGND VGND VPWR VPWR booth_b64_m38 sky130_fd_sc_hd__xor2_1
XU$$3722 t$6307 net1309 VGND VGND VPWR VPWR booth_b54_m8 sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_116_1 pp_row116_5 pp_row116_6 pp_row116_7 VGND VGND VPWR VPWR c$3388 s$3389
+ sky130_fd_sc_hd__fa_1
XTAP_4071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3733 net1200 net475 net1181 net748 VGND VGND VPWR VPWR t$6313 sky130_fd_sc_hd__a22o_1
XU$$4478 net1735 sel_0$6647 net1727 net696 VGND VGND VPWR VPWR t$6693 sky130_fd_sc_hd__a22o_1
X_1091_ clknet_leaf_59_clk net1313 VGND VGND VPWR VPWR pp_row12_7 sky130_fd_sc_hd__dfxtp_1
XTAP_4082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3744 t$6318 net1300 VGND VGND VPWR VPWR booth_b54_m19 sky130_fd_sc_hd__xor2_1
XTAP_4093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4489 t$6698 net1865 VGND VGND VPWR VPWR booth_b64_m49 sky130_fd_sc_hd__xor2_1
XU$$3755 net1085 net470 net1076 net743 VGND VGND VPWR VPWR t$6324 sky130_fd_sc_hd__a22o_1
XFILLER_92_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_109_0 c$1972 c$2702 c$2704 VGND VGND VPWR VPWR c$3344 s$3345 sky130_fd_sc_hd__fa_1
XU$$3766 t$6329 net1303 VGND VGND VPWR VPWR booth_b54_m30 sky130_fd_sc_hd__xor2_1
XTAP_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3777 net979 net473 net970 net746 VGND VGND VPWR VPWR t$6335 sky130_fd_sc_hd__a22o_1
XU$$3788 t$6340 net1305 VGND VGND VPWR VPWR booth_b54_m41 sky130_fd_sc_hd__xor2_1
XFILLER_18_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3799 net1709 net474 net1701 net747 VGND VGND VPWR VPWR t$6346 sky130_fd_sc_hd__a22o_1
XTAP_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_370 net1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_381 net1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_392 net1530 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1993_ clknet_leaf_67_clk booth_b24_m31 VGND VGND VPWR VPWR pp_row55_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_20_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0944_ clknet_leaf_180_clk booth_b64_m63 VGND VGND VPWR VPWR pp_row127_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_9_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0875_ clknet_leaf_93_clk booth_b58_m36 VGND VGND VPWR VPWR pp_row94_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_161_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_811 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_82_0 pp_row82_23 pp_row82_24 pp_row82_25 VGND VGND VPWR VPWR c$1710 s$1711
+ sky130_fd_sc_hd__fa_1
XFILLER_126_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2476_ clknet_leaf_99_clk booth_b60_m8 VGND VGND VPWR VPWR pp_row68_29 sky130_fd_sc_hd__dfxtp_1
XFILLER_134_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1427_ clknet_leaf_64_clk booth_b24_m10 VGND VGND VPWR VPWR pp_row34_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_87_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_975 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1358_ clknet_leaf_10_clk booth_b10_m21 VGND VGND VPWR VPWR pp_row31_5 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_51_6 pp_row51_18 pp_row51_19 pp_row51_20 VGND VGND VPWR VPWR c$378 s$379
+ sky130_fd_sc_hd__fa_1
XFILLER_83_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0309_ clknet_leaf_209_clk booth_b56_m17 VGND VGND VPWR VPWR pp_row73_24 sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1289_ clknet_leaf_2_clk booth_b16_m11 VGND VGND VPWR VPWR pp_row27_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_71_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_3_0 pp_row3_2 c$3900 s$3903 VGND VGND VPWR VPWR c$4158 s$4159 sky130_fd_sc_hd__fa_1
XFILLER_36_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_81_0 s$3723 c$4056 s$4059 VGND VGND VPWR VPWR c$4314 s$4315 sky130_fd_sc_hd__fa_2
Xdadda_fa_4_97_0 s$1901 c$2606 c$2608 VGND VGND VPWR VPWR c$3272 s$3273 sky130_fd_sc_hd__fa_1
XFILLER_4_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1205 net1209 VGND VGND VPWR VPWR net1205 sky130_fd_sc_hd__buf_6
Xfanout1216 net1218 VGND VGND VPWR VPWR net1216 sky130_fd_sc_hd__clkbuf_8
Xfanout1227 net1229 VGND VGND VPWR VPWR net1227 sky130_fd_sc_hd__buf_4
Xfanout1238 net64 VGND VGND VPWR VPWR net1238 sky130_fd_sc_hd__buf_4
Xfanout1249 net1252 VGND VGND VPWR VPWR net1249 sky130_fd_sc_hd__clkbuf_4
XFILLER_74_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3007 net1548 net525 net1540 net798 VGND VGND VPWR VPWR t$5941 sky130_fd_sc_hd__a22o_1
XU$$3018 notblock$5945\[2\] net39 net1369 t$5946 notblock$5945\[0\] VGND VGND VPWR
+ VPWR sel_0$5947 sky130_fd_sc_hd__a32o_1
XFILLER_189_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3029 t$5953 net1357 VGND VGND VPWR VPWR booth_b44_m4 sky130_fd_sc_hd__xor2_1
XFILLER_75_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2306 net1631 net574 net1622 net847 VGND VGND VPWR VPWR t$5583 sky130_fd_sc_hd__a22o_1
XFILLER_74_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2317 t$5588 net1437 VGND VGND VPWR VPWR booth_b32_m59 sky130_fd_sc_hd__xor2_1
XU$$2328 net1437 VGND VGND VPWR VPWR notsign$5594 sky130_fd_sc_hd__inv_1
XU$$2339 net1126 net563 net1036 net836 VGND VGND VPWR VPWR t$5601 sky130_fd_sc_hd__a22o_1
XU$$1605 net1719 net618 net1710 net891 VGND VGND VPWR VPWR t$5225 sky130_fd_sc_hd__a22o_1
XFILLER_131_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1616 t$5230 net1483 VGND VGND VPWR VPWR booth_b22_m51 sky130_fd_sc_hd__xor2_1
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1627 net1605 net617 net1597 net890 VGND VGND VPWR VPWR t$5236 sky130_fd_sc_hd__a22o_1
XFILLER_188_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1638 t$5241 net1481 VGND VGND VPWR VPWR booth_b22_m62 sky130_fd_sc_hd__xor2_1
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1649 net17 net1482 VGND VGND VPWR VPWR sel_1$5248 sky130_fd_sc_hd__xor2_4
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1080 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0660_ clknet_leaf_175_clk booth_b52_m33 VGND VGND VPWR VPWR pp_row85_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_115_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0591_ clknet_leaf_186_clk booth_b24_m59 VGND VGND VPWR VPWR pp_row83_3 sky130_fd_sc_hd__dfxtp_1
X_2330_ clknet_leaf_99_clk booth_b60_m4 VGND VGND VPWR VPWR pp_row64_30 sky130_fd_sc_hd__dfxtp_1
XFILLER_3_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2261_ clknet_leaf_199_clk booth_b2_m61 VGND VGND VPWR VPWR pp_row63_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_112_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_61_5 s$557 s$559 s$561 VGND VGND VPWR VPWR c$1468 s$1469 sky130_fd_sc_hd__fa_1
Xfanout1750 net1751 VGND VGND VPWR VPWR net1750 sky130_fd_sc_hd__buf_4
XFILLER_66_912 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1212_ clknet_leaf_49_clk booth_b22_m0 VGND VGND VPWR VPWR pp_row22_11 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_54_4 s$425 s$427 s$429 VGND VGND VPWR VPWR c$1382 s$1383 sky130_fd_sc_hd__fa_1
X_2192_ clknet_leaf_223_clk booth_b10_m51 VGND VGND VPWR VPWR pp_row61_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_133_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4220 net1651 net439 net1643 net721 VGND VGND VPWR VPWR t$6561 sky130_fd_sc_hd__a22o_1
XU$$4231 t$6566 net1265 VGND VGND VPWR VPWR booth_b60_m57 sky130_fd_sc_hd__xor2_1
XFILLER_65_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4242 net1537 net435 net1529 net717 VGND VGND VPWR VPWR t$6572 sky130_fd_sc_hd__a22o_1
XU$$4253 net1808 net421 net1233 net703 VGND VGND VPWR VPWR t$6579 sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_47_3 c$296 c$298 c$300 VGND VGND VPWR VPWR c$1296 s$1297 sky130_fd_sc_hd__fa_1
X_1143_ clknet_leaf_11_clk booth_b14_m3 VGND VGND VPWR VPWR pp_row17_7 sky130_fd_sc_hd__dfxtp_1
XU$$4264 t$6584 net1259 VGND VGND VPWR VPWR booth_b62_m5 sky130_fd_sc_hd__xor2_1
XU$$3530 t$6208 net1335 VGND VGND VPWR VPWR booth_b50_m49 sky130_fd_sc_hd__xor2_1
XU$$4275 net1222 net418 net1214 net700 VGND VGND VPWR VPWR t$6590 sky130_fd_sc_hd__a22o_1
XU$$3541 net1627 net490 net1618 net763 VGND VGND VPWR VPWR t$6214 sky130_fd_sc_hd__a22o_1
XU$$4286 t$6595 net1258 VGND VGND VPWR VPWR booth_b62_m16 sky130_fd_sc_hd__xor2_1
XU$$4297 net1112 net419 net1103 net701 VGND VGND VPWR VPWR t$6601 sky130_fd_sc_hd__a22o_1
XU$$3552 t$6219 net1334 VGND VGND VPWR VPWR booth_b50_m60 sky130_fd_sc_hd__xor2_1
XU$$3563 net48 VGND VGND VPWR VPWR notblock$6225\[1\] sky130_fd_sc_hd__inv_1
XFILLER_93_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1074_ clknet_leaf_53_clk net1415 VGND VGND VPWR VPWR pp_row10_6 sky130_fd_sc_hd__dfxtp_1
XU$$3574 net1037 net480 net938 net753 VGND VGND VPWR VPWR t$6232 sky130_fd_sc_hd__a22o_1
XU$$3585 t$6237 net1319 VGND VGND VPWR VPWR booth_b52_m8 sky130_fd_sc_hd__xor2_1
XU$$2840 net1705 net537 net1697 net810 VGND VGND VPWR VPWR t$5856 sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_17_1 s$2793 s$2795 s$2797 VGND VGND VPWR VPWR c$3466 s$3467 sky130_fd_sc_hd__fa_1
XU$$3596 net1200 net480 net1181 net753 VGND VGND VPWR VPWR t$6243 sky130_fd_sc_hd__a22o_1
XU$$2851 t$5861 net1382 VGND VGND VPWR VPWR booth_b40_m52 sky130_fd_sc_hd__xor2_1
XU$$2862 net1602 net540 net1592 net813 VGND VGND VPWR VPWR t$5867 sky130_fd_sc_hd__a22o_1
XU$$2873 t$5872 net1383 VGND VGND VPWR VPWR booth_b40_m63 sky130_fd_sc_hd__xor2_1
XU$$2884 t$5879 net1367 VGND VGND VPWR VPWR booth_b42_m0 sky130_fd_sc_hd__xor2_1
XFILLER_33_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2895 net1562 net519 net1520 net792 VGND VGND VPWR VPWR t$5885 sky130_fd_sc_hd__a22o_1
XFILLER_21_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1976_ clknet_leaf_72_clk booth_b52_m2 VGND VGND VPWR VPWR pp_row54_26 sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0927_ clknet_leaf_112_clk booth_b42_m55 VGND VGND VPWR VPWR pp_row97_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_147_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_939 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0858_ clknet_leaf_140_clk booth_b64_m29 VGND VGND VPWR VPWR pp_row93_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_162_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_4_120_1 pp_row120_3 pp_row120_4 VGND VGND VPWR VPWR c$3410 s$3411 sky130_fd_sc_hd__ha_1
XFILLER_115_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0789_ clknet_leaf_138_clk booth_b62_m28 VGND VGND VPWR VPWR pp_row90_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_143_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_1_43_4 pp_row43_12 pp_row43_13 VGND VGND VPWR VPWR c$262 s$263 sky130_fd_sc_hd__ha_1
Xdadda_ha_3_116_0_1918 VGND VGND VPWR VPWR net1918 dadda_ha_3_116_0_1918/LO sky130_fd_sc_hd__conb_1
XFILLER_25_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2459_ clknet_leaf_148_clk booth_b28_m40 VGND VGND VPWR VPWR pp_row68_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_152_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$813 final_adder.p_new$828 final_adder.g_new$861 final_adder.g_new$829
+ VGND VGND VPWR VPWR final_adder.g_new$941 sky130_fd_sc_hd__a21o_2
XFILLER_56_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_ha_4_13_2 pp_row13_6 pp_row13_7 VGND VGND VPWR VPWR c$2772 s$2773 sky130_fd_sc_hd__ha_1
XFILLER_56_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$857 final_adder.p_new$888 final_adder.g_new$953 final_adder.g_new$889
+ VGND VGND VPWR VPWR final_adder.g_new$985 sky130_fd_sc_hd__a21o_2
XFILLER_57_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$707 net1513 net406 net1505 net672 VGND VGND VPWR VPWR t$4767 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$879 final_adder.p_new$910 final_adder.g_new$863 final_adder.g_new$911
+ VGND VGND VPWR VPWR final_adder.g_new$1007 sky130_fd_sc_hd__a21o_1
XU$$718 t$4772 net1415 VGND VGND VPWR VPWR booth_b10_m13 sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_42_2 pp_row42_6 pp_row42_7 pp_row42_8 VGND VGND VPWR VPWR c$248 s$249
+ sky130_fd_sc_hd__fa_1
XU$$729 net1138 net401 net1130 net667 VGND VGND VPWR VPWR t$4778 sky130_fd_sc_hd__a22o_1
XFILLER_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_12_0 pp_row12_0 pp_row12_1 pp_row12_2 VGND VGND VPWR VPWR c$2762 s$2763
+ sky130_fd_sc_hd__fa_1
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4417_1829 VGND VGND VPWR VPWR U$$4417_1829/HI net1829 sky130_fd_sc_hd__conb_1
XFILLER_193_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1002 net1004 VGND VGND VPWR VPWR net1002 sky130_fd_sc_hd__buf_6
XFILLER_117_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1013 net1014 VGND VGND VPWR VPWR net1013 sky130_fd_sc_hd__buf_4
Xdadda_fa_3_64_3 s$1499 s$1501 s$1503 VGND VGND VPWR VPWR c$2356 s$2357 sky130_fd_sc_hd__fa_1
Xfanout1024 net1030 VGND VGND VPWR VPWR net1024 sky130_fd_sc_hd__buf_6
XFILLER_0_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1035 net1038 VGND VGND VPWR VPWR net1035 sky130_fd_sc_hd__clkbuf_4
Xfanout1046 net86 VGND VGND VPWR VPWR net1046 sky130_fd_sc_hd__buf_6
Xfanout1057 net1058 VGND VGND VPWR VPWR net1057 sky130_fd_sc_hd__buf_4
Xdadda_fa_3_57_2 c$1408 s$1411 s$1413 VGND VGND VPWR VPWR c$2298 s$2299 sky130_fd_sc_hd__fa_1
Xfanout1068 net1070 VGND VGND VPWR VPWR net1068 sky130_fd_sc_hd__clkbuf_8
Xfanout1079 net82 VGND VGND VPWR VPWR net1079 sky130_fd_sc_hd__buf_4
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_27_0 c$3500 c$3502 s$3505 VGND VGND VPWR VPWR c$3950 s$3951 sky130_fd_sc_hd__fa_2
Xclkbuf_leaf_210_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_210_clk
+ sky130_fd_sc_hd__clkbuf_16
XU$$2103 net1118 net580 net1109 net853 VGND VGND VPWR VPWR t$5480 sky130_fd_sc_hd__a22o_1
XFILLER_35_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2114 t$5485 net1442 VGND VGND VPWR VPWR booth_b30_m26 sky130_fd_sc_hd__xor2_1
XU$$2125 net1016 net576 net999 net849 VGND VGND VPWR VPWR t$5491 sky130_fd_sc_hd__a22o_1
XFILLER_16_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2136 t$5496 net1443 VGND VGND VPWR VPWR booth_b30_m37 sky130_fd_sc_hd__xor2_1
XFILLER_74_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2147 net1737 net578 net1729 net851 VGND VGND VPWR VPWR t$5502 sky130_fd_sc_hd__a22o_1
XU$$1402 net1206 net629 net1198 net902 VGND VGND VPWR VPWR t$5122 sky130_fd_sc_hd__a22o_1
XFILLER_34_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2158 t$5507 net1446 VGND VGND VPWR VPWR booth_b30_m48 sky130_fd_sc_hd__xor2_1
XU$$1413 t$5127 net1487 VGND VGND VPWR VPWR booth_b20_m18 sky130_fd_sc_hd__xor2_1
XU$$1424 net1089 net628 net1081 net901 VGND VGND VPWR VPWR t$5133 sky130_fd_sc_hd__a22o_1
XU$$2169 net1631 net578 net1622 net851 VGND VGND VPWR VPWR t$5513 sky130_fd_sc_hd__a22o_1
XU$$1435 t$5138 net1486 VGND VGND VPWR VPWR booth_b20_m29 sky130_fd_sc_hd__xor2_1
XU$$1446 net987 net630 net977 net903 VGND VGND VPWR VPWR t$5144 sky130_fd_sc_hd__a22o_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1457 t$5149 net1490 VGND VGND VPWR VPWR booth_b20_m40 sky130_fd_sc_hd__xor2_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1468 net1715 net630 net1706 net903 VGND VGND VPWR VPWR t$5155 sky130_fd_sc_hd__a22o_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1479 t$5160 net1492 VGND VGND VPWR VPWR booth_b20_m51 sky130_fd_sc_hd__xor2_1
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1830_ clknet_leaf_34_clk booth_b14_m36 VGND VGND VPWR VPWR pp_row50_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_191_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1761_ clknet_leaf_187_clk booth_b62_m44 VGND VGND VPWR VPWR pp_row106_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_184_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0712_ clknet_leaf_165_clk booth_b54_m33 VGND VGND VPWR VPWR pp_row87_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_116_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1692_ clknet_leaf_19_clk booth_b22_m23 VGND VGND VPWR VPWR pp_row45_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_144_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0643_ clknet_leaf_180_clk booth_b22_m63 VGND VGND VPWR VPWR pp_row85_1 sky130_fd_sc_hd__dfxtp_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0574_ clknet_leaf_190_clk booth_b44_m38 VGND VGND VPWR VPWR pp_row82_14 sky130_fd_sc_hd__dfxtp_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2313_ clknet_leaf_30_clk booth_b30_m34 VGND VGND VPWR VPWR pp_row64_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_97_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$109 c$4368 s$4371 VGND VGND VPWR VPWR final_adder.$signal$220 final_adder.$signal$1199
+ sky130_fd_sc_hd__ha_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2244_ clknet_leaf_30_clk booth_b40_m22 VGND VGND VPWR VPWR pp_row62_20 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_52_1 c$370 c$372 c$374 VGND VGND VPWR VPWR c$1352 s$1353 sky130_fd_sc_hd__fa_1
XFILLER_38_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1580 net1581 VGND VGND VPWR VPWR net1580 sky130_fd_sc_hd__clkbuf_4
Xfanout1591 net1592 VGND VGND VPWR VPWR net1591 sky130_fd_sc_hd__buf_4
X_2175_ clknet_leaf_224_clk booth_b44_m16 VGND VGND VPWR VPWR pp_row60_22 sky130_fd_sc_hd__dfxtp_1
XFILLER_93_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4050 t$6474 net1283 VGND VGND VPWR VPWR booth_b58_m35 sky130_fd_sc_hd__xor2_1
XFILLER_122_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4061 net929 net457 net1750 net730 VGND VGND VPWR VPWR t$6480 sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_45_0 pp_row45_17 pp_row45_18 pp_row45_19 VGND VGND VPWR VPWR c$1266 s$1267
+ sky130_fd_sc_hd__fa_1
XFILLER_93_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4072 t$6485 net1289 VGND VGND VPWR VPWR booth_b58_m46 sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_201_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_201_clk
+ sky130_fd_sc_hd__clkbuf_16
X_1126_ clknet_leaf_12_clk booth_b6_m10 VGND VGND VPWR VPWR pp_row16_3 sky130_fd_sc_hd__dfxtp_1
XU$$4083 net1651 net456 net1643 net729 VGND VGND VPWR VPWR t$6491 sky130_fd_sc_hd__a22o_1
XU$$4094 t$6496 net1288 VGND VGND VPWR VPWR booth_b58_m57 sky130_fd_sc_hd__xor2_1
XU$$3360 net1002 net494 net995 net767 VGND VGND VPWR VPWR t$6122 sky130_fd_sc_hd__a22o_1
XFILLER_81_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3371 t$6127 net1341 VGND VGND VPWR VPWR booth_b48_m38 sky130_fd_sc_hd__xor2_1
XU$$3382 net1734 net498 net1726 net771 VGND VGND VPWR VPWR t$6133 sky130_fd_sc_hd__a22o_1
XU$$3393 t$6138 net1344 VGND VGND VPWR VPWR booth_b48_m49 sky130_fd_sc_hd__xor2_1
X_1057_ clknet_leaf_58_clk net1240 VGND VGND VPWR VPWR pp_row8_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_181_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2670 t$5769 net1400 VGND VGND VPWR VPWR booth_b38_m30 sky130_fd_sc_hd__xor2_1
XFILLER_15_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2681 net974 net543 net965 net816 VGND VGND VPWR VPWR t$5775 sky130_fd_sc_hd__a22o_1
XFILLER_181_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2692 t$5780 net1396 VGND VGND VPWR VPWR booth_b38_m41 sky130_fd_sc_hd__xor2_1
XFILLER_22_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1980 net1058 net588 net1050 net861 VGND VGND VPWR VPWR t$5417 sky130_fd_sc_hd__a22o_1
XFILLER_33_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1991 t$5422 net1452 VGND VGND VPWR VPWR booth_b28_m33 sky130_fd_sc_hd__xor2_1
XFILLER_166_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_889 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1959_ clknet_leaf_63_clk booth_b22_m32 VGND VGND VPWR VPWR pp_row54_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_175_861 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_74_2 s$2433 s$2435 s$2437 VGND VGND VPWR VPWR c$3138 s$3139 sky130_fd_sc_hd__fa_1
XFILLER_163_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_67_1 c$2370 c$2372 s$2375 VGND VGND VPWR VPWR c$3094 s$3095 sky130_fd_sc_hd__fa_1
XFILLER_131_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput105 b[46] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__buf_6
Xinput116 b[56] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__buf_2
Xdadda_fa_7_44_0 s$3575 c$3982 s$3985 VGND VGND VPWR VPWR c$4240 s$4241 sky130_fd_sc_hd__fa_2
XFILLER_48_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput127 b[8] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__buf_6
Xinput138 c[108] VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_1
Xdadda_ha_1_34_0 pp_row34_0 pp_row34_1 VGND VGND VPWR VPWR c$204 s$205 sky130_fd_sc_hd__ha_1
Xinput149 c[118] VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_1
Xfinal_adder.U$$610 final_adder.p_new$622 final_adder.p_new$614 VGND VGND VPWR VPWR
+ final_adder.p_new$738 sky130_fd_sc_hd__and2_1
XFILLER_69_591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$621 final_adder.p_new$624 final_adder.g_new$633 final_adder.g_new$625
+ VGND VGND VPWR VPWR final_adder.g_new$749 sky130_fd_sc_hd__a21o_4
XTAP_3903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$632 final_adder.p_new$656 final_adder.p_new$640 VGND VGND VPWR VPWR
+ final_adder.p_new$760 sky130_fd_sc_hd__and2_1
XFILLER_5_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$643 final_adder.p_new$650 final_adder.g_new$667 final_adder.g_new$651
+ VGND VGND VPWR VPWR final_adder.g_new$771 sky130_fd_sc_hd__a21o_1
XTAP_3925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$654 final_adder.p_new$678 final_adder.p_new$662 VGND VGND VPWR VPWR
+ final_adder.p_new$782 sky130_fd_sc_hd__and2_1
XTAP_3936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$665 final_adder.p_new$672 final_adder.g_new$689 final_adder.g_new$673
+ VGND VGND VPWR VPWR final_adder.g_new$793 sky130_fd_sc_hd__a21o_1
XFILLER_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$504 t$4662 net1247 VGND VGND VPWR VPWR booth_b6_m43 sky130_fd_sc_hd__xor2_1
XFILLER_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$515 net1691 net432 net1683 net714 VGND VGND VPWR VPWR t$4668 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$676 final_adder.p_new$700 final_adder.p_new$684 VGND VGND VPWR VPWR
+ final_adder.p_new$804 sky130_fd_sc_hd__and2_1
XTAP_3958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$526 t$4673 net1247 VGND VGND VPWR VPWR booth_b6_m54 sky130_fd_sc_hd__xor2_1
XFILLER_84_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$687 final_adder.p_new$694 final_adder.g_new$711 final_adder.g_new$695
+ VGND VGND VPWR VPWR final_adder.g_new$815 sky130_fd_sc_hd__a21o_1
XTAP_3969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$698 final_adder.p_new$722 final_adder.p_new$706 VGND VGND VPWR VPWR
+ final_adder.p_new$826 sky130_fd_sc_hd__and2_1
XFILLER_45_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$537 net1582 net432 net1555 net714 VGND VGND VPWR VPWR t$4679 sky130_fd_sc_hd__a22o_1
XU$$548 net1246 VGND VGND VPWR VPWR notblock$4685\[0\] sky130_fd_sc_hd__inv_1
XU$$559 t$4691 net1239 VGND VGND VPWR VPWR booth_b8_m2 sky130_fd_sc_hd__xor2_1
XFILLER_147_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_878 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_994 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_62_0 s$581 c$1458 c$1460 VGND VGND VPWR VPWR c$2334 s$2335 sky130_fd_sc_hd__fa_1
X_0290_ clknet_leaf_199_clk booth_b20_m53 VGND VGND VPWR VPWR pp_row73_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_47_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_4_9_0 pp_row9_0 pp_row9_1 VGND VGND VPWR VPWR c$2752 s$2753 sky130_fd_sc_hd__ha_1
XU$$1210 net1630 net650 net1621 net923 VGND VGND VPWR VPWR t$5023 sky130_fd_sc_hd__a22o_1
XU$$1221 t$5028 net1012 VGND VGND VPWR VPWR booth_b16_m59 sky130_fd_sc_hd__xor2_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1232 net1013 VGND VGND VPWR VPWR notsign$5034 sky130_fd_sc_hd__inv_1
XFILLER_189_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1243 net1126 net638 net1036 net911 VGND VGND VPWR VPWR t$5041 sky130_fd_sc_hd__a22o_1
XU$$1254 t$5046 net1662 VGND VGND VPWR VPWR booth_b18_m7 sky130_fd_sc_hd__xor2_1
XU$$1265 net1201 net635 net1192 net908 VGND VGND VPWR VPWR t$5052 sky130_fd_sc_hd__a22o_1
XU$$1276 t$5057 net1664 VGND VGND VPWR VPWR booth_b18_m18 sky130_fd_sc_hd__xor2_1
XU$$1287 net1090 net636 net1080 net909 VGND VGND VPWR VPWR t$5063 sky130_fd_sc_hd__a22o_1
XFILLER_15_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1298 t$5068 net1663 VGND VGND VPWR VPWR booth_b18_m29 sky130_fd_sc_hd__xor2_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_176_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1813_ clknet_leaf_25_clk booth_b36_m13 VGND VGND VPWR VPWR pp_row49_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_191_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1744_ clknet_leaf_237_clk booth_b14_m33 VGND VGND VPWR VPWR pp_row47_7 sky130_fd_sc_hd__dfxtp_1
XU$$4439_1840 VGND VGND VPWR VPWR U$$4439_1840/HI net1840 sky130_fd_sc_hd__conb_1
XFILLER_8_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_84_1 s$3195 s$3197 s$3199 VGND VGND VPWR VPWR c$3734 s$3735 sky130_fd_sc_hd__fa_2
XFILLER_50_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1070 final_adder.$signal$1199 final_adder.g_new$1035 VGND VGND VPWR
+ VPWR net267 sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$1081 final_adder.$signal$1210 final_adder.g_new$971 VGND VGND VPWR
+ VPWR net280 sky130_fd_sc_hd__xor2_2
X_1675_ clknet_leaf_22_clk booth_b40_m4 VGND VGND VPWR VPWR pp_row44_20 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_77_0 c$3146 c$3148 c$3150 VGND VGND VPWR VPWR c$3704 s$3705 sky130_fd_sc_hd__fa_1
XFILLER_144_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0626_ clknet_leaf_176_clk booth_b38_m46 VGND VGND VPWR VPWR pp_row84_10 sky130_fd_sc_hd__dfxtp_1
Xfanout806 net807 VGND VGND VPWR VPWR net806 sky130_fd_sc_hd__buf_4
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout817 net823 VGND VGND VPWR VPWR net817 sky130_fd_sc_hd__buf_6
XFILLER_113_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout828 net829 VGND VGND VPWR VPWR net828 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_76_8 c$192 c$194 s$197 VGND VGND VPWR VPWR c$832 s$833 sky130_fd_sc_hd__fa_2
X_0557_ clknet_leaf_189_clk booth_b62_m19 VGND VGND VPWR VPWR pp_row81_23 sky130_fd_sc_hd__dfxtp_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout839 net841 VGND VGND VPWR VPWR net839 sky130_fd_sc_hd__buf_4
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_69_7 c$140 c$142 s$145 VGND VGND VPWR VPWR c$704 s$705 sky130_fd_sc_hd__fa_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0488_ clknet_leaf_129_clk booth_b60_m55 VGND VGND VPWR VPWR pp_row115_5 sky130_fd_sc_hd__dfxtp_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2227_ clknet_leaf_136_clk booth_b50_m60 VGND VGND VPWR VPWR pp_row110_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_27_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2158_ clknet_leaf_215_clk booth_b16_m44 VGND VGND VPWR VPWR pp_row60_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1109_ clknet_leaf_13_clk booth_b12_m2 VGND VGND VPWR VPWR pp_row14_6 sky130_fd_sc_hd__dfxtp_1
XU$$3190 t$6035 net1349 VGND VGND VPWR VPWR booth_b46_m16 sky130_fd_sc_hd__xor2_1
X_2089_ clknet_leaf_37_clk booth_b16_m42 VGND VGND VPWR VPWR pp_row58_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_53_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_100_3 s$1927 s$1929 s$1931 VGND VGND VPWR VPWR c$2644 s$2645 sky130_fd_sc_hd__fa_1
Xdadda_fa_1_95_0 pp_row95_0 pp_row95_1 pp_row95_2 VGND VGND VPWR VPWR c$1046 s$1047
+ sky130_fd_sc_hd__fa_1
XFILLER_1_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_558 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_2_108_0 net1917 pp_row108_1 VGND VGND VPWR VPWR c$1972 s$1973 sky130_fd_sc_hd__ha_1
XFILLER_188_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$440 final_adder.p_new$446 final_adder.p_new$442 VGND VGND VPWR VPWR
+ final_adder.p_new$568 sky130_fd_sc_hd__and2_1
XTAP_3722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$451 final_adder.p_new$452 final_adder.g_new$457 final_adder.g_new$453
+ VGND VGND VPWR VPWR final_adder.g_new$579 sky130_fd_sc_hd__a21o_1
XTAP_3733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$301 t$4559 net1279 VGND VGND VPWR VPWR booth_b4_m10 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$462 final_adder.p_new$468 final_adder.p_new$464 VGND VGND VPWR VPWR
+ final_adder.p_new$590 sky130_fd_sc_hd__and2_1
Xdadda_fa_6_107_0 c$3820 c$3822 s$3825 VGND VGND VPWR VPWR c$4110 s$4111 sky130_fd_sc_hd__fa_1
XTAP_3744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$312 net1170 net532 net1161 net805 VGND VGND VPWR VPWR t$4565 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$473 final_adder.p_new$474 final_adder.g_new$479 final_adder.g_new$475
+ VGND VGND VPWR VPWR final_adder.g_new$601 sky130_fd_sc_hd__a21o_1
XTAP_3755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$323 t$4570 net1274 VGND VGND VPWR VPWR booth_b4_m21 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$484 final_adder.p_new$490 final_adder.p_new$486 VGND VGND VPWR VPWR
+ final_adder.p_new$612 sky130_fd_sc_hd__and2_1
XTAP_3766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$334 net1063 net527 net1055 net800 VGND VGND VPWR VPWR t$4576 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$495 final_adder.p_new$496 final_adder.g_new$501 final_adder.g_new$497
+ VGND VGND VPWR VPWR final_adder.g_new$623 sky130_fd_sc_hd__a21o_1
XTAP_3777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$345 t$4581 net1279 VGND VGND VPWR VPWR booth_b4_m32 sky130_fd_sc_hd__xor2_1
XFILLER_189_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$356 net956 net527 net948 net800 VGND VGND VPWR VPWR t$4587 sky130_fd_sc_hd__a22o_1
XTAP_3799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_27_3 c$1066 s$1069 s$1071 VGND VGND VPWR VPWR c$2060 s$2061 sky130_fd_sc_hd__fa_1
XU$$367 t$4592 net1274 VGND VGND VPWR VPWR booth_b4_m43 sky130_fd_sc_hd__xor2_1
XFILLER_45_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$378 net1691 net533 net1682 net806 VGND VGND VPWR VPWR t$4598 sky130_fd_sc_hd__a22o_1
XFILLER_32_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$389 t$4603 net1280 VGND VGND VPWR VPWR booth_b4_m54 sky130_fd_sc_hd__xor2_1
XFILLER_189_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_94_0 c$3768 c$3770 s$3773 VGND VGND VPWR VPWR c$4084 s$4085 sky130_fd_sc_hd__fa_1
XFILLER_173_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1460_ clknet_leaf_40_clk booth_b6_m30 VGND VGND VPWR VPWR pp_row36_3 sky130_fd_sc_hd__dfxtp_1
X_0411_ clknet_leaf_125_clk booth_b64_m50 VGND VGND VPWR VPWR pp_row114_8 sky130_fd_sc_hd__dfxtp_1
X_1391_ clknet_leaf_244_clk net182 VGND VGND VPWR VPWR pp_row32_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_80_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0342_ clknet_leaf_202_clk booth_b58_m16 VGND VGND VPWR VPWR pp_row74_25 sky130_fd_sc_hd__dfxtp_1
XFILLER_95_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4469_1855 VGND VGND VPWR VPWR U$$4469_1855/HI net1855 sky130_fd_sc_hd__conb_1
X_0273_ clknet_leaf_226_clk booth_b52_m20 VGND VGND VPWR VPWR pp_row72_23 sky130_fd_sc_hd__dfxtp_1
XFILLER_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2012_ clknet_leaf_83_clk booth_b0_m56 VGND VGND VPWR VPWR pp_row56_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_23_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$890 net1023 net393 net1015 net659 VGND VGND VPWR VPWR t$4860 sky130_fd_sc_hd__a22o_1
XFILLER_91_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1040 t$4936 net1186 VGND VGND VPWR VPWR booth_b14_m37 sky130_fd_sc_hd__xor2_1
XU$$1051 net1741 net388 net1733 net654 VGND VGND VPWR VPWR t$4942 sky130_fd_sc_hd__a22o_1
XU$$1062 t$4947 net1190 VGND VGND VPWR VPWR booth_b14_m48 sky130_fd_sc_hd__xor2_1
XFILLER_189_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1073 net1633 net392 net1623 net658 VGND VGND VPWR VPWR t$4953 sky130_fd_sc_hd__a22o_1
XU$$1084 t$4958 net1188 VGND VGND VPWR VPWR booth_b14_m59 sky130_fd_sc_hd__xor2_1
XFILLER_52_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1095 net1188 VGND VGND VPWR VPWR notsign$4964 sky130_fd_sc_hd__inv_1
XFILLER_148_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_864 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1727_ clknet_leaf_123_clk booth_b56_m50 VGND VGND VPWR VPWR pp_row106_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1658_ clknet_leaf_6_clk booth_b10_m34 VGND VGND VPWR VPWR pp_row44_5 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_81_6 pp_row81_18 pp_row81_19 pp_row81_20 VGND VGND VPWR VPWR c$918 s$919
+ sky130_fd_sc_hd__fa_1
XFILLER_171_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout603 net604 VGND VGND VPWR VPWR net603 sky130_fd_sc_hd__clkbuf_4
X_0609_ clknet_leaf_174_clk booth_b58_m25 VGND VGND VPWR VPWR pp_row83_20 sky130_fd_sc_hd__dfxtp_1
Xfanout614 net615 VGND VGND VPWR VPWR net614 sky130_fd_sc_hd__buf_2
Xdadda_fa_1_74_5 pp_row74_23 pp_row74_24 pp_row74_25 VGND VGND VPWR VPWR c$790 s$791
+ sky130_fd_sc_hd__fa_1
X_1589_ clknet_leaf_9_clk booth_b24_m17 VGND VGND VPWR VPWR pp_row41_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_86_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout625 sel_0$4477 VGND VGND VPWR VPWR net625 sky130_fd_sc_hd__clkbuf_4
Xfanout636 net639 VGND VGND VPWR VPWR net636 sky130_fd_sc_hd__buf_6
Xfanout647 sel_0$4967 VGND VGND VPWR VPWR net647 sky130_fd_sc_hd__buf_4
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout658 sel_1$4898 VGND VGND VPWR VPWR net658 sky130_fd_sc_hd__buf_8
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_67_4 pp_row67_30 pp_row67_31 pp_row67_32 VGND VGND VPWR VPWR c$662 s$663
+ sky130_fd_sc_hd__fa_1
Xfanout669 net674 VGND VGND VPWR VPWR net669 sky130_fd_sc_hd__buf_4
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_37_2 s$2137 s$2139 s$2141 VGND VGND VPWR VPWR c$2916 s$2917 sky130_fd_sc_hd__fa_1
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_0_63_5 pp_row63_15 pp_row63_16 VGND VGND VPWR VPWR c$82 s$83 sky130_fd_sc_hd__ha_1
XFILLER_190_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_62_3 pp_row62_9 pp_row62_10 pp_row62_11 VGND VGND VPWR VPWR c$66 s$67
+ sky130_fd_sc_hd__fa_1
XFILLER_77_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3904 net1028 net463 net1020 net736 VGND VGND VPWR VPWR t$6400 sky130_fd_sc_hd__a22o_1
XU$$3915 t$6405 net1297 VGND VGND VPWR VPWR booth_b56_m36 sky130_fd_sc_hd__xor2_1
XFILLER_58_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3926 net1750 net466 net1742 net739 VGND VGND VPWR VPWR t$6411 sky130_fd_sc_hd__a22o_1
XTAP_4275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3937 t$6416 net1298 VGND VGND VPWR VPWR booth_b56_m47 sky130_fd_sc_hd__xor2_1
XTAP_3530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3948 net1643 net462 net1634 net735 VGND VGND VPWR VPWR t$6422 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$270 final_adder.p_new$272 final_adder.p_new$270 VGND VGND VPWR VPWR
+ final_adder.p_new$398 sky130_fd_sc_hd__and2_1
XTAP_4297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$281 final_adder.p_new$280 final_adder.g_new$283 final_adder.g_new$281
+ VGND VGND VPWR VPWR final_adder.g_new$409 sky130_fd_sc_hd__a21o_1
XFILLER_40_1076 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_32_1 c$1102 c$1104 c$1106 VGND VGND VPWR VPWR c$2096 s$2097 sky130_fd_sc_hd__fa_2
XFILLER_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$120 net1607 net450 net1599 net692 VGND VGND VPWR VPWR t$4467 sky130_fd_sc_hd__a22o_1
XTAP_3563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$131 t$4472 net1570 VGND VGND VPWR VPWR booth_b0_m62 sky130_fd_sc_hd__xor2_1
XU$$3959 t$6427 net1297 VGND VGND VPWR VPWR booth_b56_m58 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$292 final_adder.p_new$294 final_adder.p_new$292 VGND VGND VPWR VPWR
+ final_adder.p_new$420 sky130_fd_sc_hd__and2_1
XU$$142 net23 net1571 VGND VGND VPWR VPWR sel_1$4478 sky130_fd_sc_hd__xor2_4
XFILLER_45_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$153 net1675 net624 net1565 net897 VGND VGND VPWR VPWR t$4484 sky130_fd_sc_hd__a22o_1
XTAP_3585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$164 t$4489 net1390 VGND VGND VPWR VPWR booth_b2_m10 sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_25_0 pp_row25_5 pp_row25_6 pp_row25_7 VGND VGND VPWR VPWR c$2038 s$2039
+ sky130_fd_sc_hd__fa_1
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$175 net1166 net620 net1157 net893 VGND VGND VPWR VPWR t$4495 sky130_fd_sc_hd__a22o_1
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$186 t$4500 net1389 VGND VGND VPWR VPWR booth_b2_m21 sky130_fd_sc_hd__xor2_1
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$197 net1063 net619 net1055 net892 VGND VGND VPWR VPWR t$4506 sky130_fd_sc_hd__a22o_1
XFILLER_60_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0960_ clknet_leaf_185_clk net254 VGND VGND VPWR VPWR pp_row98_17 sky130_fd_sc_hd__dfxtp_4
XFILLER_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_984 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0891_ clknet_leaf_100_clk booth_b48_m47 VGND VGND VPWR VPWR pp_row95_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_158_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_91_5 c$1024 s$1027 s$1029 VGND VGND VPWR VPWR c$1828 s$1829 sky130_fd_sc_hd__fa_1
XFILLER_126_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1512_ clknet_leaf_44_clk booth_b16_m22 VGND VGND VPWR VPWR pp_row38_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_84_4 s$953 s$955 s$957 VGND VGND VPWR VPWR c$1742 s$1743 sky130_fd_sc_hd__fa_1
X_2492_ clknet_leaf_90_clk booth_b24_m45 VGND VGND VPWR VPWR pp_row69_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_126_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1443_ clknet_leaf_55_clk booth_b12_m23 VGND VGND VPWR VPWR pp_row35_6 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_77_3 c$832 s$835 s$837 VGND VGND VPWR VPWR c$1656 s$1657 sky130_fd_sc_hd__fa_1
XFILLER_68_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1374_ clknet_leaf_9_clk booth_b4_m28 VGND VGND VPWR VPWR pp_row32_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_68_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_47_1 s$2973 s$2975 s$2977 VGND VGND VPWR VPWR c$3586 s$3587 sky130_fd_sc_hd__fa_1
X_0325_ clknet_leaf_199_clk booth_b26_m48 VGND VGND VPWR VPWR pp_row74_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_83_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0256_ clknet_leaf_209_clk booth_b20_m52 VGND VGND VPWR VPWR pp_row72_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_51_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0187_ clknet_leaf_148_clk booth_b18_m52 VGND VGND VPWR VPWR pp_row70_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_36_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_100_2 pp_row100_6 pp_row100_7 pp_row100_8 VGND VGND VPWR VPWR c$1928 s$1929
+ sky130_fd_sc_hd__fa_1
XFILLER_91_692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_121_1 c$3408 c$3410 s$3413 VGND VGND VPWR VPWR c$3882 s$3883 sky130_fd_sc_hd__fa_1
XFILLER_17_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_114_0 c$3368 c$3370 c$3372 VGND VGND VPWR VPWR c$3852 s$3853 sky130_fd_sc_hd__fa_1
XFILLER_178_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout400 sel_0$4827 VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__buf_6
Xclkbuf_2_2_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_2_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_133_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout411 net412 VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__buf_4
Xfanout1409 net1411 VGND VGND VPWR VPWR net1409 sky130_fd_sc_hd__buf_6
XFILLER_99_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout422 net425 VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_72_2 pp_row72_17 pp_row72_18 pp_row72_19 VGND VGND VPWR VPWR c$748 s$749
+ sky130_fd_sc_hd__fa_1
Xfanout433 sel_0$4617 VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__buf_6
XFILLER_171_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout444 net445 VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__buf_4
Xfanout455 net458 VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_65_1 pp_row65_21 pp_row65_22 pp_row65_23 VGND VGND VPWR VPWR c$620 s$621
+ sky130_fd_sc_hd__fa_1
Xfanout466 net467 VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout477 net479 VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__buf_4
XFILLER_19_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout488 net492 VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__buf_4
Xdadda_fa_4_42_0 s$1241 c$2166 c$2168 VGND VGND VPWR VPWR c$2942 s$2943 sky130_fd_sc_hd__fa_1
XFILLER_74_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout499 net500 VGND VGND VPWR VPWR net499 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_58_0 pp_row58_11 pp_row58_12 pp_row58_13 VGND VGND VPWR VPWR c$492 s$493
+ sky130_fd_sc_hd__fa_2
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1809 net1224 net596 net1216 net869 VGND VGND VPWR VPWR t$5330 sky130_fd_sc_hd__a22o_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_948 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_94_3 s$1859 s$1861 s$1863 VGND VGND VPWR VPWR c$2596 s$2597 sky130_fd_sc_hd__fa_1
XFILLER_124_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_87_2 c$1768 s$1771 s$1773 VGND VGND VPWR VPWR c$2538 s$2539 sky130_fd_sc_hd__fa_1
Xdadda_ha_0_54_1 pp_row54_3 pp_row54_4 VGND VGND VPWR VPWR c$6 s$7 sky130_fd_sc_hd__ha_1
Xdadda_fa_6_57_0 c$3620 c$3622 s$3625 VGND VGND VPWR VPWR c$4010 s$4011 sky130_fd_sc_hd__fa_1
XFILLER_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4402 net1563 sel_0$6647 net125 net695 VGND VGND VPWR VPWR t$6655 sky130_fd_sc_hd__a22o_1
XU$$4413 t$6660 net1827 VGND VGND VPWR VPWR booth_b64_m11 sky130_fd_sc_hd__xor2_1
XFILLER_93_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4424 net1159 sel_0$6647 net1152 net693 VGND VGND VPWR VPWR t$6666 sky130_fd_sc_hd__a22o_1
XFILLER_49_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_0_60_0 pp_row60_0 pp_row60_1 pp_row60_2 VGND VGND VPWR VPWR c$40 s$41 sky130_fd_sc_hd__fa_1
XU$$4435 t$6671 net1838 VGND VGND VPWR VPWR booth_b64_m22 sky130_fd_sc_hd__xor2_1
XU$$4446 net84 sel_0$6647 net1054 net698 VGND VGND VPWR VPWR t$6677 sky130_fd_sc_hd__a22o_1
XFILLER_64_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3701 net1301 VGND VGND VPWR VPWR notblock$6295\[2\] sky130_fd_sc_hd__inv_1
XTAP_4050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3712 t$6302 net1305 VGND VGND VPWR VPWR booth_b54_m3 sky130_fd_sc_hd__xor2_1
XTAP_4061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4457 t$6682 net1849 VGND VGND VPWR VPWR booth_b64_m33 sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_116_2 pp_row116_8 c$2746 s$2749 VGND VGND VPWR VPWR c$3390 s$3391 sky130_fd_sc_hd__fa_2
XTAP_4072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4468 net954 sel_0$6647 net945 net699 VGND VGND VPWR VPWR t$6688 sky130_fd_sc_hd__a22o_1
XU$$3723 net1507 net468 net1498 net741 VGND VGND VPWR VPWR t$6308 sky130_fd_sc_hd__a22o_1
Xclkbuf_5_24__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_5_24__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_1090_ clknet_leaf_58_clk booth_b12_m0 VGND VGND VPWR VPWR pp_row12_6 sky130_fd_sc_hd__dfxtp_1
XU$$3734 t$6313 net1304 VGND VGND VPWR VPWR booth_b54_m14 sky130_fd_sc_hd__xor2_1
XU$$4479 t$6693 net1860 VGND VGND VPWR VPWR booth_b64_m44 sky130_fd_sc_hd__xor2_1
XTAP_4083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3745 net1136 net468 net1120 net741 VGND VGND VPWR VPWR t$6319 sky130_fd_sc_hd__a22o_1
XTAP_4094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3756 t$6324 net1301 VGND VGND VPWR VPWR booth_b54_m25 sky130_fd_sc_hd__xor2_1
XU$$3767 net1028 net469 net1020 net742 VGND VGND VPWR VPWR t$6330 sky130_fd_sc_hd__a22o_1
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_109_1 c$2706 c$2708 s$2711 VGND VGND VPWR VPWR c$3346 s$3347 sky130_fd_sc_hd__fa_1
XTAP_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3778 t$6335 net1306 VGND VGND VPWR VPWR booth_b54_m36 sky130_fd_sc_hd__xor2_1
XTAP_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3789 net1750 net474 net1742 net747 VGND VGND VPWR VPWR t$6341 sky130_fd_sc_hd__a22o_1
XFILLER_166_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_360 net997 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_371 net1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_382 net1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_393 net1530 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1992_ clknet_leaf_69_clk booth_b22_m33 VGND VGND VPWR VPWR pp_row55_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_14_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0943_ clknet_leaf_130_clk booth_b58_m63 VGND VGND VPWR VPWR pp_row121_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0874_ clknet_leaf_93_clk booth_b56_m38 VGND VGND VPWR VPWR pp_row94_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_134_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_82_1 c$906 c$908 c$910 VGND VGND VPWR VPWR c$1712 s$1713 sky130_fd_sc_hd__fa_1
XFILLER_138_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2475_ clknet_leaf_99_clk booth_b58_m10 VGND VGND VPWR VPWR pp_row68_28 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_75_0 s$195 c$780 c$782 VGND VGND VPWR VPWR c$1626 s$1627 sky130_fd_sc_hd__fa_1
XFILLER_114_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1426_ clknet_leaf_64_clk booth_b22_m12 VGND VGND VPWR VPWR pp_row34_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_69_987 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1357_ clknet_leaf_2_clk booth_b8_m23 VGND VGND VPWR VPWR pp_row31_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_51_7 pp_row51_21 pp_row51_22 pp_row51_23 VGND VGND VPWR VPWR c$380 s$381
+ sky130_fd_sc_hd__fa_1
X_0308_ clknet_leaf_226_clk booth_b54_m19 VGND VGND VPWR VPWR pp_row73_23 sky130_fd_sc_hd__dfxtp_1
X_1288_ clknet_leaf_1_clk booth_b14_m13 VGND VGND VPWR VPWR pp_row27_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_83_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0239_ clknet_leaf_150_clk booth_b50_m21 VGND VGND VPWR VPWR pp_row71_22 sky130_fd_sc_hd__dfxtp_1
XFILLER_52_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_97_1 c$2610 c$2612 s$2615 VGND VGND VPWR VPWR c$3274 s$3275 sky130_fd_sc_hd__fa_1
XFILLER_4_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_74_0 s$3695 c$4042 s$4045 VGND VGND VPWR VPWR c$4300 s$4301 sky130_fd_sc_hd__fa_1
XFILLER_146_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1206 net1208 VGND VGND VPWR VPWR net1206 sky130_fd_sc_hd__buf_6
Xfanout1217 net1218 VGND VGND VPWR VPWR net1217 sky130_fd_sc_hd__buf_4
XFILLER_121_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1228 net1229 VGND VGND VPWR VPWR net1228 sky130_fd_sc_hd__buf_4
Xfanout1239 net1243 VGND VGND VPWR VPWR net1239 sky130_fd_sc_hd__buf_6
XFILLER_75_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3008 t$5941 net1374 VGND VGND VPWR VPWR booth_b42_m62 sky130_fd_sc_hd__xor2_1
XU$$3019 net39 net1370 VGND VGND VPWR VPWR sel_1$5948 sky130_fd_sc_hd__xor2_1
XFILLER_74_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2307 t$5583 net1435 VGND VGND VPWR VPWR booth_b32_m54 sky130_fd_sc_hd__xor2_1
XU$$2318 net1584 net575 net1557 net848 VGND VGND VPWR VPWR t$5589 sky130_fd_sc_hd__a22o_1
XU$$2329 net1435 VGND VGND VPWR VPWR notblock$5595\[0\] sky130_fd_sc_hd__inv_1
XU$$1606 t$5225 net1484 VGND VGND VPWR VPWR booth_b22_m46 sky130_fd_sc_hd__xor2_1
XU$$1617 net1646 net616 net1638 net889 VGND VGND VPWR VPWR t$5231 sky130_fd_sc_hd__a22o_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1628 t$5236 net1481 VGND VGND VPWR VPWR booth_b22_m57 sky130_fd_sc_hd__xor2_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1639 net1536 net617 net1528 net890 VGND VGND VPWR VPWR t$5242 sky130_fd_sc_hd__a22o_1
XFILLER_15_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_789 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_92_0 s$1037 c$1818 c$1820 VGND VGND VPWR VPWR c$2574 s$2575 sky130_fd_sc_hd__fa_1
XFILLER_143_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_748 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0590_ clknet_leaf_186_clk booth_b22_m61 VGND VGND VPWR VPWR pp_row83_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_136_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2260_ clknet_leaf_137_clk booth_b56_m54 VGND VGND VPWR VPWR pp_row110_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1740 net101 VGND VGND VPWR VPWR net1740 sky130_fd_sc_hd__clkbuf_4
X_1211_ clknet_leaf_49_clk booth_b20_m2 VGND VGND VPWR VPWR pp_row22_10 sky130_fd_sc_hd__dfxtp_1
Xfanout1751 net1752 VGND VGND VPWR VPWR net1751 sky130_fd_sc_hd__buf_4
X_2191_ clknet_leaf_223_clk booth_b8_m53 VGND VGND VPWR VPWR pp_row61_4 sky130_fd_sc_hd__dfxtp_1
XU$$4210 net1710 net439 net1702 net721 VGND VGND VPWR VPWR t$6556 sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_54_5 s$431 s$433 s$435 VGND VGND VPWR VPWR c$1384 s$1385 sky130_fd_sc_hd__fa_1
Xdadda_fa_4_121_0 pp_row121_0 pp_row121_1 pp_row121_2 VGND VGND VPWR VPWR c$3412 s$3413
+ sky130_fd_sc_hd__fa_1
XU$$4221 t$6561 net1270 VGND VGND VPWR VPWR booth_b60_m52 sky130_fd_sc_hd__xor2_1
XU$$4232 net1601 net435 net1592 net717 VGND VGND VPWR VPWR t$6567 sky130_fd_sc_hd__a22o_1
X_1142_ clknet_leaf_11_clk booth_b12_m5 VGND VGND VPWR VPWR pp_row17_6 sky130_fd_sc_hd__dfxtp_1
XU$$4243 t$6572 net1266 VGND VGND VPWR VPWR booth_b60_m63 sky130_fd_sc_hd__xor2_1
XFILLER_65_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4254 t$6579 net1254 VGND VGND VPWR VPWR booth_b62_m0 sky130_fd_sc_hd__xor2_1
XU$$4265 net1567 net422 net1526 net704 VGND VGND VPWR VPWR t$6585 sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_47_4 s$303 s$305 s$307 VGND VGND VPWR VPWR c$1298 s$1299 sky130_fd_sc_hd__fa_2
XU$$3520 t$6203 net1334 VGND VGND VPWR VPWR booth_b50_m44 sky130_fd_sc_hd__xor2_1
XU$$3531 net1686 net490 net1661 net763 VGND VGND VPWR VPWR t$6209 sky130_fd_sc_hd__a22o_1
XU$$4276 t$6590 net1254 VGND VGND VPWR VPWR booth_b62_m11 sky130_fd_sc_hd__xor2_1
XFILLER_65_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3542 t$6214 net1336 VGND VGND VPWR VPWR booth_b50_m55 sky130_fd_sc_hd__xor2_1
XU$$4287 net1159 net418 net1152 net700 VGND VGND VPWR VPWR t$6596 sky130_fd_sc_hd__a22o_1
XFILLER_92_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4298 t$6601 net1255 VGND VGND VPWR VPWR booth_b62_m22 sky130_fd_sc_hd__xor2_1
XU$$3553 net1556 net491 net1549 net764 VGND VGND VPWR VPWR t$6220 sky130_fd_sc_hd__a22o_1
X_1073_ clknet_leaf_52_clk booth_b10_m0 VGND VGND VPWR VPWR pp_row10_5 sky130_fd_sc_hd__dfxtp_1
XU$$3564 net1321 VGND VGND VPWR VPWR notblock$6225\[2\] sky130_fd_sc_hd__inv_1
XU$$3575 t$6232 net1324 VGND VGND VPWR VPWR booth_b52_m3 sky130_fd_sc_hd__xor2_1
XU$$2830 net1747 net537 net1739 net810 VGND VGND VPWR VPWR t$5851 sky130_fd_sc_hd__a22o_1
XU$$2841 t$5856 net1379 VGND VGND VPWR VPWR booth_b40_m47 sky130_fd_sc_hd__xor2_1
XU$$3586 net1507 net479 net1498 net752 VGND VGND VPWR VPWR t$6238 sky130_fd_sc_hd__a22o_1
XU$$2852 net1644 net540 net1635 net813 VGND VGND VPWR VPWR t$5862 sky130_fd_sc_hd__a22o_1
XFILLER_34_843 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3597 t$6243 net1324 VGND VGND VPWR VPWR booth_b52_m14 sky130_fd_sc_hd__xor2_1
XU$$2863 t$5867 net1382 VGND VGND VPWR VPWR booth_b40_m58 sky130_fd_sc_hd__xor2_1
XFILLER_34_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2874 net1532 net541 net1784 net814 VGND VGND VPWR VPWR t$5873 sky130_fd_sc_hd__a22o_1
XU$$2885 net1227 net519 net1122 net792 VGND VGND VPWR VPWR t$5880 sky130_fd_sc_hd__a22o_1
XU$$2896 t$5885 net1367 VGND VGND VPWR VPWR booth_b42_m6 sky130_fd_sc_hd__xor2_1
XFILLER_178_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_190 net981 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1975_ clknet_leaf_72_clk booth_b50_m4 VGND VGND VPWR VPWR pp_row54_25 sky130_fd_sc_hd__dfxtp_1
XFILLER_119_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0926_ clknet_leaf_112_clk booth_b40_m57 VGND VGND VPWR VPWR pp_row97_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0857_ clknet_leaf_142_clk booth_b62_m31 VGND VGND VPWR VPWR pp_row93_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0788_ clknet_leaf_132_clk notsign$6364 VGND VGND VPWR VPWR pp_row119_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_143_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2458_ clknet_leaf_128_clk booth_b50_m62 VGND VGND VPWR VPWR pp_row112_2 sky130_fd_sc_hd__dfxtp_1
X_1409_ clknet_leaf_57_clk booth_b26_m7 VGND VGND VPWR VPWR pp_row33_13 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$803 final_adder.p_new$818 final_adder.g_new$851 final_adder.g_new$819
+ VGND VGND VPWR VPWR final_adder.g_new$931 sky130_fd_sc_hd__a21o_1
X_2389_ clknet_leaf_96_clk booth_b36_m30 VGND VGND VPWR VPWR pp_row66_18 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$825 final_adder.p_new$840 final_adder.g_new$753 final_adder.g_new$841
+ VGND VGND VPWR VPWR final_adder.g_new$953 sky130_fd_sc_hd__a21o_2
Xfinal_adder.U$$847 final_adder.p_new$878 final_adder.g_new$943 final_adder.g_new$879
+ VGND VGND VPWR VPWR final_adder.g_new$975 sky130_fd_sc_hd__a21o_2
XFILLER_112_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$708 t$4767 net1415 VGND VGND VPWR VPWR booth_b10_m8 sky130_fd_sc_hd__xor2_1
XFILLER_112_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$869 final_adder.p_new$900 final_adder.g_new$853 final_adder.g_new$901
+ VGND VGND VPWR VPWR final_adder.g_new$997 sky130_fd_sc_hd__a21o_1
XU$$719 net1194 net402 net1175 net668 VGND VGND VPWR VPWR t$4773 sky130_fd_sc_hd__a22o_1
Xdadda_fa_1_42_3 pp_row42_9 pp_row42_10 pp_row42_11 VGND VGND VPWR VPWR c$250 s$251
+ sky130_fd_sc_hd__fa_1
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_12_1 pp_row12_3 pp_row12_4 pp_row12_5 VGND VGND VPWR VPWR c$2764 s$2765
+ sky130_fd_sc_hd__fa_1
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_109_0 pp_row109_0 pp_row109_1 pp_row109_2 VGND VGND VPWR VPWR c$2710 s$2711
+ sky130_fd_sc_hd__fa_1
XFILLER_4_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1003 net1004 VGND VGND VPWR VPWR net1003 sky130_fd_sc_hd__buf_4
Xfanout1014 net9 VGND VGND VPWR VPWR net1014 sky130_fd_sc_hd__buf_6
XFILLER_120_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1025 net1026 VGND VGND VPWR VPWR net1025 sky130_fd_sc_hd__buf_4
Xfanout1036 net1038 VGND VGND VPWR VPWR net1036 sky130_fd_sc_hd__buf_4
XFILLER_66_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1047 net1048 VGND VGND VPWR VPWR net1047 sky130_fd_sc_hd__clkbuf_8
XFILLER_94_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_57_3 s$1415 s$1417 s$1419 VGND VGND VPWR VPWR c$2300 s$2301 sky130_fd_sc_hd__fa_1
Xfanout1058 net1059 VGND VGND VPWR VPWR net1058 sky130_fd_sc_hd__buf_6
XFILLER_47_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1069 net1070 VGND VGND VPWR VPWR net1069 sky130_fd_sc_hd__clkbuf_4
XFILLER_102_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2104 t$5480 net1441 VGND VGND VPWR VPWR booth_b30_m21 sky130_fd_sc_hd__xor2_1
XU$$2115 net1066 net581 net1057 net854 VGND VGND VPWR VPWR t$5486 sky130_fd_sc_hd__a22o_1
XU$$2126 t$5491 net1440 VGND VGND VPWR VPWR booth_b30_m32 sky130_fd_sc_hd__xor2_1
XU$$2137 net958 net582 net950 net855 VGND VGND VPWR VPWR t$5497 sky130_fd_sc_hd__a22o_1
XU$$2148 t$5502 net1440 VGND VGND VPWR VPWR booth_b30_m43 sky130_fd_sc_hd__xor2_1
XU$$1403 t$5122 net1488 VGND VGND VPWR VPWR booth_b20_m13 sky130_fd_sc_hd__xor2_1
XFILLER_188_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2159 net1688 net579 net1680 net852 VGND VGND VPWR VPWR t$5508 sky130_fd_sc_hd__a22o_1
XU$$1414 net1139 net627 net1131 net900 VGND VGND VPWR VPWR t$5128 sky130_fd_sc_hd__a22o_1
XFILLER_90_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1425 t$5133 net1486 VGND VGND VPWR VPWR booth_b20_m24 sky130_fd_sc_hd__xor2_1
XU$$1436 net1041 net631 net1025 net904 VGND VGND VPWR VPWR t$5139 sky130_fd_sc_hd__a22o_1
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1447 t$5144 net1489 VGND VGND VPWR VPWR booth_b20_m35 sky130_fd_sc_hd__xor2_1
XFILLER_187_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1023 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1458 net925 net628 net1745 net901 VGND VGND VPWR VPWR t$5150 sky130_fd_sc_hd__a22o_1
XU$$1469 t$5155 net1489 VGND VGND VPWR VPWR booth_b20_m46 sky130_fd_sc_hd__xor2_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1760_ clknet_leaf_23_clk booth_b44_m3 VGND VGND VPWR VPWR pp_row47_22 sky130_fd_sc_hd__dfxtp_1
XFILLER_128_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0711_ clknet_leaf_165_clk booth_b52_m35 VGND VGND VPWR VPWR pp_row87_15 sky130_fd_sc_hd__dfxtp_1
X_1691_ clknet_leaf_19_clk booth_b20_m25 VGND VGND VPWR VPWR pp_row45_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_116_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0642_ clknet_leaf_183_clk notsign$5174 VGND VGND VPWR VPWR pp_row85_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_131_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0573_ clknet_leaf_190_clk booth_b42_m40 VGND VGND VPWR VPWR pp_row82_13 sky130_fd_sc_hd__dfxtp_1
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2312_ clknet_leaf_87_clk booth_b28_m36 VGND VGND VPWR VPWR pp_row64_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_987 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2243_ clknet_leaf_150_clk booth_b38_m24 VGND VGND VPWR VPWR pp_row62_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_78_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_52_2 c$376 c$378 c$380 VGND VGND VPWR VPWR c$1354 s$1355 sky130_fd_sc_hd__fa_1
Xfanout1570 net1572 VGND VGND VPWR VPWR net1570 sky130_fd_sc_hd__buf_6
Xfanout1581 net119 VGND VGND VPWR VPWR net1581 sky130_fd_sc_hd__buf_4
Xfanout1592 net1593 VGND VGND VPWR VPWR net1592 sky130_fd_sc_hd__clkbuf_8
XFILLER_38_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2174_ clknet_leaf_224_clk booth_b42_m18 VGND VGND VPWR VPWR pp_row60_21 sky130_fd_sc_hd__dfxtp_1
XU$$4040 t$6469 net1284 VGND VGND VPWR VPWR booth_b58_m30 sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_45_1 pp_row45_20 pp_row45_21 pp_row45_22 VGND VGND VPWR VPWR c$1268 s$1269
+ sky130_fd_sc_hd__fa_1
XU$$4051 net979 net455 net970 net728 VGND VGND VPWR VPWR t$6475 sky130_fd_sc_hd__a22o_1
XU$$4062 t$6480 net1289 VGND VGND VPWR VPWR booth_b58_m41 sky130_fd_sc_hd__xor2_1
XU$$4073 net1708 net456 net1700 net729 VGND VGND VPWR VPWR t$6486 sky130_fd_sc_hd__a22o_1
XFILLER_53_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1125_ clknet_leaf_11_clk booth_b4_m12 VGND VGND VPWR VPWR pp_row16_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_81_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4084 t$6491 net1288 VGND VGND VPWR VPWR booth_b58_m52 sky130_fd_sc_hd__xor2_1
XFILLER_20_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3350 net1060 net494 net1051 net767 VGND VGND VPWR VPWR t$6117 sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_22_0 c$2816 c$2818 c$2820 VGND VGND VPWR VPWR c$3484 s$3485 sky130_fd_sc_hd__fa_1
XU$$4095 net1601 net456 net1592 net729 VGND VGND VPWR VPWR t$6497 sky130_fd_sc_hd__a22o_1
XU$$3361 t$6122 net1341 VGND VGND VPWR VPWR booth_b48_m33 sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_38_0 pp_row38_8 pp_row38_9 pp_row38_10 VGND VGND VPWR VPWR c$1182 s$1183
+ sky130_fd_sc_hd__fa_1
XFILLER_65_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3372 net951 net494 net943 net767 VGND VGND VPWR VPWR t$6128 sky130_fd_sc_hd__a22o_1
XU$$3383 t$6133 net1344 VGND VGND VPWR VPWR booth_b48_m44 sky130_fd_sc_hd__xor2_1
X_1056_ clknet_leaf_56_clk booth_b8_m0 VGND VGND VPWR VPWR pp_row8_4 sky130_fd_sc_hd__dfxtp_1
XU$$3394 net1684 net498 net1660 net771 VGND VGND VPWR VPWR t$6139 sky130_fd_sc_hd__a22o_1
XU$$2660 t$5764 net1395 VGND VGND VPWR VPWR booth_b38_m25 sky130_fd_sc_hd__xor2_1
XU$$2671 net1029 net547 net1021 net820 VGND VGND VPWR VPWR t$5770 sky130_fd_sc_hd__a22o_1
XFILLER_55_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2682 t$5775 net1394 VGND VGND VPWR VPWR booth_b38_m36 sky130_fd_sc_hd__xor2_1
XU$$2693 net1748 net546 net1740 net819 VGND VGND VPWR VPWR t$5781 sky130_fd_sc_hd__a22o_1
XFILLER_181_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1970 net1101 net587 net1091 net860 VGND VGND VPWR VPWR t$5412 sky130_fd_sc_hd__a22o_1
XU$$1981 t$5417 net1452 VGND VGND VPWR VPWR booth_b28_m28 sky130_fd_sc_hd__xor2_1
XU$$1992 net991 net586 net982 net859 VGND VGND VPWR VPWR t$5423 sky130_fd_sc_hd__a22o_1
XFILLER_21_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1958_ clknet_leaf_66_clk booth_b20_m34 VGND VGND VPWR VPWR pp_row54_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_193_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0909_ clknet_leaf_104_clk booth_b46_m50 VGND VGND VPWR VPWR pp_row96_8 sky130_fd_sc_hd__dfxtp_1
X_1889_ clknet_leaf_39_clk booth_b10_m42 VGND VGND VPWR VPWR pp_row52_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_162_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_67_2 s$2377 s$2379 s$2381 VGND VGND VPWR VPWR c$3096 s$3097 sky130_fd_sc_hd__fa_1
XFILLER_142_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput106 b[47] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__buf_6
Xinput117 b[57] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__buf_2
Xinput128 b[9] VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_2
Xinput139 c[109] VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_1
Xfinal_adder.U$$600 final_adder.p_new$612 final_adder.p_new$604 VGND VGND VPWR VPWR
+ final_adder.p_new$728 sky130_fd_sc_hd__and2_1
Xdadda_fa_7_37_0 s$3547 c$3968 s$3971 VGND VGND VPWR VPWR c$4226 s$4227 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$611 final_adder.p_new$614 final_adder.g_new$623 final_adder.g_new$615
+ VGND VGND VPWR VPWR final_adder.g_new$739 sky130_fd_sc_hd__a21o_1
XTAP_3904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$633 final_adder.p_new$640 final_adder.g_new$657 final_adder.g_new$641
+ VGND VGND VPWR VPWR final_adder.g_new$761 sky130_fd_sc_hd__a21o_1
XTAP_3915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$644 final_adder.p_new$668 final_adder.p_new$652 VGND VGND VPWR VPWR
+ final_adder.p_new$772 sky130_fd_sc_hd__and2_1
XTAP_3926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$655 final_adder.p_new$662 final_adder.g_new$679 final_adder.g_new$663
+ VGND VGND VPWR VPWR final_adder.g_new$783 sky130_fd_sc_hd__a21o_1
XTAP_3937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$666 final_adder.p_new$690 final_adder.p_new$674 VGND VGND VPWR VPWR
+ final_adder.p_new$794 sky130_fd_sc_hd__and2_1
XU$$505 net1729 net428 net1720 net710 VGND VGND VPWR VPWR t$4663 sky130_fd_sc_hd__a22o_1
XTAP_3948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$516 t$4668 net1251 VGND VGND VPWR VPWR booth_b6_m49 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$677 final_adder.p_new$684 final_adder.g_new$701 final_adder.g_new$685
+ VGND VGND VPWR VPWR final_adder.g_new$805 sky130_fd_sc_hd__a21o_1
Xdadda_fa_1_40_0 pp_row40_0 pp_row40_1 pp_row40_2 VGND VGND VPWR VPWR c$228 s$229
+ sky130_fd_sc_hd__fa_1
XTAP_3959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$688 final_adder.p_new$712 final_adder.p_new$696 VGND VGND VPWR VPWR
+ final_adder.p_new$816 sky130_fd_sc_hd__and2_1
XU$$527 net1620 net428 net1612 net710 VGND VGND VPWR VPWR t$4674 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$699 final_adder.p_new$706 final_adder.g_new$723 final_adder.g_new$707
+ VGND VGND VPWR VPWR final_adder.g_new$827 sky130_fd_sc_hd__a21o_1
XU$$538 t$4679 net1251 VGND VGND VPWR VPWR booth_b6_m60 sky130_fd_sc_hd__xor2_1
XU$$549 net63 VGND VGND VPWR VPWR notblock$4685\[1\] sky130_fd_sc_hd__inv_1
XFILLER_25_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_90 net530 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_1114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_62_1 c$1462 c$1464 c$1466 VGND VGND VPWR VPWR c$2336 s$2337 sky130_fd_sc_hd__fa_1
XFILLER_0_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_55_0 s$455 c$1374 c$1376 VGND VGND VPWR VPWR c$2278 s$2279 sky130_fd_sc_hd__fa_1
XFILLER_0_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_195_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_195_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_46_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1200 net1690 net650 net1682 net923 VGND VGND VPWR VPWR t$5018 sky130_fd_sc_hd__a22o_1
XFILLER_189_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1211 t$5023 net1014 VGND VGND VPWR VPWR booth_b16_m54 sky130_fd_sc_hd__xor2_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_960 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1222 net1578 net648 net1551 net921 VGND VGND VPWR VPWR t$5029 sky130_fd_sc_hd__a22o_1
XU$$1233 net1013 VGND VGND VPWR VPWR notblock$5035\[0\] sky130_fd_sc_hd__inv_1
XFILLER_50_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1244 t$5041 net1664 VGND VGND VPWR VPWR booth_b18_m2 sky130_fd_sc_hd__xor2_1
XFILLER_189_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1255 net1511 net635 net1503 net908 VGND VGND VPWR VPWR t$5047 sky130_fd_sc_hd__a22o_1
XU$$1266 t$5052 net1662 VGND VGND VPWR VPWR booth_b18_m13 sky130_fd_sc_hd__xor2_1
XFILLER_149_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1277 net1139 net637 net1130 net910 VGND VGND VPWR VPWR t$5058 sky130_fd_sc_hd__a22o_1
XFILLER_188_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1288 t$5063 net1663 VGND VGND VPWR VPWR booth_b18_m24 sky130_fd_sc_hd__xor2_1
XU$$1299 net1040 net636 net1023 net909 VGND VGND VPWR VPWR t$5069 sky130_fd_sc_hd__a22o_1
XFILLER_176_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1812_ clknet_leaf_26_clk booth_b34_m15 VGND VGND VPWR VPWR pp_row49_17 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_7_112_0 s$3847 c$4118 s$4121 VGND VGND VPWR VPWR c$4376 s$4377 sky130_fd_sc_hd__fa_1
XFILLER_30_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1743_ clknet_leaf_237_clk booth_b12_m35 VGND VGND VPWR VPWR pp_row47_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1060 final_adder.$signal$1189 final_adder.g_new$1040 VGND VGND VPWR
+ VPWR net383 sky130_fd_sc_hd__xor2_1
X_1674_ clknet_leaf_240_clk booth_b38_m6 VGND VGND VPWR VPWR pp_row44_19 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$1071 final_adder.$signal$1200 final_adder.g_new$981 VGND VGND VPWR
+ VPWR net269 sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$1082 final_adder.$signal$1211 final_adder.g_new$1029 VGND VGND VPWR
+ VPWR net281 sky130_fd_sc_hd__xor2_2
Xdadda_fa_5_77_1 s$3153 s$3155 s$3157 VGND VGND VPWR VPWR c$3706 s$3707 sky130_fd_sc_hd__fa_1
XFILLER_89_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0625_ clknet_leaf_176_clk booth_b36_m48 VGND VGND VPWR VPWR pp_row84_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_144_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout807 sel_1$4548 VGND VGND VPWR VPWR net807 sky130_fd_sc_hd__buf_4
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0556_ clknet_leaf_189_clk booth_b60_m21 VGND VGND VPWR VPWR pp_row81_22 sky130_fd_sc_hd__dfxtp_1
Xfanout818 net819 VGND VGND VPWR VPWR net818 sky130_fd_sc_hd__buf_6
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout829 net831 VGND VGND VPWR VPWR net829 sky130_fd_sc_hd__buf_6
XFILLER_112_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0487_ clknet_leaf_205_clk booth_b42_m37 VGND VGND VPWR VPWR pp_row79_14 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_69_8 s$147 s$149 s$151 VGND VGND VPWR VPWR c$706 s$707 sky130_fd_sc_hd__fa_2
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2226_ clknet_leaf_227_clk booth_b8_m54 VGND VGND VPWR VPWR pp_row62_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_39_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_186_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_186_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_39_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2157_ clknet_leaf_215_clk booth_b14_m46 VGND VGND VPWR VPWR pp_row60_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_81_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1108_ clknet_leaf_13_clk booth_b10_m4 VGND VGND VPWR VPWR pp_row14_5 sky130_fd_sc_hd__dfxtp_1
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2088_ clknet_leaf_37_clk booth_b14_m44 VGND VGND VPWR VPWR pp_row58_7 sky130_fd_sc_hd__dfxtp_1
XU$$3180 t$6030 net1354 VGND VGND VPWR VPWR booth_b46_m11 sky130_fd_sc_hd__xor2_1
XU$$3191 net1159 net501 net1151 net774 VGND VGND VPWR VPWR t$6036 sky130_fd_sc_hd__a22o_1
Xdadda_fa_6_9_0 c$3428 c$3430 s$3433 VGND VGND VPWR VPWR c$3914 s$3915 sky130_fd_sc_hd__fa_1
XFILLER_179_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1039_ clknet_leaf_248_clk net212 VGND VGND VPWR VPWR pp_row5_3 sky130_fd_sc_hd__dfxtp_4
XU$$2490 net1504 net551 net1497 net824 VGND VGND VPWR VPWR t$5678 sky130_fd_sc_hd__a22o_1
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_840 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_110_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_110_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_174_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_72_0 s$1601 c$2406 c$2408 VGND VGND VPWR VPWR c$3122 s$3123 sky130_fd_sc_hd__fa_1
XFILLER_116_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_88_0 net1900 pp_row88_1 pp_row88_2 VGND VGND VPWR VPWR c$1000 s$1001 sky130_fd_sc_hd__fa_1
XFILLER_107_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_5_5__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_5_5__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_3701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$430 final_adder.p_new$436 final_adder.p_new$432 VGND VGND VPWR VPWR
+ final_adder.p_new$558 sky130_fd_sc_hd__and2_1
XFILLER_188_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$441 final_adder.p_new$442 final_adder.g_new$447 final_adder.g_new$443
+ VGND VGND VPWR VPWR final_adder.g_new$569 sky130_fd_sc_hd__a21o_1
XTAP_3723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$452 final_adder.p_new$458 final_adder.p_new$454 VGND VGND VPWR VPWR
+ final_adder.p_new$580 sky130_fd_sc_hd__and2_1
XTAP_3734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_177_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_177_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_85_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$302 net1221 net532 net1211 net805 VGND VGND VPWR VPWR t$4560 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$463 final_adder.p_new$464 final_adder.g_new$469 final_adder.g_new$465
+ VGND VGND VPWR VPWR final_adder.g_new$591 sky130_fd_sc_hd__a21o_1
XTAP_3745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$313 t$4565 net1279 VGND VGND VPWR VPWR booth_b4_m16 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$474 final_adder.p_new$480 final_adder.p_new$476 VGND VGND VPWR VPWR
+ final_adder.p_new$602 sky130_fd_sc_hd__and2_1
XTAP_3756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$324 net1105 net527 net1097 net800 VGND VGND VPWR VPWR t$4571 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$485 final_adder.p_new$486 final_adder.g_new$491 final_adder.g_new$487
+ VGND VGND VPWR VPWR final_adder.g_new$613 sky130_fd_sc_hd__a21o_1
XTAP_3767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$496 final_adder.p_new$502 final_adder.p_new$498 VGND VGND VPWR VPWR
+ final_adder.p_new$624 sky130_fd_sc_hd__and2_1
XU$$335 t$4576 net1273 VGND VGND VPWR VPWR booth_b4_m27 sky130_fd_sc_hd__xor2_1
XFILLER_29_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$346 net998 net527 net990 net800 VGND VGND VPWR VPWR t$4582 sky130_fd_sc_hd__a22o_1
XFILLER_45_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$357 t$4587 net1273 VGND VGND VPWR VPWR booth_b4_m38 sky130_fd_sc_hd__xor2_1
XFILLER_189_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$368 net1729 net529 net1720 net802 VGND VGND VPWR VPWR t$4593 sky130_fd_sc_hd__a22o_1
XU$$379 t$4598 net1280 VGND VGND VPWR VPWR booth_b4_m49 sky130_fd_sc_hd__xor2_1
XFILLER_185_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_87_0 c$3740 c$3742 s$3745 VGND VGND VPWR VPWR c$4070 s$4071 sky130_fd_sc_hd__fa_2
XFILLER_172_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_101_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_101_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_5_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0410_ clknet_leaf_197_clk net230 VGND VGND VPWR VPWR pp_row76_28 sky130_fd_sc_hd__dfxtp_1
X_1390_ clknet_leaf_5_clk net1430 VGND VGND VPWR VPWR pp_row32_17 sky130_fd_sc_hd__dfxtp_1
X_0341_ clknet_leaf_202_clk booth_b56_m18 VGND VGND VPWR VPWR pp_row74_24 sky130_fd_sc_hd__dfxtp_1
XFILLER_171_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0272_ clknet_leaf_217_clk booth_b50_m22 VGND VGND VPWR VPWR pp_row72_22 sky130_fd_sc_hd__dfxtp_1
X_2011_ clknet_leaf_231_clk net207 VGND VGND VPWR VPWR pp_row55_28 sky130_fd_sc_hd__dfxtp_4
Xclkbuf_leaf_168_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_168_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$880 net1074 net396 net1066 net662 VGND VGND VPWR VPWR t$4855 sky130_fd_sc_hd__a22o_1
XFILLER_23_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1030 t$4931 net1184 VGND VGND VPWR VPWR booth_b14_m32 sky130_fd_sc_hd__xor2_1
XU$$891 t$4860 net1311 VGND VGND VPWR VPWR booth_b12_m31 sky130_fd_sc_hd__xor2_1
XU$$1041 net961 net388 net955 net654 VGND VGND VPWR VPWR t$4937 sky130_fd_sc_hd__a22o_1
XU$$1052 t$4942 net1187 VGND VGND VPWR VPWR booth_b14_m43 sky130_fd_sc_hd__xor2_1
XFILLER_177_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1063 net1687 net390 net1679 net656 VGND VGND VPWR VPWR t$4948 sky130_fd_sc_hd__a22o_1
XU$$1074 t$4953 net1191 VGND VGND VPWR VPWR booth_b14_m54 sky130_fd_sc_hd__xor2_1
XU$$1085 net1578 net391 net1551 net657 VGND VGND VPWR VPWR t$4959 sky130_fd_sc_hd__a22o_1
XU$$1096 net1188 VGND VGND VPWR VPWR notblock$4965\[0\] sky130_fd_sc_hd__inv_1
XFILLER_148_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1726_ clknet_leaf_23_clk booth_b36_m10 VGND VGND VPWR VPWR pp_row46_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_137_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1657_ clknet_leaf_6_clk booth_b8_m36 VGND VGND VPWR VPWR pp_row44_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_160_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4517_1879 VGND VGND VPWR VPWR U$$4517_1879/HI net1879 sky130_fd_sc_hd__conb_1
Xdadda_fa_1_81_7 pp_row81_21 pp_row81_22 pp_row81_23 VGND VGND VPWR VPWR c$920 s$921
+ sky130_fd_sc_hd__fa_1
XFILLER_176_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout604 sel_0$5247 VGND VGND VPWR VPWR net604 sky130_fd_sc_hd__buf_4
X_0608_ clknet_leaf_172_clk booth_b56_m27 VGND VGND VPWR VPWR pp_row83_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_98_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1588_ clknet_leaf_9_clk booth_b22_m19 VGND VGND VPWR VPWR pp_row41_11 sky130_fd_sc_hd__dfxtp_1
Xfanout615 sel_0$5177 VGND VGND VPWR VPWR net615 sky130_fd_sc_hd__buf_4
Xfanout626 sel_0$4477 VGND VGND VPWR VPWR net626 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_74_6 pp_row74_26 pp_row74_27 pp_row74_28 VGND VGND VPWR VPWR c$792 s$793
+ sky130_fd_sc_hd__fa_1
XFILLER_101_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout637 net638 VGND VGND VPWR VPWR net637 sky130_fd_sc_hd__buf_4
XFILLER_99_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout648 net650 VGND VGND VPWR VPWR net648 sky130_fd_sc_hd__buf_6
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0539_ clknet_leaf_163_clk booth_b30_m51 VGND VGND VPWR VPWR pp_row81_7 sky130_fd_sc_hd__dfxtp_1
Xfanout659 net660 VGND VGND VPWR VPWR net659 sky130_fd_sc_hd__buf_4
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_67_5 pp_row67_33 c$108 c$110 VGND VGND VPWR VPWR c$664 s$665 sky130_fd_sc_hd__fa_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_159_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_159_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2209_ clknet_leaf_212_clk booth_b40_m21 VGND VGND VPWR VPWR pp_row61_20 sky130_fd_sc_hd__dfxtp_1
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_1051 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_62_4 pp_row62_12 pp_row62_13 pp_row62_14 VGND VGND VPWR VPWR c$68 s$69
+ sky130_fd_sc_hd__fa_1
XFILLER_76_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3905 t$6400 net1292 VGND VGND VPWR VPWR booth_b56_m31 sky130_fd_sc_hd__xor2_1
XTAP_4254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3916 net970 net462 net962 net735 VGND VGND VPWR VPWR t$6406 sky130_fd_sc_hd__a22o_1
Xdadda_ha_3_19_2 pp_row19_6 pp_row19_7 VGND VGND VPWR VPWR c$1996 s$1997 sky130_fd_sc_hd__ha_1
XTAP_4265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3927 t$6411 net1298 VGND VGND VPWR VPWR booth_b56_m42 sky130_fd_sc_hd__xor2_1
XTAP_3531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$260 final_adder.p_new$262 final_adder.p_new$260 VGND VGND VPWR VPWR
+ final_adder.p_new$388 sky130_fd_sc_hd__and2_1
XTAP_4276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$110 net1650 net449 net1641 net691 VGND VGND VPWR VPWR t$4462 sky130_fd_sc_hd__a22o_1
XU$$3938 net1701 net466 net1694 net739 VGND VGND VPWR VPWR t$6417 sky130_fd_sc_hd__a22o_1
XTAP_4287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3949 t$6422 net1293 VGND VGND VPWR VPWR booth_b56_m53 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$271 final_adder.p_new$270 final_adder.g_new$273 final_adder.g_new$271
+ VGND VGND VPWR VPWR final_adder.g_new$399 sky130_fd_sc_hd__a21o_1
XTAP_4298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$282 final_adder.p_new$284 final_adder.p_new$282 VGND VGND VPWR VPWR
+ final_adder.p_new$410 sky130_fd_sc_hd__and2_1
Xdadda_fa_3_32_2 c$1108 s$1111 s$1113 VGND VGND VPWR VPWR c$2098 s$2099 sky130_fd_sc_hd__fa_2
XU$$121 t$4467 net1576 VGND VGND VPWR VPWR booth_b0_m57 sky130_fd_sc_hd__xor2_1
XTAP_3564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$132 net1535 net444 net1527 net686 VGND VGND VPWR VPWR t$4473 sky130_fd_sc_hd__a22o_1
XFILLER_40_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$293 final_adder.p_new$292 final_adder.g_new$295 final_adder.g_new$293
+ VGND VGND VPWR VPWR final_adder.g_new$421 sky130_fd_sc_hd__a21o_1
XU$$143 net1761 net624 net1231 net897 VGND VGND VPWR VPWR t$4479 sky130_fd_sc_hd__a22o_1
XTAP_3575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$154 t$4484 net1390 VGND VGND VPWR VPWR booth_b2_m5 sky130_fd_sc_hd__xor2_1
XTAP_3586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_25_1 pp_row25_8 pp_row25_9 pp_row25_10 VGND VGND VPWR VPWR c$2040 s$2041
+ sky130_fd_sc_hd__fa_1
XFILLER_75_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$165 net1224 net625 net1216 net898 VGND VGND VPWR VPWR t$4490 sky130_fd_sc_hd__a22o_1
XFILLER_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$176 t$4495 net1386 VGND VGND VPWR VPWR booth_b2_m16 sky130_fd_sc_hd__xor2_1
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$187 net1106 net620 net1099 net893 VGND VGND VPWR VPWR t$4501 sky130_fd_sc_hd__a22o_1
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$198 t$4506 net1385 VGND VGND VPWR VPWR booth_b2_m27 sky130_fd_sc_hd__xor2_1
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_18_0 pp_row18_0 pp_row18_1 pp_row18_2 VGND VGND VPWR VPWR c$1986 s$1987
+ sky130_fd_sc_hd__fa_1
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_996 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0890_ clknet_leaf_100_clk booth_b46_m49 VGND VGND VPWR VPWR pp_row95_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_158_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_776 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1511_ clknet_leaf_44_clk booth_b14_m24 VGND VGND VPWR VPWR pp_row38_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_142_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2491_ clknet_leaf_125_clk booth_b56_m56 VGND VGND VPWR VPWR pp_row112_5 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_84_5 s$959 s$961 s$963 VGND VGND VPWR VPWR c$1744 s$1745 sky130_fd_sc_hd__fa_2
X_1442_ clknet_leaf_54_clk booth_b10_m25 VGND VGND VPWR VPWR pp_row35_5 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_77_4 s$839 s$841 s$843 VGND VGND VPWR VPWR c$1658 s$1659 sky130_fd_sc_hd__fa_1
X_1373_ clknet_leaf_7_clk booth_b2_m30 VGND VGND VPWR VPWR pp_row32_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_68_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0324_ clknet_leaf_199_clk booth_b24_m50 VGND VGND VPWR VPWR pp_row74_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_96_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0255_ clknet_leaf_124_clk booth_b54_m59 VGND VGND VPWR VPWR pp_row113_3 sky130_fd_sc_hd__dfxtp_1
X_0186_ clknet_leaf_148_clk booth_b16_m54 VGND VGND VPWR VPWR pp_row70_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_63_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_100_3 pp_row100_9 pp_row100_10 pp_row100_11 VGND VGND VPWR VPWR c$1930
+ s$1931 sky130_fd_sc_hd__fa_1
XFILLER_51_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1082 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_114_1 s$3375 s$3377 s$3379 VGND VGND VPWR VPWR c$3854 s$3855 sky130_fd_sc_hd__fa_1
XFILLER_191_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_107_0 c$3326 c$3328 c$3330 VGND VGND VPWR VPWR c$3824 s$3825 sky130_fd_sc_hd__fa_1
XFILLER_173_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1709_ clknet_leaf_236_clk booth_b4_m42 VGND VGND VPWR VPWR pp_row46_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_145_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout401 net402 VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__buf_4
Xfanout412 net417 VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_72_3 pp_row72_20 pp_row72_21 pp_row72_22 VGND VGND VPWR VPWR c$750 s$751
+ sky130_fd_sc_hd__fa_1
Xfanout423 net425 VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__buf_4
Xfanout434 net437 VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__buf_4
Xfanout445 net450 VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__buf_4
XFILLER_171_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout456 net458 VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_65_2 pp_row65_24 pp_row65_25 pp_row65_26 VGND VGND VPWR VPWR c$622 s$623
+ sky130_fd_sc_hd__fa_1
Xfanout467 sel_0$6367 VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__buf_6
XFILLER_59_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout478 net479 VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__buf_2
Xfanout489 net491 VGND VGND VPWR VPWR net489 sky130_fd_sc_hd__buf_4
Xdadda_fa_4_42_1 c$2170 c$2172 s$2175 VGND VGND VPWR VPWR c$2944 s$2945 sky130_fd_sc_hd__fa_1
XFILLER_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_58_1 pp_row58_14 pp_row58_15 pp_row58_16 VGND VGND VPWR VPWR c$494 s$495
+ sky130_fd_sc_hd__fa_1
Xdadda_fa_1_82_0_1897 VGND VGND VPWR VPWR net1897 dadda_fa_1_82_0_1897/LO sky130_fd_sc_hd__conb_1
Xdadda_fa_4_35_0 s$1157 c$2110 c$2112 VGND VGND VPWR VPWR c$2900 s$2901 sky130_fd_sc_hd__fa_1
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_87_3 s$1775 s$1777 s$1779 VGND VGND VPWR VPWR c$2540 s$2541 sky130_fd_sc_hd__fa_2
XFILLER_123_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4403 t$6655 net1822 VGND VGND VPWR VPWR booth_b64_m6 sky130_fd_sc_hd__xor2_1
XU$$4414 net1214 sel_0$6647 net1205 net694 VGND VGND VPWR VPWR t$6661 sky130_fd_sc_hd__a22o_1
XU$$4425 t$6666 net1833 VGND VGND VPWR VPWR booth_b64_m17 sky130_fd_sc_hd__xor2_1
Xdadda_fa_0_60_1 pp_row60_3 pp_row60_4 pp_row60_5 VGND VGND VPWR VPWR c$42 s$43 sky130_fd_sc_hd__fa_1
Xfanout990 net991 VGND VGND VPWR VPWR net990 sky130_fd_sc_hd__buf_4
XTAP_4040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4436 net1103 sel_0$6647 net1095 net693 VGND VGND VPWR VPWR t$6672 sky130_fd_sc_hd__a22o_1
XU$$4447 t$6677 net1844 VGND VGND VPWR VPWR booth_b64_m28 sky130_fd_sc_hd__xor2_1
XU$$3702 net1301 notblock$6295\[1\] VGND VGND VPWR VPWR t$6296 sky130_fd_sc_hd__and2_1
XFILLER_93_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4458 net997 sel_0$6647 net989 net697 VGND VGND VPWR VPWR t$6683 sky130_fd_sc_hd__a22o_1
XFILLER_64_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3713 net938 net472 net1677 net745 VGND VGND VPWR VPWR t$6303 sky130_fd_sc_hd__a22o_1
XTAP_4062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4469 t$6688 net1855 VGND VGND VPWR VPWR booth_b64_m39 sky130_fd_sc_hd__xor2_1
XU$$3724 t$6308 net1300 VGND VGND VPWR VPWR booth_b54_m9 sky130_fd_sc_hd__xor2_1
XTAP_4073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3735 net1182 net475 net1172 net748 VGND VGND VPWR VPWR t$6314 sky130_fd_sc_hd__a22o_1
XTAP_4084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3746 t$6319 net1300 VGND VGND VPWR VPWR booth_b54_m20 sky130_fd_sc_hd__xor2_1
XTAP_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3757 net1077 net469 net1068 net742 VGND VGND VPWR VPWR t$6325 sky130_fd_sc_hd__a22o_1
XU$$3768 t$6330 net1303 VGND VGND VPWR VPWR booth_b54_m31 sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_109_2 s$2713 s$2715 s$2717 VGND VGND VPWR VPWR c$3348 s$3349 sky130_fd_sc_hd__fa_1
XTAP_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3779 net970 net472 net962 net745 VGND VGND VPWR VPWR t$6336 sky130_fd_sc_hd__a22o_1
XTAP_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_350 net888 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_361 net1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_372 net1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_383 net1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_394 net1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1991_ clknet_leaf_81_clk booth_b20_m35 VGND VGND VPWR VPWR pp_row55_10 sky130_fd_sc_hd__dfxtp_1
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0942_ clknet_leaf_113_clk booth_b36_m62 VGND VGND VPWR VPWR pp_row98_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_158_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0873_ clknet_leaf_141_clk booth_b54_m40 VGND VGND VPWR VPWR pp_row94_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_146_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_82_2 c$912 c$914 c$916 VGND VGND VPWR VPWR c$1714 s$1715 sky130_fd_sc_hd__fa_1
XFILLER_142_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2474_ clknet_leaf_99_clk booth_b56_m12 VGND VGND VPWR VPWR pp_row68_27 sky130_fd_sc_hd__dfxtp_1
XFILLER_87_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_75_1 c$784 c$786 c$788 VGND VGND VPWR VPWR c$1628 s$1629 sky130_fd_sc_hd__fa_1
XFILLER_141_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1425_ clknet_leaf_56_clk booth_b20_m14 VGND VGND VPWR VPWR pp_row34_10 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_52_0 c$2996 c$2998 c$3000 VGND VGND VPWR VPWR c$3604 s$3605 sky130_fd_sc_hd__fa_2
XFILLER_123_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_68_0 s$143 c$654 c$656 VGND VGND VPWR VPWR c$1542 s$1543 sky130_fd_sc_hd__fa_1
X_1356_ clknet_leaf_10_clk booth_b6_m25 VGND VGND VPWR VPWR pp_row31_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_84_903 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0307_ clknet_leaf_226_clk booth_b52_m21 VGND VGND VPWR VPWR pp_row73_22 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_0_70_0_1892 VGND VGND VPWR VPWR net1892 dadda_fa_0_70_0_1892/LO sky130_fd_sc_hd__conb_1
X_1287_ clknet_leaf_1_clk booth_b12_m15 VGND VGND VPWR VPWR pp_row27_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_37_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0238_ clknet_leaf_150_clk booth_b48_m23 VGND VGND VPWR VPWR pp_row71_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_110_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0169_ clknet_leaf_97_clk booth_b46_m23 VGND VGND VPWR VPWR pp_row69_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_36_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_90_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_90_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_19_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_97_2 s$2617 s$2619 s$2621 VGND VGND VPWR VPWR c$3276 s$3277 sky130_fd_sc_hd__fa_1
XFILLER_192_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_5_30__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_5_30__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_65_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_67_0 s$3667 c$4028 s$4031 VGND VGND VPWR VPWR c$4286 s$4287 sky130_fd_sc_hd__fa_1
XFILLER_182_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1207 net1208 VGND VGND VPWR VPWR net1207 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_1_70_0 pp_row70_14 pp_row70_15 pp_row70_16 VGND VGND VPWR VPWR c$708 s$709
+ sky130_fd_sc_hd__fa_1
Xfanout1218 net67 VGND VGND VPWR VPWR net1218 sky130_fd_sc_hd__buf_6
Xfanout1229 net1234 VGND VGND VPWR VPWR net1229 sky130_fd_sc_hd__buf_4
XFILLER_132_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3009 net1542 net524 net1534 net797 VGND VGND VPWR VPWR t$5942 sky130_fd_sc_hd__a22o_1
XFILLER_59_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2308 net1622 net574 net1613 net847 VGND VGND VPWR VPWR t$5584 sky130_fd_sc_hd__a22o_1
XU$$2319 t$5589 net1437 VGND VGND VPWR VPWR booth_b32_m60 sky130_fd_sc_hd__xor2_1
XFILLER_55_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1607 net1706 net618 net1698 net891 VGND VGND VPWR VPWR t$5226 sky130_fd_sc_hd__a22o_1
XFILLER_188_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1618 t$5231 net1483 VGND VGND VPWR VPWR booth_b22_m52 sky130_fd_sc_hd__xor2_1
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1629 net1597 net616 net1588 net889 VGND VGND VPWR VPWR t$5237 sky130_fd_sc_hd__a22o_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_81_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_81_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_131_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_92_1 c$1822 c$1824 c$1826 VGND VGND VPWR VPWR c$2576 s$2577 sky130_fd_sc_hd__fa_1
XFILLER_6_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_85_0 s$977 c$1734 c$1736 VGND VGND VPWR VPWR c$2518 s$2519 sky130_fd_sc_hd__fa_1
XFILLER_97_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1730 net1732 VGND VGND VPWR VPWR net1730 sky130_fd_sc_hd__clkbuf_4
X_1210_ clknet_leaf_49_clk booth_b18_m4 VGND VGND VPWR VPWR pp_row22_9 sky130_fd_sc_hd__dfxtp_1
Xfanout1741 net1744 VGND VGND VPWR VPWR net1741 sky130_fd_sc_hd__buf_6
X_2190_ clknet_leaf_223_clk booth_b6_m55 VGND VGND VPWR VPWR pp_row61_3 sky130_fd_sc_hd__dfxtp_1
Xfanout1752 net100 VGND VGND VPWR VPWR net1752 sky130_fd_sc_hd__buf_12
XU$$4200 net1750 net440 net1743 net722 VGND VGND VPWR VPWR t$6551 sky130_fd_sc_hd__a22o_1
XFILLER_66_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4211 t$6556 net1270 VGND VGND VPWR VPWR booth_b60_m47 sky130_fd_sc_hd__xor2_1
XU$$4222 net1643 net439 net1634 net721 VGND VGND VPWR VPWR t$6562 sky130_fd_sc_hd__a22o_1
XFILLER_65_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1141_ clknet_leaf_11_clk booth_b10_m7 VGND VGND VPWR VPWR pp_row17_5 sky130_fd_sc_hd__dfxtp_1
XU$$4233 t$6567 net1265 VGND VGND VPWR VPWR booth_b60_m58 sky130_fd_sc_hd__xor2_1
XU$$4244 net1529 net435 net1807 net717 VGND VGND VPWR VPWR t$6573 sky130_fd_sc_hd__a22o_1
XU$$3510 t$6198 net1330 VGND VGND VPWR VPWR booth_b50_m39 sky130_fd_sc_hd__xor2_1
XFILLER_92_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_47_5 s$309 s$311 s$313 VGND VGND VPWR VPWR c$1300 s$1301 sky130_fd_sc_hd__fa_2
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4255 net1234 net421 net1125 net703 VGND VGND VPWR VPWR t$6580 sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_114_0 pp_row114_5 pp_row114_6 pp_row114_7 VGND VGND VPWR VPWR c$3374 s$3375
+ sky130_fd_sc_hd__fa_1
XU$$4266 t$6585 net1259 VGND VGND VPWR VPWR booth_b62_m6 sky130_fd_sc_hd__xor2_1
XU$$3521 net1725 net492 net1715 net765 VGND VGND VPWR VPWR t$6204 sky130_fd_sc_hd__a22o_1
XU$$3532 t$6209 net1335 VGND VGND VPWR VPWR booth_b50_m50 sky130_fd_sc_hd__xor2_1
XFILLER_168_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4277 net1214 net418 net1205 net700 VGND VGND VPWR VPWR t$6591 sky130_fd_sc_hd__a22o_1
X_1072_ clknet_leaf_120_clk booth_b50_m52 VGND VGND VPWR VPWR pp_row102_7 sky130_fd_sc_hd__dfxtp_1
XU$$4288 t$6596 net1254 VGND VGND VPWR VPWR booth_b62_m17 sky130_fd_sc_hd__xor2_1
XFILLER_81_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3543 net1616 net489 net1608 net762 VGND VGND VPWR VPWR t$6215 sky130_fd_sc_hd__a22o_1
XFILLER_168_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3554 t$6220 net1334 VGND VGND VPWR VPWR booth_b50_m61 sky130_fd_sc_hd__xor2_1
XU$$4299 net1103 net419 net1095 net701 VGND VGND VPWR VPWR t$6602 sky130_fd_sc_hd__a22o_1
XU$$2820 net967 net537 net958 net810 VGND VGND VPWR VPWR t$5846 sky130_fd_sc_hd__a22o_1
XU$$3565 net1321 notblock$6225\[1\] VGND VGND VPWR VPWR t$6226 sky130_fd_sc_hd__and2_1
XU$$2831 t$5851 net1378 VGND VGND VPWR VPWR booth_b40_m42 sky130_fd_sc_hd__xor2_1
XFILLER_74_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3576 net938 net481 net1677 net754 VGND VGND VPWR VPWR t$6233 sky130_fd_sc_hd__a22o_1
XTAP_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3587 t$6238 net1319 VGND VGND VPWR VPWR booth_b52_m9 sky130_fd_sc_hd__xor2_1
XU$$2842 net1702 net538 net1692 net811 VGND VGND VPWR VPWR t$5857 sky130_fd_sc_hd__a22o_1
XU$$3598 net1181 net480 net1172 net753 VGND VGND VPWR VPWR t$6244 sky130_fd_sc_hd__a22o_1
XU$$2853 t$5862 net1382 VGND VGND VPWR VPWR booth_b40_m53 sky130_fd_sc_hd__xor2_1
XTAP_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2864 net1592 net541 net1584 net814 VGND VGND VPWR VPWR t$5868 sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_72_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_72_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_34_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2875 t$5873 net1383 VGND VGND VPWR VPWR booth_b40_m64 sky130_fd_sc_hd__xor2_1
XU$$2886 t$5880 net1367 VGND VGND VPWR VPWR booth_b42_m1 sky130_fd_sc_hd__xor2_1
XFILLER_61_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2897 net1522 net519 net1514 net792 VGND VGND VPWR VPWR t$5886 sky130_fd_sc_hd__a22o_1
XANTENNA_180 net952 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_191 net1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_1_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_1_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_18_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1974_ clknet_leaf_71_clk booth_b48_m6 VGND VGND VPWR VPWR pp_row54_24 sky130_fd_sc_hd__dfxtp_1
XFILLER_147_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0925_ clknet_leaf_112_clk booth_b38_m59 VGND VGND VPWR VPWR pp_row97_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0856_ clknet_leaf_142_clk booth_b60_m33 VGND VGND VPWR VPWR pp_row93_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_134_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0787_ clknet_leaf_139_clk booth_b60_m30 VGND VGND VPWR VPWR pp_row90_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_170_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2457_ clknet_leaf_145_clk booth_b26_m42 VGND VGND VPWR VPWR pp_row68_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_102_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1408_ clknet_leaf_57_clk booth_b24_m9 VGND VGND VPWR VPWR pp_row33_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_152_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2388_ clknet_leaf_77_clk booth_b34_m32 VGND VGND VPWR VPWR pp_row66_17 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$815 final_adder.p_new$830 final_adder.g_new$863 final_adder.g_new$831
+ VGND VGND VPWR VPWR final_adder.g_new$943 sky130_fd_sc_hd__a21o_1
XFILLER_21_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$837 final_adder.p_new$868 final_adder.g_new$933 final_adder.g_new$869
+ VGND VGND VPWR VPWR final_adder.g_new$965 sky130_fd_sc_hd__a21o_2
X_1339_ clknet_leaf_0_clk booth_b10_m20 VGND VGND VPWR VPWR pp_row30_5 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$859 final_adder.p_new$890 final_adder.g_new$955 final_adder.g_new$891
+ VGND VGND VPWR VPWR final_adder.g_new$987 sky130_fd_sc_hd__a21o_2
XU$$709 net1508 net404 net1499 net670 VGND VGND VPWR VPWR t$4768 sky130_fd_sc_hd__a22o_1
XFILLER_83_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_63_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_63_clk sky130_fd_sc_hd__clkbuf_16
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_109_1 pp_row109_3 pp_row109_4 pp_row109_5 VGND VGND VPWR VPWR c$2712 s$2713
+ sky130_fd_sc_hd__fa_1
XFILLER_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1004 net1005 VGND VGND VPWR VPWR net1004 sky130_fd_sc_hd__buf_6
Xfanout1015 net1016 VGND VGND VPWR VPWR net1015 sky130_fd_sc_hd__buf_4
XFILLER_126_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1026 net1030 VGND VGND VPWR VPWR net1026 sky130_fd_sc_hd__buf_6
XFILLER_121_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1037 net1038 VGND VGND VPWR VPWR net1037 sky130_fd_sc_hd__buf_4
Xfanout1048 net1054 VGND VGND VPWR VPWR net1048 sky130_fd_sc_hd__buf_6
Xfanout1059 net84 VGND VGND VPWR VPWR net1059 sky130_fd_sc_hd__buf_4
XFILLER_48_947 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2105 net1108 net580 net1100 net853 VGND VGND VPWR VPWR t$5481 sky130_fd_sc_hd__a22o_1
XU$$2116 t$5486 net1441 VGND VGND VPWR VPWR booth_b30_m27 sky130_fd_sc_hd__xor2_1
XU$$2127 net999 net579 net991 net852 VGND VGND VPWR VPWR t$5492 sky130_fd_sc_hd__a22o_1
XU$$2138 t$5497 net1446 VGND VGND VPWR VPWR booth_b30_m38 sky130_fd_sc_hd__xor2_1
XU$$2149 net1729 net576 net1720 net849 VGND VGND VPWR VPWR t$5503 sky130_fd_sc_hd__a22o_1
XU$$1404 net1198 net629 net1179 net902 VGND VGND VPWR VPWR t$5123 sky130_fd_sc_hd__a22o_1
XFILLER_27_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1415 t$5128 net1486 VGND VGND VPWR VPWR booth_b20_m19 sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_54_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_54_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_167_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1426 net1081 net628 net1072 net901 VGND VGND VPWR VPWR t$5134 sky130_fd_sc_hd__a22o_1
XFILLER_37_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1437 t$5139 net1487 VGND VGND VPWR VPWR booth_b20_m30 sky130_fd_sc_hd__xor2_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1448 net977 net630 net969 net903 VGND VGND VPWR VPWR t$5145 sky130_fd_sc_hd__a22o_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1459 t$5150 net1490 VGND VGND VPWR VPWR booth_b20_m41 sky130_fd_sc_hd__xor2_1
XFILLER_163_1035 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0710_ clknet_leaf_132_clk booth_b54_m64 VGND VGND VPWR VPWR pp_row118_1 sky130_fd_sc_hd__dfxtp_1
X_1690_ clknet_leaf_19_clk booth_b18_m27 VGND VGND VPWR VPWR pp_row45_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_167_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0641_ clknet_leaf_185_clk net239 VGND VGND VPWR VPWR pp_row84_24 sky130_fd_sc_hd__dfxtp_1
XFILLER_7_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0572_ clknet_leaf_189_clk booth_b40_m42 VGND VGND VPWR VPWR pp_row82_12 sky130_fd_sc_hd__dfxtp_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2311_ clknet_leaf_85_clk booth_b26_m38 VGND VGND VPWR VPWR pp_row64_13 sky130_fd_sc_hd__dfxtp_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2242_ clknet_leaf_150_clk booth_b36_m26 VGND VGND VPWR VPWR pp_row62_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_100_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1560 net1562 VGND VGND VPWR VPWR net1560 sky130_fd_sc_hd__clkbuf_4
XFILLER_78_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_52_3 c$382 s$385 s$387 VGND VGND VPWR VPWR c$1356 s$1357 sky130_fd_sc_hd__fa_2
Xfanout1571 net1572 VGND VGND VPWR VPWR net1571 sky130_fd_sc_hd__buf_2
X_2173_ clknet_leaf_224_clk booth_b40_m20 VGND VGND VPWR VPWR pp_row60_20 sky130_fd_sc_hd__dfxtp_1
Xfanout1582 net1585 VGND VGND VPWR VPWR net1582 sky130_fd_sc_hd__clkbuf_8
XU$$4030 t$6464 net1286 VGND VGND VPWR VPWR booth_b58_m25 sky130_fd_sc_hd__xor2_1
XFILLER_66_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1593 net1594 VGND VGND VPWR VPWR net1593 sky130_fd_sc_hd__buf_4
XU$$4041 net1028 net453 net1020 net726 VGND VGND VPWR VPWR t$6470 sky130_fd_sc_hd__a22o_1
XFILLER_38_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4052 t$6475 net1287 VGND VGND VPWR VPWR booth_b58_m36 sky130_fd_sc_hd__xor2_1
XU$$4063 net1750 net457 net1742 net730 VGND VGND VPWR VPWR t$6481 sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_45_2 pp_row45_23 c$264 c$266 VGND VGND VPWR VPWR c$1270 s$1271 sky130_fd_sc_hd__fa_1
X_1124_ clknet_leaf_11_clk booth_b2_m14 VGND VGND VPWR VPWR pp_row16_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_81_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4074 t$6486 net1289 VGND VGND VPWR VPWR booth_b58_m47 sky130_fd_sc_hd__xor2_1
XU$$3340 net1102 net496 net1094 net769 VGND VGND VPWR VPWR t$6112 sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_22_1 s$2823 s$2825 s$2827 VGND VGND VPWR VPWR c$3486 s$3487 sky130_fd_sc_hd__fa_1
XU$$4085 net1643 net456 net1634 net729 VGND VGND VPWR VPWR t$6492 sky130_fd_sc_hd__a22o_1
XU$$3351 t$6117 net1341 VGND VGND VPWR VPWR booth_b48_m28 sky130_fd_sc_hd__xor2_1
XU$$4096 t$6497 net1288 VGND VGND VPWR VPWR booth_b58_m58 sky130_fd_sc_hd__xor2_1
XFILLER_0_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3362 net994 net494 net984 net767 VGND VGND VPWR VPWR t$6123 sky130_fd_sc_hd__a22o_1
XFILLER_47_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_38_1 pp_row38_11 pp_row38_12 pp_row38_13 VGND VGND VPWR VPWR c$1184 s$1185
+ sky130_fd_sc_hd__fa_1
X_1055_ clknet_leaf_58_clk booth_b6_m2 VGND VGND VPWR VPWR pp_row8_3 sky130_fd_sc_hd__dfxtp_1
XU$$3373 t$6128 net1341 VGND VGND VPWR VPWR booth_b48_m39 sky130_fd_sc_hd__xor2_1
XU$$3384 net1726 net498 net1717 net771 VGND VGND VPWR VPWR t$6134 sky130_fd_sc_hd__a22o_1
XFILLER_0_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_15_0 c$2774 c$2776 c$2778 VGND VGND VPWR VPWR c$3456 s$3457 sky130_fd_sc_hd__fa_1
Xclkbuf_leaf_45_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_45_clk sky130_fd_sc_hd__clkbuf_16
XU$$3395 t$6139 net1344 VGND VGND VPWR VPWR booth_b48_m50 sky130_fd_sc_hd__xor2_1
XU$$2650 t$5759 net1402 VGND VGND VPWR VPWR booth_b38_m20 sky130_fd_sc_hd__xor2_1
XFILLER_179_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2661 net1075 net549 net1067 net822 VGND VGND VPWR VPWR t$5765 sky130_fd_sc_hd__a22o_1
XFILLER_34_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2672 t$5770 net1400 VGND VGND VPWR VPWR booth_b38_m31 sky130_fd_sc_hd__xor2_1
XU$$2683 net966 net545 net959 net818 VGND VGND VPWR VPWR t$5776 sky130_fd_sc_hd__a22o_1
XU$$2694 t$5781 net1397 VGND VGND VPWR VPWR booth_b38_m42 sky130_fd_sc_hd__xor2_1
XU$$1960 net1148 net585 net1138 net858 VGND VGND VPWR VPWR t$5407 sky130_fd_sc_hd__a22o_1
XFILLER_181_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1971 t$5412 net1451 VGND VGND VPWR VPWR booth_b28_m23 sky130_fd_sc_hd__xor2_1
XFILLER_61_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1982 net1049 net587 net1041 net860 VGND VGND VPWR VPWR t$5418 sky130_fd_sc_hd__a22o_1
XFILLER_166_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1993 t$5423 net1450 VGND VGND VPWR VPWR booth_b28_m34 sky130_fd_sc_hd__xor2_1
XFILLER_193_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1957_ clknet_leaf_66_clk booth_b18_m36 VGND VGND VPWR VPWR pp_row54_9 sky130_fd_sc_hd__dfxtp_1
X_0908_ clknet_leaf_103_clk booth_b44_m52 VGND VGND VPWR VPWR pp_row96_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_174_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1888_ clknet_leaf_39_clk booth_b8_m44 VGND VGND VPWR VPWR pp_row52_4 sky130_fd_sc_hd__dfxtp_1
X_0839_ clknet_leaf_105_clk booth_b30_m63 VGND VGND VPWR VPWR pp_row93_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_116_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_719 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput107 b[48] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__buf_6
Xdadda_ha_1_41_3 pp_row41_9 pp_row41_10 VGND VGND VPWR VPWR c$242 s$243 sky130_fd_sc_hd__ha_1
Xinput118 b[58] VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput129 c[0] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_1
Xfinal_adder.U$$601 final_adder.p_new$604 final_adder.g_new$613 final_adder.g_new$605
+ VGND VGND VPWR VPWR final_adder.g_new$729 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$612 final_adder.p_new$624 final_adder.p_new$616 VGND VGND VPWR VPWR
+ final_adder.p_new$740 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$623 final_adder.p_new$626 final_adder.g_new$509 final_adder.g_new$627
+ VGND VGND VPWR VPWR final_adder.g_new$751 sky130_fd_sc_hd__a21o_4
XTAP_3905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$634 final_adder.p_new$658 final_adder.p_new$642 VGND VGND VPWR VPWR
+ final_adder.p_new$762 sky130_fd_sc_hd__and2_1
Xdadda_ha_4_11_1 pp_row11_3 pp_row11_4 VGND VGND VPWR VPWR c$2760 s$2761 sky130_fd_sc_hd__ha_1
XTAP_3916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$645 final_adder.p_new$652 final_adder.g_new$669 final_adder.g_new$653
+ VGND VGND VPWR VPWR final_adder.g_new$773 sky130_fd_sc_hd__a21o_1
XTAP_3927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$656 final_adder.p_new$680 final_adder.p_new$664 VGND VGND VPWR VPWR
+ final_adder.p_new$784 sky130_fd_sc_hd__and2_1
XTAP_3938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$667 final_adder.p_new$674 final_adder.g_new$691 final_adder.g_new$675
+ VGND VGND VPWR VPWR final_adder.g_new$795 sky130_fd_sc_hd__a21o_1
XU$$506 t$4663 net1246 VGND VGND VPWR VPWR booth_b6_m44 sky130_fd_sc_hd__xor2_1
XTAP_3949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$517 net1682 net432 net1657 net714 VGND VGND VPWR VPWR t$4669 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$678 final_adder.p_new$702 final_adder.p_new$686 VGND VGND VPWR VPWR
+ final_adder.p_new$806 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$689 final_adder.p_new$696 final_adder.g_new$713 final_adder.g_new$697
+ VGND VGND VPWR VPWR final_adder.g_new$817 sky130_fd_sc_hd__a21o_1
XU$$528 t$4674 net1246 VGND VGND VPWR VPWR booth_b6_m55 sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_40_1 pp_row40_3 pp_row40_4 pp_row40_5 VGND VGND VPWR VPWR c$230 s$231
+ sky130_fd_sc_hd__fa_1
XU$$539 net1559 net432 net122 net714 VGND VGND VPWR VPWR t$4680 sky130_fd_sc_hd__a22o_1
XFILLER_56_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_36_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_71_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_80 net487 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_91 net530 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_62_2 c$1468 s$1471 s$1473 VGND VGND VPWR VPWR c$2338 s$2339 sky130_fd_sc_hd__fa_1
XFILLER_122_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_1031 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_55_1 c$1378 c$1380 c$1382 VGND VGND VPWR VPWR c$2280 s$2281 sky130_fd_sc_hd__fa_1
XFILLER_94_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_32_0 c$3520 c$3522 s$3525 VGND VGND VPWR VPWR c$3960 s$3961 sky130_fd_sc_hd__fa_2
XFILLER_48_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_48_0 s$331 c$1290 c$1292 VGND VGND VPWR VPWR c$2222 s$2223 sky130_fd_sc_hd__fa_1
XFILLER_130_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_27_clk clknet_5_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_16
XU$$1201 t$5018 net1014 VGND VGND VPWR VPWR booth_b16_m49 sky130_fd_sc_hd__xor2_1
XU$$1212 net1620 net649 net1612 net922 VGND VGND VPWR VPWR t$5024 sky130_fd_sc_hd__a22o_1
XFILLER_189_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1223 t$5029 net1012 VGND VGND VPWR VPWR booth_b16_m60 sky130_fd_sc_hd__xor2_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1234 net10 VGND VGND VPWR VPWR notblock$5035\[1\] sky130_fd_sc_hd__inv_1
XFILLER_62_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1245 net1036 net638 net936 net911 VGND VGND VPWR VPWR t$5042 sky130_fd_sc_hd__a22o_1
XU$$1256 t$5047 net1662 VGND VGND VPWR VPWR booth_b18_m8 sky130_fd_sc_hd__xor2_1
XFILLER_189_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1267 net1195 net637 net1175 net910 VGND VGND VPWR VPWR t$5053 sky130_fd_sc_hd__a22o_1
XU$$1278 t$5058 net1664 VGND VGND VPWR VPWR booth_b18_m19 sky130_fd_sc_hd__xor2_1
XU$$1289 net1081 net636 net1072 net909 VGND VGND VPWR VPWR t$5064 sky130_fd_sc_hd__a22o_1
XFILLER_30_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1811_ clknet_leaf_26_clk booth_b32_m17 VGND VGND VPWR VPWR pp_row49_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_31_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_105_0 s$3819 c$4104 s$4107 VGND VGND VPWR VPWR c$4362 s$4363 sky130_fd_sc_hd__fa_1
X_1742_ clknet_leaf_237_clk booth_b10_m37 VGND VGND VPWR VPWR pp_row47_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_117_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1050 final_adder.$signal$1179 final_adder.g_new$1045 VGND VGND VPWR
+ VPWR net372 sky130_fd_sc_hd__xor2_2
XFILLER_183_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1061 final_adder.$signal$1190 final_adder.g_new$991 VGND VGND VPWR
+ VPWR net258 sky130_fd_sc_hd__xor2_1
XFILLER_7_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1673_ clknet_leaf_4_clk booth_b36_m8 VGND VGND VPWR VPWR pp_row44_18 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$1072 final_adder.$signal$1201 final_adder.g_new$1034 VGND VGND VPWR
+ VPWR net270 sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$1083 final_adder.$signal$1212 final_adder.g_new$969 VGND VGND VPWR
+ VPWR net282 sky130_fd_sc_hd__xor2_2
X_0624_ clknet_leaf_187_clk booth_b34_m50 VGND VGND VPWR VPWR pp_row84_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_113_900 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout808 net809 VGND VGND VPWR VPWR net808 sky130_fd_sc_hd__buf_4
XFILLER_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout819 net823 VGND VGND VPWR VPWR net819 sky130_fd_sc_hd__buf_6
X_0555_ clknet_leaf_126_clk booth_b56_m60 VGND VGND VPWR VPWR pp_row116_3 sky130_fd_sc_hd__dfxtp_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0486_ clknet_leaf_205_clk booth_b40_m39 VGND VGND VPWR VPWR pp_row79_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_98_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2225_ clknet_leaf_227_clk booth_b6_m56 VGND VGND VPWR VPWR pp_row62_3 sky130_fd_sc_hd__dfxtp_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_50_0 pp_row50_26 pp_row50_27 c$332 VGND VGND VPWR VPWR c$1326 s$1327 sky130_fd_sc_hd__fa_1
XFILLER_38_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1390 net1391 VGND VGND VPWR VPWR net1390 sky130_fd_sc_hd__clkbuf_8
X_2156_ clknet_leaf_215_clk booth_b12_m48 VGND VGND VPWR VPWR pp_row60_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1107_ clknet_leaf_14_clk booth_b8_m6 VGND VGND VPWR VPWR pp_row14_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3170 t$6025 net1353 VGND VGND VPWR VPWR booth_b46_m6 sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_18_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_16
X_2087_ clknet_leaf_37_clk booth_b12_m46 VGND VGND VPWR VPWR pp_row58_6 sky130_fd_sc_hd__dfxtp_1
XU$$3181 net1212 net502 net1204 net775 VGND VGND VPWR VPWR t$6031 sky130_fd_sc_hd__a22o_1
XU$$3192 t$6036 net1349 VGND VGND VPWR VPWR booth_b46_m17 sky130_fd_sc_hd__xor2_1
X_1038_ clknet_leaf_120_clk booth_b44_m58 VGND VGND VPWR VPWR pp_row102_4 sky130_fd_sc_hd__dfxtp_1
XU$$2480 net933 net552 net1672 net825 VGND VGND VPWR VPWR t$5673 sky130_fd_sc_hd__a22o_1
XU$$2491 t$5678 net1403 VGND VGND VPWR VPWR booth_b36_m9 sky130_fd_sc_hd__xor2_1
XU$$1790 t$5320 net1457 VGND VGND VPWR VPWR booth_b26_m1 sky130_fd_sc_hd__xor2_1
XFILLER_50_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_72_1 c$2410 c$2412 s$2415 VGND VGND VPWR VPWR c$3124 s$3125 sky130_fd_sc_hd__fa_1
Xdadda_fa_1_88_1 pp_row88_3 pp_row88_4 pp_row88_5 VGND VGND VPWR VPWR c$1002 s$1003
+ sky130_fd_sc_hd__fa_1
XFILLER_192_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_65_0 s$1517 c$2350 c$2352 VGND VGND VPWR VPWR c$3080 s$3081 sky130_fd_sc_hd__fa_1
XFILLER_67_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$420 final_adder.p_new$426 final_adder.p_new$422 VGND VGND VPWR VPWR
+ final_adder.p_new$548 sky130_fd_sc_hd__and2_1
XTAP_3702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$431 final_adder.p_new$432 final_adder.g_new$437 final_adder.g_new$433
+ VGND VGND VPWR VPWR final_adder.g_new$559 sky130_fd_sc_hd__a21o_1
XTAP_3713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$442 final_adder.p_new$448 final_adder.p_new$444 VGND VGND VPWR VPWR
+ final_adder.p_new$570 sky130_fd_sc_hd__and2_1
XTAP_3724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$453 final_adder.p_new$454 final_adder.g_new$459 final_adder.g_new$455
+ VGND VGND VPWR VPWR final_adder.g_new$581 sky130_fd_sc_hd__a21o_1
XTAP_3735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$303 t$4560 net1279 VGND VGND VPWR VPWR booth_b4_m11 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$464 final_adder.p_new$470 final_adder.p_new$466 VGND VGND VPWR VPWR
+ final_adder.p_new$592 sky130_fd_sc_hd__and2_1
XFILLER_177_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$314 net1161 net532 net1149 net805 VGND VGND VPWR VPWR t$4566 sky130_fd_sc_hd__a22o_1
XFILLER_123_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$475 final_adder.p_new$476 final_adder.g_new$481 final_adder.g_new$477
+ VGND VGND VPWR VPWR final_adder.g_new$603 sky130_fd_sc_hd__a21o_1
XTAP_3757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$325 t$4571 net1273 VGND VGND VPWR VPWR booth_b4_m22 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$486 final_adder.p_new$492 final_adder.p_new$488 VGND VGND VPWR VPWR
+ final_adder.p_new$614 sky130_fd_sc_hd__and2_1
XTAP_3768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$336 net1056 net528 net1048 net801 VGND VGND VPWR VPWR t$4577 sky130_fd_sc_hd__a22o_1
XFILLER_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$497 final_adder.p_new$498 final_adder.g_new$503 final_adder.g_new$499
+ VGND VGND VPWR VPWR final_adder.g_new$625 sky130_fd_sc_hd__a21o_1
XTAP_3779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$347 t$4582 net1273 VGND VGND VPWR VPWR booth_b4_m33 sky130_fd_sc_hd__xor2_1
XFILLER_17_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$358 net948 net529 net940 net802 VGND VGND VPWR VPWR t$4588 sky130_fd_sc_hd__a22o_1
XU$$369 t$4593 net1274 VGND VGND VPWR VPWR booth_b4_m44 sky130_fd_sc_hd__xor2_1
XFILLER_26_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0340_ clknet_leaf_202_clk booth_b54_m20 VGND VGND VPWR VPWR pp_row74_23 sky130_fd_sc_hd__dfxtp_1
XFILLER_110_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0271_ clknet_leaf_217_clk booth_b48_m24 VGND VGND VPWR VPWR pp_row72_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_76_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2010_ clknet_leaf_75_clk booth_b54_m1 VGND VGND VPWR VPWR pp_row55_27 sky130_fd_sc_hd__dfxtp_1
XFILLER_48_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$828_1887 VGND VGND VPWR VPWR U$$828_1887/HI net1887 sky130_fd_sc_hd__conb_1
XFILLER_36_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$870 net1117 net397 net1108 net663 VGND VGND VPWR VPWR t$4850 sky130_fd_sc_hd__a22o_1
XU$$1020 t$4926 net1184 VGND VGND VPWR VPWR booth_b14_m27 sky130_fd_sc_hd__xor2_1
XU$$881 t$4855 net1312 VGND VGND VPWR VPWR booth_b12_m26 sky130_fd_sc_hd__xor2_1
XFILLER_189_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1031 net998 net386 net990 net652 VGND VGND VPWR VPWR t$4932 sky130_fd_sc_hd__a22o_1
XU$$892 net1016 net394 net999 net660 VGND VGND VPWR VPWR t$4861 sky130_fd_sc_hd__a22o_1
XU$$1042 t$4937 net1186 VGND VGND VPWR VPWR booth_b14_m38 sky130_fd_sc_hd__xor2_1
XU$$1053 net1733 net391 net1724 net657 VGND VGND VPWR VPWR t$4943 sky130_fd_sc_hd__a22o_1
XFILLER_188_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1064 t$4948 net1190 VGND VGND VPWR VPWR booth_b14_m49 sky130_fd_sc_hd__xor2_1
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1075 net1623 net391 net1615 net657 VGND VGND VPWR VPWR t$4954 sky130_fd_sc_hd__a22o_1
XU$$1086 t$4959 net1188 VGND VGND VPWR VPWR booth_b14_m60 sky130_fd_sc_hd__xor2_1
XU$$1097 net8 VGND VGND VPWR VPWR notblock$4965\[1\] sky130_fd_sc_hd__inv_1
XFILLER_149_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1725_ clknet_leaf_21_clk booth_b34_m12 VGND VGND VPWR VPWR pp_row46_17 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_82_0 c$3176 c$3178 c$3180 VGND VGND VPWR VPWR c$3724 s$3725 sky130_fd_sc_hd__fa_1
Xdadda_fa_2_98_0 net1908 pp_row98_1 pp_row98_2 VGND VGND VPWR VPWR c$1902 s$1903 sky130_fd_sc_hd__fa_1
Xclkbuf_leaf_7_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_144_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1656_ clknet_leaf_6_clk booth_b6_m38 VGND VGND VPWR VPWR pp_row44_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0607_ clknet_leaf_174_clk booth_b54_m29 VGND VGND VPWR VPWR pp_row83_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_132_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1587_ clknet_leaf_4_clk booth_b20_m21 VGND VGND VPWR VPWR pp_row41_10 sky130_fd_sc_hd__dfxtp_1
Xfanout605 net606 VGND VGND VPWR VPWR net605 sky130_fd_sc_hd__buf_4
Xfanout616 net618 VGND VGND VPWR VPWR net616 sky130_fd_sc_hd__buf_4
XFILLER_98_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout627 net628 VGND VGND VPWR VPWR net627 sky130_fd_sc_hd__buf_4
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_74_7 pp_row74_29 c$180 c$182 VGND VGND VPWR VPWR c$794 s$795 sky130_fd_sc_hd__fa_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout638 net639 VGND VGND VPWR VPWR net638 sky130_fd_sc_hd__buf_6
XFILLER_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout649 net650 VGND VGND VPWR VPWR net649 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0538_ clknet_leaf_166_clk booth_b28_m53 VGND VGND VPWR VPWR pp_row81_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_113_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_67_6 c$112 c$114 c$116 VGND VGND VPWR VPWR c$666 s$667 sky130_fd_sc_hd__fa_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0469_ clknet_leaf_155_clk booth_b62_m16 VGND VGND VPWR VPWR pp_row78_25 sky130_fd_sc_hd__dfxtp_1
XFILLER_85_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2208_ clknet_leaf_29_clk booth_b38_m23 VGND VGND VPWR VPWR pp_row61_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_160_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2139_ clknet_leaf_26_clk booth_b42_m17 VGND VGND VPWR VPWR pp_row59_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_183_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_ha_1_94_1 pp_row94_3 pp_row94_4 VGND VGND VPWR VPWR c$1044 s$1045 sky130_fd_sc_hd__ha_1
Xdadda_fa_7_97_0 s$3787 c$4088 s$4091 VGND VGND VPWR VPWR c$4346 s$4347 sky130_fd_sc_hd__fa_1
XFILLER_33_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_803 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_112_0 c$3840 c$3842 s$3845 VGND VGND VPWR VPWR c$4120 s$4121 sky130_fd_sc_hd__fa_1
XFILLER_134_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3906 net1020 net462 net1003 net735 VGND VGND VPWR VPWR t$6401 sky130_fd_sc_hd__a22o_1
XTAP_4255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3917 t$6406 net1293 VGND VGND VPWR VPWR booth_b56_m37 sky130_fd_sc_hd__xor2_1
XFILLER_131_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3928 net1742 net466 net1734 net739 VGND VGND VPWR VPWR t$6412 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$250 final_adder.$signal$1094 final_adder.$signal$1095 VGND VGND VPWR
+ VPWR final_adder.p_new$378 sky130_fd_sc_hd__and2_1
XTAP_3521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3939 t$6417 net1298 VGND VGND VPWR VPWR booth_b56_m48 sky130_fd_sc_hd__xor2_1
XU$$100 net1703 net444 net1695 net686 VGND VGND VPWR VPWR t$4457 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$261 final_adder.p_new$260 final_adder.g_new$263 final_adder.g_new$261
+ VGND VGND VPWR VPWR final_adder.g_new$389 sky130_fd_sc_hd__a21o_1
XTAP_4288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$111 t$4462 net1576 VGND VGND VPWR VPWR booth_b0_m52 sky130_fd_sc_hd__xor2_1
XTAP_3543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$272 final_adder.p_new$274 final_adder.p_new$272 VGND VGND VPWR VPWR
+ final_adder.p_new$400 sky130_fd_sc_hd__and2_1
XTAP_3554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$283 final_adder.p_new$282 final_adder.g_new$285 final_adder.g_new$283
+ VGND VGND VPWR VPWR final_adder.g_new$411 sky130_fd_sc_hd__a21o_1
XFILLER_27_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_32_3 s$1115 s$1117 s$1119 VGND VGND VPWR VPWR c$2100 s$2101 sky130_fd_sc_hd__fa_2
XU$$122 net1599 net449 net1590 net691 VGND VGND VPWR VPWR t$4468 sky130_fd_sc_hd__a22o_1
XTAP_4299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$133 t$4473 net1570 VGND VGND VPWR VPWR booth_b0_m63 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$294 final_adder.p_new$296 final_adder.p_new$294 VGND VGND VPWR VPWR
+ final_adder.p_new$422 sky130_fd_sc_hd__and2_1
XU$$144 t$4479 net1390 VGND VGND VPWR VPWR booth_b2_m0 sky130_fd_sc_hd__xor2_1
XTAP_3576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$155 net1564 net624 net1523 net897 VGND VGND VPWR VPWR t$4485 sky130_fd_sc_hd__a22o_1
XTAP_3598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$166 t$4490 net1391 VGND VGND VPWR VPWR booth_b2_m11 sky130_fd_sc_hd__xor2_1
XFILLER_33_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_25_2 pp_row25_11 pp_row25_12 pp_row25_13 VGND VGND VPWR VPWR c$2042 s$2043
+ sky130_fd_sc_hd__fa_1
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$177 net1157 net623 net1149 net896 VGND VGND VPWR VPWR t$4496 sky130_fd_sc_hd__a22o_1
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$188 t$4501 net1386 VGND VGND VPWR VPWR booth_b2_m22 sky130_fd_sc_hd__xor2_1
XU$$199 net1055 net619 net1047 net892 VGND VGND VPWR VPWR t$4507 sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_18_1 pp_row18_3 pp_row18_4 pp_row18_5 VGND VGND VPWR VPWR c$1988 s$1989
+ sky130_fd_sc_hd__fa_1
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_942 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_788 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1510_ clknet_leaf_44_clk booth_b12_m26 VGND VGND VPWR VPWR pp_row38_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_99_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2490_ clknet_leaf_90_clk booth_b22_m47 VGND VGND VPWR VPWR pp_row69_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_153_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1441_ clknet_leaf_54_clk booth_b8_m27 VGND VGND VPWR VPWR pp_row35_4 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_77_5 s$845 s$847 s$849 VGND VGND VPWR VPWR c$1660 s$1661 sky130_fd_sc_hd__fa_2
X_1372_ clknet_leaf_7_clk booth_b0_m32 VGND VGND VPWR VPWR pp_row32_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_122_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0323_ clknet_leaf_201_clk booth_b22_m52 VGND VGND VPWR VPWR pp_row74_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_110_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0254_ clknet_leaf_209_clk booth_b18_m54 VGND VGND VPWR VPWR pp_row72_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0185_ clknet_leaf_90_clk booth_b14_m56 VGND VGND VPWR VPWR pp_row70_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_107_1 s$3333 s$3335 s$3337 VGND VGND VPWR VPWR c$3826 s$3827 sky130_fd_sc_hd__fa_1
XFILLER_191_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1708_ clknet_leaf_236_clk booth_b2_m44 VGND VGND VPWR VPWR pp_row46_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_117_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1639_ clknet_leaf_184_clk net135 VGND VGND VPWR VPWR pp_row105_13 sky130_fd_sc_hd__dfxtp_2
XFILLER_133_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout402 net408 VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__buf_4
XFILLER_160_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout413 net414 VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__buf_4
XFILLER_87_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_72_4 pp_row72_23 pp_row72_24 pp_row72_25 VGND VGND VPWR VPWR c$752 s$753
+ sky130_fd_sc_hd__fa_1
Xfanout424 net425 VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__clkbuf_4
Xfanout435 net436 VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__clkbuf_4
XFILLER_115_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout446 net447 VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__clkbuf_4
Xfanout457 net458 VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__clkbuf_4
Xfanout468 net471 VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_65_3 pp_row65_27 pp_row65_28 pp_row65_29 VGND VGND VPWR VPWR c$624 s$625
+ sky130_fd_sc_hd__fa_1
XFILLER_171_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout479 sel_0$6227 VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__buf_4
XFILLER_115_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_42_2 s$2177 s$2179 s$2181 VGND VGND VPWR VPWR c$2946 s$2947 sky130_fd_sc_hd__fa_1
XFILLER_86_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_58_2 pp_row58_17 pp_row58_18 pp_row58_19 VGND VGND VPWR VPWR c$496 s$497
+ sky130_fd_sc_hd__fa_1
XFILLER_27_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_35_1 c$2114 c$2116 s$2119 VGND VGND VPWR VPWR c$2902 s$2903 sky130_fd_sc_hd__fa_1
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_12_0 s$3447 c$3918 s$3921 VGND VGND VPWR VPWR c$4176 s$4177 sky130_fd_sc_hd__fa_1
Xdadda_fa_4_28_0 s$1081 c$2054 c$2056 VGND VGND VPWR VPWR c$2858 s$2859 sky130_fd_sc_hd__fa_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_0_61_4 pp_row61_12 pp_row61_13 VGND VGND VPWR VPWR c$58 s$59 sky130_fd_sc_hd__ha_1
XFILLER_124_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4404 net125 sel_0$6647 net1518 net696 VGND VGND VPWR VPWR t$6656 sky130_fd_sc_hd__a22o_1
XU$$4415 t$6661 net1828 VGND VGND VPWR VPWR booth_b64_m12 sky130_fd_sc_hd__xor2_1
Xfanout980 net981 VGND VGND VPWR VPWR net980 sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_240_clk clknet_5_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_240_clk
+ sky130_fd_sc_hd__clkbuf_16
XU$$4426 net1152 sel_0$6647 net1141 net693 VGND VGND VPWR VPWR t$6667 sky130_fd_sc_hd__a22o_1
Xdadda_fa_0_60_2 pp_row60_6 pp_row60_7 pp_row60_8 VGND VGND VPWR VPWR c$44 s$45 sky130_fd_sc_hd__fa_1
XTAP_4030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4437 t$6672 net1839 VGND VGND VPWR VPWR booth_b64_m23 sky130_fd_sc_hd__xor2_1
Xfanout991 net91 VGND VGND VPWR VPWR net991 sky130_fd_sc_hd__buf_6
XTAP_4041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3703 notblock$6295\[2\] net50 net1321 t$6296 notblock$6295\[0\] VGND VGND VPWR
+ VPWR sel_0$6297 sky130_fd_sc_hd__a32o_2
XTAP_4052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4448 net1054 sel_0$6647 net1046 net696 VGND VGND VPWR VPWR t$6678 sky130_fd_sc_hd__a22o_1
XTAP_4063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4459 t$6683 net1850 VGND VGND VPWR VPWR booth_b64_m34 sky130_fd_sc_hd__xor2_1
XFILLER_64_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3714 t$6303 net1305 VGND VGND VPWR VPWR booth_b54_m4 sky130_fd_sc_hd__xor2_1
XU$$3725 net1501 net472 net1226 net745 VGND VGND VPWR VPWR t$6309 sky130_fd_sc_hd__a22o_1
XFILLER_46_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3736 t$6314 net1304 VGND VGND VPWR VPWR booth_b54_m15 sky130_fd_sc_hd__xor2_1
XTAP_4085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3747 net1120 net468 net1111 net741 VGND VGND VPWR VPWR t$6320 sky130_fd_sc_hd__a22o_1
XTAP_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_30_0 pp_row30_14 pp_row30_15 pp_row30_16 VGND VGND VPWR VPWR c$2078 s$2079
+ sky130_fd_sc_hd__fa_1
XU$$3758 t$6325 net1303 VGND VGND VPWR VPWR booth_b54_m26 sky130_fd_sc_hd__xor2_1
XFILLER_92_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3769 net1020 net469 net1003 net742 VGND VGND VPWR VPWR t$6331 sky130_fd_sc_hd__a22o_1
XTAP_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_340 net782 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_351 net888 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_362 net1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_373 net1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_384 net1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_395 net1546 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1990_ clknet_leaf_81_clk booth_b18_m37 VGND VGND VPWR VPWR pp_row55_9 sky130_fd_sc_hd__dfxtp_1
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0941_ clknet_leaf_113_clk booth_b34_m64 VGND VGND VPWR VPWR pp_row98_1 sky130_fd_sc_hd__dfxtp_1
XU$$4403_1822 VGND VGND VPWR VPWR U$$4403_1822/HI net1822 sky130_fd_sc_hd__conb_1
X_0872_ clknet_leaf_141_clk booth_b52_m42 VGND VGND VPWR VPWR pp_row94_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_158_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_82_3 c$918 c$920 s$923 VGND VGND VPWR VPWR c$1716 s$1717 sky130_fd_sc_hd__fa_1
X_2473_ clknet_leaf_98_clk booth_b54_m14 VGND VGND VPWR VPWR pp_row68_26 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_75_2 c$790 c$792 c$794 VGND VGND VPWR VPWR c$1630 s$1631 sky130_fd_sc_hd__fa_1
X_1424_ clknet_leaf_56_clk booth_b18_m16 VGND VGND VPWR VPWR pp_row34_9 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_52_1 s$3003 s$3005 s$3007 VGND VGND VPWR VPWR c$3606 s$3607 sky130_fd_sc_hd__fa_1
Xdadda_fa_2_68_1 c$658 c$660 c$662 VGND VGND VPWR VPWR c$1544 s$1545 sky130_fd_sc_hd__fa_2
XFILLER_110_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1355_ clknet_leaf_3_clk booth_b4_m27 VGND VGND VPWR VPWR pp_row31_2 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_45_0 c$2954 c$2956 c$2958 VGND VGND VPWR VPWR c$3576 s$3577 sky130_fd_sc_hd__fa_1
XFILLER_84_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_231_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_231_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0306_ clknet_leaf_226_clk booth_b50_m23 VGND VGND VPWR VPWR pp_row73_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_56_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1286_ clknet_leaf_1_clk booth_b10_m17 VGND VGND VPWR VPWR pp_row27_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0237_ clknet_leaf_211_clk booth_b46_m25 VGND VGND VPWR VPWR pp_row71_20 sky130_fd_sc_hd__dfxtp_1
XFILLER_92_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0168_ clknet_leaf_147_clk booth_b44_m25 VGND VGND VPWR VPWR pp_row69_20 sky130_fd_sc_hd__dfxtp_1
XFILLER_34_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1208 net1209 VGND VGND VPWR VPWR net1208 sky130_fd_sc_hd__buf_4
Xfanout1219 net1220 VGND VGND VPWR VPWR net1219 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_70_1 pp_row70_17 pp_row70_18 pp_row70_19 VGND VGND VPWR VPWR c$710 s$711
+ sky130_fd_sc_hd__fa_1
XFILLER_113_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_63_0 pp_row63_17 pp_row63_18 pp_row63_19 VGND VGND VPWR VPWR c$582 s$583
+ sky130_fd_sc_hd__fa_1
XFILLER_115_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_222_clk clknet_5_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_222_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_75_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2309 t$5584 net1435 VGND VGND VPWR VPWR booth_b32_m55 sky130_fd_sc_hd__xor2_1
XFILLER_28_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1608 t$5226 net1484 VGND VGND VPWR VPWR booth_b22_m47 sky130_fd_sc_hd__xor2_1
XU$$1619 net1638 net616 net1629 net889 VGND VGND VPWR VPWR t$5232 sky130_fd_sc_hd__a22o_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_580 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_92_2 c$1828 s$1831 s$1833 VGND VGND VPWR VPWR c$2578 s$2579 sky130_fd_sc_hd__fa_1
XFILLER_170_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_85_1 c$1738 c$1740 c$1742 VGND VGND VPWR VPWR c$2520 s$2521 sky130_fd_sc_hd__fa_1
XFILLER_156_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_62_0 c$3640 c$3642 s$3645 VGND VGND VPWR VPWR c$4020 s$4021 sky130_fd_sc_hd__fa_1
Xdadda_fa_3_78_0 s$869 c$1650 c$1652 VGND VGND VPWR VPWR c$2462 s$2463 sky130_fd_sc_hd__fa_2
XU$$4433_1837 VGND VGND VPWR VPWR U$$4433_1837/HI net1837 sky130_fd_sc_hd__conb_1
XFILLER_97_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_ha_0_52_0 pp_row52_0 pp_row52_1 VGND VGND VPWR VPWR c$1 s sky130_fd_sc_hd__ha_1
XFILLER_124_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1720 net1723 VGND VGND VPWR VPWR net1720 sky130_fd_sc_hd__buf_4
Xfanout1731 net1732 VGND VGND VPWR VPWR net1731 sky130_fd_sc_hd__buf_4
Xfanout1742 net1743 VGND VGND VPWR VPWR net1742 sky130_fd_sc_hd__buf_4
XU$$4201 t$6551 net1271 VGND VGND VPWR VPWR booth_b60_m42 sky130_fd_sc_hd__xor2_1
XFILLER_77_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_213_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_213_clk
+ sky130_fd_sc_hd__clkbuf_16
XU$$4212 net1702 net435 net1692 net717 VGND VGND VPWR VPWR t$6557 sky130_fd_sc_hd__a22o_1
XFILLER_133_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1140_ clknet_leaf_15_clk booth_b8_m9 VGND VGND VPWR VPWR pp_row17_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_78_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4223 t$6562 net1270 VGND VGND VPWR VPWR booth_b60_m53 sky130_fd_sc_hd__xor2_1
XU$$4234 net1589 net435 net1580 net717 VGND VGND VPWR VPWR t$6568 sky130_fd_sc_hd__a22o_1
XU$$3500 t$6193 net1331 VGND VGND VPWR VPWR booth_b50_m34 sky130_fd_sc_hd__xor2_1
XU$$4245 t$6573 net1265 VGND VGND VPWR VPWR booth_b60_m64 sky130_fd_sc_hd__xor2_1
XU$$4256 t$6580 net1254 VGND VGND VPWR VPWR booth_b62_m1 sky130_fd_sc_hd__xor2_1
XU$$3511 net946 net489 net930 net762 VGND VGND VPWR VPWR t$6199 sky130_fd_sc_hd__a22o_1
XU$$4267 net1526 net422 net1518 net704 VGND VGND VPWR VPWR t$6586 sky130_fd_sc_hd__a22o_1
XU$$3522 t$6204 net1337 VGND VGND VPWR VPWR booth_b50_m45 sky130_fd_sc_hd__xor2_1
XFILLER_92_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_114_1 pp_row114_8 pp_row114_9 c$2738 VGND VGND VPWR VPWR c$3376 s$3377
+ sky130_fd_sc_hd__fa_1
XU$$3533 net1661 net491 net1653 net764 VGND VGND VPWR VPWR t$6210 sky130_fd_sc_hd__a22o_1
XU$$4278 t$6591 net1254 VGND VGND VPWR VPWR booth_b62_m12 sky130_fd_sc_hd__xor2_1
XFILLER_19_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1071_ clknet_leaf_52_clk booth_b8_m2 VGND VGND VPWR VPWR pp_row10_4 sky130_fd_sc_hd__dfxtp_1
XU$$4289 net1152 net420 net1142 net702 VGND VGND VPWR VPWR t$6597 sky130_fd_sc_hd__a22o_1
XU$$3544 t$6215 net1334 VGND VGND VPWR VPWR booth_b50_m56 sky130_fd_sc_hd__xor2_1
XU$$2810 net1016 net535 net999 net808 VGND VGND VPWR VPWR t$5841 sky130_fd_sc_hd__a22o_1
XU$$3555 net1549 net489 net1541 net762 VGND VGND VPWR VPWR t$6221 sky130_fd_sc_hd__a22o_1
XU$$2821 t$5846 net1378 VGND VGND VPWR VPWR booth_b40_m37 sky130_fd_sc_hd__xor2_1
XFILLER_74_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3566 notblock$6225\[2\] net48 net1332 t$6226 notblock$6225\[0\] VGND VGND VPWR
+ VPWR sel_0$6227 sky130_fd_sc_hd__a32o_4
Xdadda_fa_4_107_0 s$1971 c$2686 c$2688 VGND VGND VPWR VPWR c$3332 s$3333 sky130_fd_sc_hd__fa_1
XU$$2832 net1739 net537 net1731 net810 VGND VGND VPWR VPWR t$5852 sky130_fd_sc_hd__a22o_1
XFILLER_52_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3577 t$6233 net1325 VGND VGND VPWR VPWR booth_b52_m4 sky130_fd_sc_hd__xor2_1
XTAP_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2843 t$5857 net1380 VGND VGND VPWR VPWR booth_b40_m48 sky130_fd_sc_hd__xor2_1
XTAP_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3588 net1498 net479 net1222 net752 VGND VGND VPWR VPWR t$6239 sky130_fd_sc_hd__a22o_1
XTAP_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3599 t$6244 net1324 VGND VGND VPWR VPWR booth_b52_m15 sky130_fd_sc_hd__xor2_1
XU$$2854 net1635 net540 net1626 net813 VGND VGND VPWR VPWR t$5863 sky130_fd_sc_hd__a22o_1
XFILLER_73_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2865 t$5868 net1382 VGND VGND VPWR VPWR booth_b40_m59 sky130_fd_sc_hd__xor2_1
XU$$2876 net1383 VGND VGND VPWR VPWR notsign$5874 sky130_fd_sc_hd__inv_1
XANTENNA_170 net901 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2887 net1124 net519 net1033 net792 VGND VGND VPWR VPWR t$5881 sky130_fd_sc_hd__a22o_1
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2898 t$5886 net1367 VGND VGND VPWR VPWR booth_b42_m7 sky130_fd_sc_hd__xor2_1
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_181 net963 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_192 net1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1973_ clknet_leaf_71_clk booth_b46_m8 VGND VGND VPWR VPWR pp_row54_23 sky130_fd_sc_hd__dfxtp_1
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0924_ clknet_leaf_113_clk booth_b36_m61 VGND VGND VPWR VPWR pp_row97_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_147_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0855_ clknet_leaf_181_clk net150 VGND VGND VPWR VPWR pp_row119_6 sky130_fd_sc_hd__dfxtp_2
XFILLER_162_717 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0786_ clknet_leaf_140_clk booth_b58_m32 VGND VGND VPWR VPWR pp_row90_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_143_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_80_0 pp_row80_26 c$870 c$872 VGND VGND VPWR VPWR c$1686 s$1687 sky130_fd_sc_hd__fa_2
Xdadda_ha_1_50_8 pp_row50_24 pp_row50_25 VGND VGND VPWR VPWR c$364 s$365 sky130_fd_sc_hd__ha_2
XFILLER_143_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_783 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2456_ clknet_leaf_92_clk booth_b24_m44 VGND VGND VPWR VPWR pp_row68_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_102_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1407_ clknet_leaf_54_clk booth_b22_m11 VGND VGND VPWR VPWR pp_row33_11 sky130_fd_sc_hd__dfxtp_1
X_2387_ clknet_leaf_77_clk booth_b32_m34 VGND VGND VPWR VPWR pp_row66_16 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_204_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_204_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_84_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$805 final_adder.p_new$820 final_adder.g_new$853 final_adder.g_new$821
+ VGND VGND VPWR VPWR final_adder.g_new$933 sky130_fd_sc_hd__a21o_2
XFILLER_151_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$827 final_adder.p_new$842 final_adder.g_new$631 final_adder.g_new$843
+ VGND VGND VPWR VPWR final_adder.g_new$955 sky130_fd_sc_hd__a21o_2
X_1338_ clknet_leaf_123_clk booth_b40_m64 VGND VGND VPWR VPWR pp_row104_1 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$849 final_adder.p_new$880 final_adder.g_new$945 final_adder.g_new$881
+ VGND VGND VPWR VPWR final_adder.g_new$977 sky130_fd_sc_hd__a21o_2
XFILLER_68_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1269_ clknet_leaf_1_clk booth_b14_m12 VGND VGND VPWR VPWR pp_row26_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_25_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_95_0 s$1877 c$2590 c$2592 VGND VGND VPWR VPWR c$3260 s$3261 sky130_fd_sc_hd__fa_1
XFILLER_193_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_109_2 pp_row109_6 pp_row109_7 pp_row109_8 VGND VGND VPWR VPWR c$2714 s$2715
+ sky130_fd_sc_hd__fa_1
XFILLER_105_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput380 net380 VGND VGND VPWR VPWR o[96] sky130_fd_sc_hd__buf_2
XFILLER_10_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1005 net90 VGND VGND VPWR VPWR net1005 sky130_fd_sc_hd__buf_6
Xfanout1016 net1022 VGND VGND VPWR VPWR net1016 sky130_fd_sc_hd__buf_6
Xfanout1027 net1029 VGND VGND VPWR VPWR net1027 sky130_fd_sc_hd__buf_4
XFILLER_86_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1038 net87 VGND VGND VPWR VPWR net1038 sky130_fd_sc_hd__buf_4
XFILLER_126_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1049 net1050 VGND VGND VPWR VPWR net1049 sky130_fd_sc_hd__buf_4
XFILLER_86_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$965_1889 VGND VGND VPWR VPWR U$$965_1889/HI net1889 sky130_fd_sc_hd__conb_1
XFILLER_48_959 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_756 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2106 t$5481 net1441 VGND VGND VPWR VPWR booth_b30_m22 sky130_fd_sc_hd__xor2_1
XFILLER_142_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2117 net1058 net581 net1050 net854 VGND VGND VPWR VPWR t$5487 sky130_fd_sc_hd__a22o_1
XFILLER_15_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2128 t$5492 net1440 VGND VGND VPWR VPWR booth_b30_m33 sky130_fd_sc_hd__xor2_1
XU$$2139 net954 net583 net946 net856 VGND VGND VPWR VPWR t$5498 sky130_fd_sc_hd__a22o_1
XU$$1405 t$5123 net1488 VGND VGND VPWR VPWR booth_b20_m14 sky130_fd_sc_hd__xor2_1
XU$$1416 net1130 net627 net1114 net900 VGND VGND VPWR VPWR t$5129 sky130_fd_sc_hd__a22o_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1427 t$5134 net1486 VGND VGND VPWR VPWR booth_b20_m25 sky130_fd_sc_hd__xor2_1
XU$$1438 net1025 net630 net1017 net903 VGND VGND VPWR VPWR t$5140 sky130_fd_sc_hd__a22o_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1449 t$5145 net1489 VGND VGND VPWR VPWR booth_b20_m36 sky130_fd_sc_hd__xor2_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1099 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_2_106_0_1907 VGND VGND VPWR VPWR net1907 dadda_fa_2_106_0_1907/LO sky130_fd_sc_hd__conb_1
XFILLER_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0640_ clknet_leaf_186_clk booth_b64_m20 VGND VGND VPWR VPWR pp_row84_23 sky130_fd_sc_hd__dfxtp_1
XFILLER_171_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0571_ clknet_leaf_188_clk booth_b38_m44 VGND VGND VPWR VPWR pp_row82_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_83_1015 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2310_ clknet_leaf_84_clk booth_b24_m40 VGND VGND VPWR VPWR pp_row64_12 sky130_fd_sc_hd__dfxtp_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_934 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2241_ clknet_leaf_148_clk booth_b34_m28 VGND VGND VPWR VPWR pp_row62_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_39_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1550 net122 VGND VGND VPWR VPWR net1550 sky130_fd_sc_hd__buf_4
Xfanout1561 net1562 VGND VGND VPWR VPWR net1561 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_52_4 s$389 s$391 s$393 VGND VGND VPWR VPWR c$1358 s$1359 sky130_fd_sc_hd__fa_1
Xfanout1572 net1577 VGND VGND VPWR VPWR net1572 sky130_fd_sc_hd__buf_4
XU$$4020 t$6459 net1282 VGND VGND VPWR VPWR booth_b58_m20 sky130_fd_sc_hd__xor2_1
X_2172_ clknet_leaf_163_clk booth_b64_m60 VGND VGND VPWR VPWR pp_row124_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4031 net1077 net454 net1069 net727 VGND VGND VPWR VPWR t$6465 sky130_fd_sc_hd__a22o_1
Xfanout1583 net1584 VGND VGND VPWR VPWR net1583 sky130_fd_sc_hd__buf_4
Xfanout1594 net118 VGND VGND VPWR VPWR net1594 sky130_fd_sc_hd__buf_6
XU$$4042 t$6470 net1285 VGND VGND VPWR VPWR booth_b58_m31 sky130_fd_sc_hd__xor2_1
XU$$4053 net970 net455 net962 net728 VGND VGND VPWR VPWR t$6476 sky130_fd_sc_hd__a22o_1
X_1123_ clknet_leaf_11_clk booth_b0_m16 VGND VGND VPWR VPWR pp_row16_0 sky130_fd_sc_hd__dfxtp_1
XU$$4064 t$6481 net1289 VGND VGND VPWR VPWR booth_b58_m42 sky130_fd_sc_hd__xor2_1
XFILLER_38_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_45_3 c$268 c$270 c$272 VGND VGND VPWR VPWR c$1272 s$1273 sky130_fd_sc_hd__fa_1
XU$$3330 net1153 net497 net1145 net770 VGND VGND VPWR VPWR t$6107 sky130_fd_sc_hd__a22o_1
XFILLER_66_789 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4075 net1700 net456 net1693 net729 VGND VGND VPWR VPWR t$6487 sky130_fd_sc_hd__a22o_1
XFILLER_25_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3341 t$6112 net1339 VGND VGND VPWR VPWR booth_b48_m23 sky130_fd_sc_hd__xor2_1
XU$$4086 t$6492 net1288 VGND VGND VPWR VPWR booth_b58_m53 sky130_fd_sc_hd__xor2_1
XU$$3352 net1051 net495 net1043 net768 VGND VGND VPWR VPWR t$6118 sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_38_2 pp_row38_14 pp_row38_15 pp_row38_16 VGND VGND VPWR VPWR c$1186 s$1187
+ sky130_fd_sc_hd__fa_1
XU$$4097 net1589 net453 net1580 net726 VGND VGND VPWR VPWR t$6498 sky130_fd_sc_hd__a22o_1
XU$$3363 t$6123 net1341 VGND VGND VPWR VPWR booth_b48_m34 sky130_fd_sc_hd__xor2_1
X_1054_ clknet_leaf_56_clk booth_b4_m4 VGND VGND VPWR VPWR pp_row8_2 sky130_fd_sc_hd__dfxtp_1
XU$$3374 net943 net495 net927 net768 VGND VGND VPWR VPWR t$6129 sky130_fd_sc_hd__a22o_1
XU$$2640 t$5754 net1399 VGND VGND VPWR VPWR booth_b38_m15 sky130_fd_sc_hd__xor2_1
XU$$3385 t$6134 net1344 VGND VGND VPWR VPWR booth_b48_m45 sky130_fd_sc_hd__xor2_1
XFILLER_20_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_15_1 s$2781 s$2783 s$2785 VGND VGND VPWR VPWR c$3458 s$3459 sky130_fd_sc_hd__fa_2
XU$$3396 net1660 net498 net1652 net771 VGND VGND VPWR VPWR t$6140 sky130_fd_sc_hd__a22o_1
XFILLER_20_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2651 net1116 net544 net1107 net817 VGND VGND VPWR VPWR t$5760 sky130_fd_sc_hd__a22o_1
XU$$2662 t$5765 net1399 VGND VGND VPWR VPWR booth_b38_m26 sky130_fd_sc_hd__xor2_1
XFILLER_34_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2673 net1019 net546 net1002 net819 VGND VGND VPWR VPWR t$5771 sky130_fd_sc_hd__a22o_1
XU$$2684 t$5776 net1396 VGND VGND VPWR VPWR booth_b38_m37 sky130_fd_sc_hd__xor2_1
XU$$1950 net1201 net584 net1192 net857 VGND VGND VPWR VPWR t$5402 sky130_fd_sc_hd__a22o_1
XU$$2695 net1740 net545 net1732 net818 VGND VGND VPWR VPWR t$5782 sky130_fd_sc_hd__a22o_1
XU$$1961 t$5407 net1449 VGND VGND VPWR VPWR booth_b28_m18 sky130_fd_sc_hd__xor2_1
XU$$1972 net1091 net587 net1083 net860 VGND VGND VPWR VPWR t$5413 sky130_fd_sc_hd__a22o_1
XU$$1983 t$5418 net1451 VGND VGND VPWR VPWR booth_b28_m29 sky130_fd_sc_hd__xor2_1
XU$$1994 net983 net586 net974 net859 VGND VGND VPWR VPWR t$5424 sky130_fd_sc_hd__a22o_1
X_1956_ clknet_leaf_66_clk booth_b16_m38 VGND VGND VPWR VPWR pp_row54_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_159_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0907_ clknet_leaf_103_clk booth_b42_m54 VGND VGND VPWR VPWR pp_row96_6 sky130_fd_sc_hd__dfxtp_1
X_1887_ clknet_leaf_80_clk booth_b6_m46 VGND VGND VPWR VPWR pp_row52_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_174_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0838_ clknet_leaf_105_clk notsign$5454 VGND VGND VPWR VPWR pp_row93_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0769_ clknet_leaf_138_clk booth_b26_m64 VGND VGND VPWR VPWR pp_row90_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput108 b[49] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__buf_4
Xinput119 b[59] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__buf_2
X_2439_ clknet_leaf_75_clk booth_b56_m11 VGND VGND VPWR VPWR pp_row67_28 sky130_fd_sc_hd__dfxtp_1
XFILLER_102_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$602 final_adder.p_new$614 final_adder.p_new$606 VGND VGND VPWR VPWR
+ final_adder.p_new$730 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$613 final_adder.p_new$616 final_adder.g_new$625 final_adder.g_new$617
+ VGND VGND VPWR VPWR final_adder.g_new$741 sky130_fd_sc_hd__a21o_1
XTAP_3906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$635 final_adder.p_new$642 final_adder.g_new$659 final_adder.g_new$643
+ VGND VGND VPWR VPWR final_adder.g_new$763 sky130_fd_sc_hd__a21o_1
XTAP_3917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$646 final_adder.p_new$670 final_adder.p_new$654 VGND VGND VPWR VPWR
+ final_adder.p_new$774 sky130_fd_sc_hd__and2_1
XTAP_3928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$657 final_adder.p_new$664 final_adder.g_new$681 final_adder.g_new$665
+ VGND VGND VPWR VPWR final_adder.g_new$785 sky130_fd_sc_hd__a21o_1
XFILLER_45_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$507 net1725 net432 net1716 net714 VGND VGND VPWR VPWR t$4664 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$668 final_adder.p_new$692 final_adder.p_new$676 VGND VGND VPWR VPWR
+ final_adder.p_new$796 sky130_fd_sc_hd__and2_1
XU$$518 t$4669 net1251 VGND VGND VPWR VPWR booth_b6_m50 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$679 final_adder.p_new$686 final_adder.g_new$703 final_adder.g_new$687
+ VGND VGND VPWR VPWR final_adder.g_new$807 sky130_fd_sc_hd__a21o_1
XU$$529 net1612 net428 net1604 net710 VGND VGND VPWR VPWR t$4675 sky130_fd_sc_hd__a22o_1
Xdadda_fa_1_40_2 pp_row40_6 pp_row40_7 pp_row40_8 VGND VGND VPWR VPWR c$232 s$233
+ sky130_fd_sc_hd__fa_1
XFILLER_72_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$90 net1745 net444 net1737 net686 VGND VGND VPWR VPWR t$4452 sky130_fd_sc_hd__a22o_1
XFILLER_13_804 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_10_0 pp_row10_0 pp_row10_1 pp_row10_2 VGND VGND VPWR VPWR c$2754 s$2755
+ sky130_fd_sc_hd__fa_1
XFILLER_188_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_70 net433 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_81 net492 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_92 net530 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_114_0 net1911 pp_row114_1 pp_row114_2 VGND VGND VPWR VPWR c$2742 s$2743
+ sky130_fd_sc_hd__fa_1
XFILLER_107_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_0_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_0_0_clk sky130_fd_sc_hd__clkbuf_8
Xdadda_fa_3_62_3 s$1475 s$1477 s$1479 VGND VGND VPWR VPWR c$2340 s$2341 sky130_fd_sc_hd__fa_1
XFILLER_122_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_55_2 c$1384 s$1387 s$1389 VGND VGND VPWR VPWR c$2282 s$2283 sky130_fd_sc_hd__fa_1
XFILLER_0_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1043 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_48_1 c$1294 c$1296 c$1298 VGND VGND VPWR VPWR c$2224 s$2225 sky130_fd_sc_hd__fa_1
XFILLER_48_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_25_0 c$3492 c$3494 s$3497 VGND VGND VPWR VPWR c$3946 s$3947 sky130_fd_sc_hd__fa_1
XU$$1202 net1682 net650 net1657 net923 VGND VGND VPWR VPWR t$5019 sky130_fd_sc_hd__a22o_1
XU$$1213 t$5024 net1012 VGND VGND VPWR VPWR booth_b16_m55 sky130_fd_sc_hd__xor2_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1224 net1551 net648 net1543 net921 VGND VGND VPWR VPWR t$5030 sky130_fd_sc_hd__a22o_1
XFILLER_189_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1235 net1668 VGND VGND VPWR VPWR notblock$5035\[2\] sky130_fd_sc_hd__inv_1
XFILLER_16_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1246 t$5042 net1665 VGND VGND VPWR VPWR booth_b18_m3 sky130_fd_sc_hd__xor2_1
XFILLER_188_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1257 net1503 net635 net1494 net908 VGND VGND VPWR VPWR t$5048 sky130_fd_sc_hd__a22o_1
XFILLER_71_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1268 t$5053 net1664 VGND VGND VPWR VPWR booth_b18_m14 sky130_fd_sc_hd__xor2_1
XFILLER_189_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1279 net1131 net637 net1115 net910 VGND VGND VPWR VPWR t$5059 sky130_fd_sc_hd__a22o_1
XFILLER_188_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1810_ clknet_leaf_26_clk booth_b30_m19 VGND VGND VPWR VPWR pp_row49_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_62_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1741_ clknet_leaf_237_clk booth_b8_m39 VGND VGND VPWR VPWR pp_row47_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1040 final_adder.$signal$1169 final_adder.g_new$1050 VGND VGND VPWR
+ VPWR net361 sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$1051 final_adder.$signal$1180 final_adder.g_new$1001 VGND VGND VPWR
+ VPWR net374 sky130_fd_sc_hd__xor2_2
X_1672_ clknet_leaf_123_clk booth_b46_m60 VGND VGND VPWR VPWR pp_row106_3 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$1062 final_adder.$signal$1191 final_adder.g_new$1039 VGND VGND VPWR
+ VPWR net259 sky130_fd_sc_hd__xor2_1
XFILLER_183_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1073 final_adder.$signal$1202 final_adder.g_new$979 VGND VGND VPWR
+ VPWR net271 sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$1084 final_adder.$signal$1213 final_adder.g_new$1028 VGND VGND VPWR
+ VPWR net283 sky130_fd_sc_hd__xor2_2
X_0623_ clknet_leaf_187_clk booth_b32_m52 VGND VGND VPWR VPWR pp_row84_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_98_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_912 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0554_ clknet_leaf_189_clk booth_b58_m23 VGND VGND VPWR VPWR pp_row81_21 sky130_fd_sc_hd__dfxtp_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout809 net815 VGND VGND VPWR VPWR net809 sky130_fd_sc_hd__buf_4
XFILLER_98_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0485_ clknet_leaf_205_clk booth_b38_m41 VGND VGND VPWR VPWR pp_row79_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_61_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2224_ clknet_leaf_227_clk booth_b4_m58 VGND VGND VPWR VPWR pp_row62_2 sky130_fd_sc_hd__dfxtp_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_50_1 c$334 c$336 c$338 VGND VGND VPWR VPWR c$1328 s$1329 sky130_fd_sc_hd__fa_1
Xfanout1380 net1384 VGND VGND VPWR VPWR net1380 sky130_fd_sc_hd__buf_6
Xfanout1391 net1393 VGND VGND VPWR VPWR net1391 sky130_fd_sc_hd__buf_4
XFILLER_22_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2155_ clknet_leaf_214_clk booth_b10_m50 VGND VGND VPWR VPWR pp_row60_5 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_43_0 pp_row43_14 pp_row43_15 pp_row43_16 VGND VGND VPWR VPWR c$1242 s$1243
+ sky130_fd_sc_hd__fa_1
XU$$4485_1863 VGND VGND VPWR VPWR U$$4485_1863/HI net1863 sky130_fd_sc_hd__conb_1
XFILLER_66_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1106_ clknet_leaf_14_clk booth_b6_m8 VGND VGND VPWR VPWR pp_row14_3 sky130_fd_sc_hd__dfxtp_1
XU$$3160 t$6020 net1348 VGND VGND VPWR VPWR booth_b46_m1 sky130_fd_sc_hd__xor2_1
X_2086_ clknet_leaf_32_clk booth_b10_m48 VGND VGND VPWR VPWR pp_row58_5 sky130_fd_sc_hd__dfxtp_1
XU$$3171 net1525 net505 net1517 net778 VGND VGND VPWR VPWR t$6026 sky130_fd_sc_hd__a22o_1
XFILLER_35_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3182 t$6031 net1349 VGND VGND VPWR VPWR booth_b46_m12 sky130_fd_sc_hd__xor2_1
X_1037_ clknet_leaf_60_clk booth_b4_m1 VGND VGND VPWR VPWR pp_row5_2 sky130_fd_sc_hd__dfxtp_1
XU$$3193 net1153 net505 net1145 net778 VGND VGND VPWR VPWR t$6037 sky130_fd_sc_hd__a22o_1
XFILLER_146_1020 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2470 notblock$5665\[2\] net30 net1426 t$5666 notblock$5665\[0\] VGND VGND VPWR
+ VPWR sel_0$5667 sky130_fd_sc_hd__a32o_1
XU$$2481 t$5673 net1404 VGND VGND VPWR VPWR booth_b36_m4 sky130_fd_sc_hd__xor2_1
XU$$2492 net1497 net551 net1223 net824 VGND VGND VPWR VPWR t$5679 sky130_fd_sc_hd__a22o_1
XFILLER_167_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1780 net1474 VGND VGND VPWR VPWR notsign$5314 sky130_fd_sc_hd__inv_1
XU$$1791 net1122 net593 net1031 net866 VGND VGND VPWR VPWR t$5321 sky130_fd_sc_hd__a22o_1
XFILLER_139_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1939_ clknet_leaf_70_clk booth_b42_m11 VGND VGND VPWR VPWR pp_row53_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_135_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput90 b[32] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_72_2 s$2417 s$2419 s$2421 VGND VGND VPWR VPWR c$3126 s$3127 sky130_fd_sc_hd__fa_1
XFILLER_104_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_88_2 pp_row88_6 pp_row88_7 pp_row88_8 VGND VGND VPWR VPWR c$1004 s$1005
+ sky130_fd_sc_hd__fa_1
XFILLER_192_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_65_1 c$2354 c$2356 s$2359 VGND VGND VPWR VPWR c$3082 s$3083 sky130_fd_sc_hd__fa_1
XFILLER_115_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_42_0 s$3567 c$3978 s$3981 VGND VGND VPWR VPWR c$4236 s$4237 sky130_fd_sc_hd__fa_2
XFILLER_88_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_58_0 s$1433 c$2294 c$2296 VGND VGND VPWR VPWR c$3038 s$3039 sky130_fd_sc_hd__fa_1
XTAP_4404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$410 final_adder.p_new$416 final_adder.p_new$412 VGND VGND VPWR VPWR
+ final_adder.p_new$538 sky130_fd_sc_hd__and2_1
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$421 final_adder.p_new$422 final_adder.g_new$427 final_adder.g_new$423
+ VGND VGND VPWR VPWR final_adder.g_new$549 sky130_fd_sc_hd__a21o_1
XTAP_3703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$432 final_adder.p_new$438 final_adder.p_new$434 VGND VGND VPWR VPWR
+ final_adder.p_new$560 sky130_fd_sc_hd__and2_1
XTAP_3714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$443 final_adder.p_new$444 final_adder.g_new$449 final_adder.g_new$445
+ VGND VGND VPWR VPWR final_adder.g_new$571 sky130_fd_sc_hd__a21o_1
XTAP_3725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$454 final_adder.p_new$460 final_adder.p_new$456 VGND VGND VPWR VPWR
+ final_adder.p_new$582 sky130_fd_sc_hd__and2_1
XTAP_3736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$304 net1211 net528 net1203 net801 VGND VGND VPWR VPWR t$4561 sky130_fd_sc_hd__a22o_1
XFILLER_72_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$465 final_adder.p_new$466 final_adder.g_new$471 final_adder.g_new$467
+ VGND VGND VPWR VPWR final_adder.g_new$593 sky130_fd_sc_hd__a21o_1
XTAP_3747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$315 t$4566 net1279 VGND VGND VPWR VPWR booth_b4_m17 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$476 final_adder.p_new$482 final_adder.p_new$478 VGND VGND VPWR VPWR
+ final_adder.p_new$604 sky130_fd_sc_hd__and2_1
XTAP_3758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$326 net1097 net527 net1088 net800 VGND VGND VPWR VPWR t$4572 sky130_fd_sc_hd__a22o_1
XFILLER_17_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$487 final_adder.p_new$488 final_adder.g_new$493 final_adder.g_new$489
+ VGND VGND VPWR VPWR final_adder.g_new$615 sky130_fd_sc_hd__a21o_1
XFILLER_123_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$498 final_adder.p_new$504 final_adder.p_new$500 VGND VGND VPWR VPWR
+ final_adder.p_new$626 sky130_fd_sc_hd__and2_1
XU$$337 t$4577 net1276 VGND VGND VPWR VPWR booth_b4_m28 sky130_fd_sc_hd__xor2_1
XU$$348 net991 net528 net983 net801 VGND VGND VPWR VPWR t$4583 sky130_fd_sc_hd__a22o_1
XU$$359 t$4588 net1274 VGND VGND VPWR VPWR booth_b4_m39 sky130_fd_sc_hd__xor2_1
XFILLER_72_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_1120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1025 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1007 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_60_0 s$545 c$1434 c$1436 VGND VGND VPWR VPWR c$2318 s$2319 sky130_fd_sc_hd__fa_1
XFILLER_95_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_76_0 net1895 pp_row76_1 pp_row76_2 VGND VGND VPWR VPWR c$196 s$197 sky130_fd_sc_hd__fa_1
XFILLER_67_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0270_ clknet_leaf_217_clk booth_b46_m26 VGND VGND VPWR VPWR pp_row72_20 sky130_fd_sc_hd__dfxtp_1
XFILLER_48_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$860 net1164 net393 net1155 net659 VGND VGND VPWR VPWR t$4845 sky130_fd_sc_hd__a22o_1
XU$$1010 t$4921 net1186 VGND VGND VPWR VPWR booth_b14_m22 sky130_fd_sc_hd__xor2_1
XU$$871 t$4850 net1313 VGND VGND VPWR VPWR booth_b12_m21 sky130_fd_sc_hd__xor2_1
XU$$1021 net1055 net386 net1047 net652 VGND VGND VPWR VPWR t$4927 sky130_fd_sc_hd__a22o_1
XU$$882 net1064 net394 net1056 net660 VGND VGND VPWR VPWR t$4856 sky130_fd_sc_hd__a22o_1
XFILLER_91_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1032 t$4932 net1184 VGND VGND VPWR VPWR booth_b14_m33 sky130_fd_sc_hd__xor2_1
XFILLER_16_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$893 t$4861 net1311 VGND VGND VPWR VPWR booth_b12_m32 sky130_fd_sc_hd__xor2_1
XFILLER_189_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1043 net955 net388 net944 net654 VGND VGND VPWR VPWR t$4938 sky130_fd_sc_hd__a22o_1
XU$$1054 t$4943 net1187 VGND VGND VPWR VPWR booth_b14_m44 sky130_fd_sc_hd__xor2_1
XU$$1065 net1682 net391 net1657 net657 VGND VGND VPWR VPWR t$4949 sky130_fd_sc_hd__a22o_1
XFILLER_149_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1076 t$4954 net1191 VGND VGND VPWR VPWR booth_b14_m55 sky130_fd_sc_hd__xor2_1
XFILLER_176_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1087 net1551 net391 net1543 net657 VGND VGND VPWR VPWR t$4960 sky130_fd_sc_hd__a22o_1
XU$$1098 net1012 VGND VGND VPWR VPWR notblock$4965\[2\] sky130_fd_sc_hd__inv_1
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1724_ clknet_leaf_22_clk booth_b32_m14 VGND VGND VPWR VPWR pp_row46_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_82_1 s$3183 s$3185 s$3187 VGND VGND VPWR VPWR c$3726 s$3727 sky130_fd_sc_hd__fa_1
Xdadda_fa_2_98_1 pp_row98_3 pp_row98_4 pp_row98_5 VGND VGND VPWR VPWR c$1904 s$1905
+ sky130_fd_sc_hd__fa_1
XFILLER_172_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1655_ clknet_leaf_221_clk booth_b4_m40 VGND VGND VPWR VPWR pp_row44_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_75_0 c$3134 c$3136 c$3138 VGND VGND VPWR VPWR c$3696 s$3697 sky130_fd_sc_hd__fa_1
XFILLER_144_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0606_ clknet_leaf_173_clk booth_b52_m31 VGND VGND VPWR VPWR pp_row83_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_113_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1586_ clknet_leaf_4_clk booth_b18_m23 VGND VGND VPWR VPWR pp_row41_9 sky130_fd_sc_hd__dfxtp_1
Xfanout606 sel_0$5247 VGND VGND VPWR VPWR net606 sky130_fd_sc_hd__buf_6
Xfanout617 net618 VGND VGND VPWR VPWR net617 sky130_fd_sc_hd__clkbuf_4
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout628 net631 VGND VGND VPWR VPWR net628 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_74_8 c$184 s$187 s$189 VGND VGND VPWR VPWR c$796 s$797 sky130_fd_sc_hd__fa_2
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0537_ clknet_leaf_163_clk booth_b26_m55 VGND VGND VPWR VPWR pp_row81_5 sky130_fd_sc_hd__dfxtp_1
Xfanout639 sel_0$5037 VGND VGND VPWR VPWR net639 sky130_fd_sc_hd__buf_6
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_67_7 c$118 s$121 s$123 VGND VGND VPWR VPWR c$668 s$669 sky130_fd_sc_hd__fa_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0468_ clknet_leaf_155_clk booth_b60_m18 VGND VGND VPWR VPWR pp_row78_24 sky130_fd_sc_hd__dfxtp_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2207_ clknet_leaf_29_clk booth_b36_m25 VGND VGND VPWR VPWR pp_row61_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_85_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_1041 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0399_ clknet_leaf_191_clk booth_b46_m30 VGND VGND VPWR VPWR pp_row76_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_67_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2138_ clknet_leaf_143_clk booth_b56_m53 VGND VGND VPWR VPWR pp_row109_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_148_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2069_ clknet_leaf_35_clk booth_b40_m17 VGND VGND VPWR VPWR pp_row57_20 sky130_fd_sc_hd__dfxtp_1
XFILLER_23_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_93_0 pp_row93_0 pp_row93_1 pp_row93_2 VGND VGND VPWR VPWR c$1038 s$1039
+ sky130_fd_sc_hd__fa_1
XFILLER_150_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_5_13__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_5_13__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_2_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3907 t$6401 net1292 VGND VGND VPWR VPWR booth_b56_m32 sky130_fd_sc_hd__xor2_1
XTAP_4256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$240 final_adder.$signal$1104 final_adder.$signal$1105 VGND VGND VPWR
+ VPWR final_adder.p_new$368 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$251 final_adder.$signal$1095 final_adder.$signal$10 final_adder.$signal$12
+ VGND VGND VPWR VPWR final_adder.g_new$379 sky130_fd_sc_hd__a21o_1
XTAP_3522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3918 net962 net464 net954 net737 VGND VGND VPWR VPWR t$6407 sky130_fd_sc_hd__a22o_1
XTAP_4267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3929 t$6412 net1298 VGND VGND VPWR VPWR booth_b56_m43 sky130_fd_sc_hd__xor2_1
XU$$101 t$4457 net1570 VGND VGND VPWR VPWR booth_b0_m47 sky130_fd_sc_hd__xor2_1
XTAP_4278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_105_0 c$3812 c$3814 s$3817 VGND VGND VPWR VPWR c$4106 s$4107 sky130_fd_sc_hd__fa_1
XTAP_3533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$262 final_adder.p_new$264 final_adder.p_new$262 VGND VGND VPWR VPWR
+ final_adder.p_new$390 sky130_fd_sc_hd__and2_1
XTAP_4289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$112 net1642 net449 net1633 net691 VGND VGND VPWR VPWR t$4463 sky130_fd_sc_hd__a22o_1
XTAP_3544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$273 final_adder.p_new$272 final_adder.g_new$275 final_adder.g_new$273
+ VGND VGND VPWR VPWR final_adder.g_new$401 sky130_fd_sc_hd__a21o_1
XTAP_3555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$284 final_adder.p_new$286 final_adder.p_new$284 VGND VGND VPWR VPWR
+ final_adder.p_new$412 sky130_fd_sc_hd__and2_1
XU$$123 t$4468 net1576 VGND VGND VPWR VPWR booth_b0_m58 sky130_fd_sc_hd__xor2_1
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$134 net1527 net444 net1758 net686 VGND VGND VPWR VPWR t$4474 sky130_fd_sc_hd__a22o_1
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$295 final_adder.p_new$294 final_adder.g_new$297 final_adder.g_new$295
+ VGND VGND VPWR VPWR final_adder.g_new$423 sky130_fd_sc_hd__a21o_1
XU$$145 net1231 net624 net1127 net897 VGND VGND VPWR VPWR t$4480 sky130_fd_sc_hd__a22o_1
XTAP_3577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_25_3 c$1054 c$1056 s$1059 VGND VGND VPWR VPWR c$2044 s$2045 sky130_fd_sc_hd__fa_1
XU$$156 t$4485 net1390 VGND VGND VPWR VPWR booth_b2_m6 sky130_fd_sc_hd__xor2_1
XTAP_3599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$167 net1211 net623 net1203 net896 VGND VGND VPWR VPWR t$4491 sky130_fd_sc_hd__a22o_1
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$178 t$4496 net1389 VGND VGND VPWR VPWR booth_b2_m17 sky130_fd_sc_hd__xor2_1
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$189 net1097 net620 net1088 net893 VGND VGND VPWR VPWR t$4502 sky130_fd_sc_hd__a22o_1
XFILLER_60_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_92_0 c$3760 c$3762 s$3765 VGND VGND VPWR VPWR c$4080 s$4081 sky130_fd_sc_hd__fa_1
XFILLER_127_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1440_ clknet_leaf_54_clk booth_b6_m29 VGND VGND VPWR VPWR pp_row35_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_141_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1371_ clknet_leaf_110_clk booth_b46_m58 VGND VGND VPWR VPWR pp_row104_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_110_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0322_ clknet_leaf_182_clk net144 VGND VGND VPWR VPWR pp_row113_9 sky130_fd_sc_hd__dfxtp_2
XFILLER_96_957 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0253_ clknet_leaf_210_clk booth_b16_m56 VGND VGND VPWR VPWR pp_row72_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0184_ clknet_leaf_147_clk booth_b12_m58 VGND VGND VPWR VPWR pp_row70_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_91_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$690 net2 net1238 VGND VGND VPWR VPWR sel_1$4758 sky130_fd_sc_hd__xor2_1
XFILLER_63_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_1_80_8 pp_row80_24 pp_row80_25 VGND VGND VPWR VPWR c$904 s$905 sky130_fd_sc_hd__ha_1
XFILLER_129_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1707_ clknet_leaf_236_clk booth_b0_m46 VGND VGND VPWR VPWR pp_row46_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_144_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1638_ clknet_leaf_240_clk booth_b20_m23 VGND VGND VPWR VPWR pp_row43_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout403 net408 VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__clkbuf_8
Xfanout414 net415 VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__clkbuf_4
X_1569_ clknet_leaf_20_clk booth_b34_m6 VGND VGND VPWR VPWR pp_row40_17 sky130_fd_sc_hd__dfxtp_1
Xfanout425 sel_0$6577 VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_72_5 pp_row72_26 pp_row72_27 pp_row72_28 VGND VGND VPWR VPWR c$754 s$755
+ sky130_fd_sc_hd__fa_1
Xfanout436 net437 VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__buf_4
XFILLER_58_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout447 net449 VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__buf_2
Xfanout458 net459 VGND VGND VPWR VPWR net458 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_65_4 pp_row65_30 pp_row65_31 pp_row65_32 VGND VGND VPWR VPWR c$626 s$627
+ sky130_fd_sc_hd__fa_1
Xfanout469 net471 VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__buf_4
XFILLER_101_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_58_3 pp_row58_20 pp_row58_21 pp_row58_22 VGND VGND VPWR VPWR c$498 s$499
+ sky130_fd_sc_hd__fa_1
Xdadda_fa_4_35_2 s$2121 s$2123 s$2125 VGND VGND VPWR VPWR c$2904 s$2905 sky130_fd_sc_hd__fa_1
XFILLER_73_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_28_1 c$2058 c$2060 s$2063 VGND VGND VPWR VPWR c$2860 s$2861 sky130_fd_sc_hd__fa_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_846 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_892 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4405 t$6656 net1823 VGND VGND VPWR VPWR booth_b64_m7 sky130_fd_sc_hd__xor2_1
XFILLER_77_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4416 net1209 sel_0$6647 net1197 net695 VGND VGND VPWR VPWR t$6662 sky130_fd_sc_hd__a22o_1
Xfanout970 net972 VGND VGND VPWR VPWR net970 sky130_fd_sc_hd__buf_6
XTAP_4020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout981 net93 VGND VGND VPWR VPWR net981 sky130_fd_sc_hd__buf_8
XFILLER_65_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_0_60_3 pp_row60_9 pp_row60_10 pp_row60_11 VGND VGND VPWR VPWR c$46 s$47
+ sky130_fd_sc_hd__fa_1
XTAP_4031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4427 t$6667 net1834 VGND VGND VPWR VPWR booth_b64_m18 sky130_fd_sc_hd__xor2_1
XFILLER_37_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout992 net993 VGND VGND VPWR VPWR net992 sky130_fd_sc_hd__buf_4
XU$$4438 net1095 sel_0$6647 net1086 net695 VGND VGND VPWR VPWR t$6673 sky130_fd_sc_hd__a22o_1
XTAP_4042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_ha_3_17_1 pp_row17_3 pp_row17_4 VGND VGND VPWR VPWR c$1984 s$1985 sky130_fd_sc_hd__ha_1
XU$$3704 net50 net1321 VGND VGND VPWR VPWR sel_1$6298 sky130_fd_sc_hd__xor2_4
XFILLER_92_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4449 t$6678 net1845 VGND VGND VPWR VPWR booth_b64_m29 sky130_fd_sc_hd__xor2_1
XTAP_4053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3715 net1674 net468 net1563 net741 VGND VGND VPWR VPWR t$6304 sky130_fd_sc_hd__a22o_1
XTAP_4064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3726 t$6309 net1304 VGND VGND VPWR VPWR booth_b54_m10 sky130_fd_sc_hd__xor2_1
XFILLER_58_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3737 net1169 net468 net1160 net741 VGND VGND VPWR VPWR t$6315 sky130_fd_sc_hd__a22o_1
XTAP_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_30_1 pp_row30_17 c$1082 c$1084 VGND VGND VPWR VPWR c$2080 s$2081 sky130_fd_sc_hd__fa_1
XU$$3748 t$6320 net1300 VGND VGND VPWR VPWR booth_b54_m21 sky130_fd_sc_hd__xor2_1
XTAP_4097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3759 net1069 net469 net1061 net742 VGND VGND VPWR VPWR t$6326 sky130_fd_sc_hd__a22o_1
XTAP_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_330 net687 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdadda_fa_3_23_0 pp_row23_2 pp_row23_3 pp_row23_4 VGND VGND VPWR VPWR c$2022 s$2023
+ sky130_fd_sc_hd__fa_1
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_341 net782 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_352 net915 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_363 net1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_374 net1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_385 net1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_396 net1552 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0940_ clknet_leaf_184_clk net253 VGND VGND VPWR VPWR pp_row97_17 sky130_fd_sc_hd__dfxtp_4
XFILLER_186_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0871_ clknet_leaf_141_clk booth_b50_m44 VGND VGND VPWR VPWR pp_row94_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_173_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_848 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2472_ clknet_leaf_98_clk booth_b52_m16 VGND VGND VPWR VPWR pp_row68_25 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_82_4 s$925 s$927 s$929 VGND VGND VPWR VPWR c$1718 s$1719 sky130_fd_sc_hd__fa_1
XFILLER_5_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1423_ clknet_leaf_56_clk booth_b16_m18 VGND VGND VPWR VPWR pp_row34_8 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_75_3 c$796 s$799 s$801 VGND VGND VPWR VPWR c$1632 s$1633 sky130_fd_sc_hd__fa_1
XFILLER_130_829 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1354_ clknet_leaf_4_clk booth_b2_m29 VGND VGND VPWR VPWR pp_row31_1 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_68_2 c$664 c$666 c$668 VGND VGND VPWR VPWR c$1546 s$1547 sky130_fd_sc_hd__fa_1
XFILLER_96_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_45_1 s$2961 s$2963 s$2965 VGND VGND VPWR VPWR c$3578 s$3579 sky130_fd_sc_hd__fa_1
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0305_ clknet_leaf_225_clk booth_b48_m25 VGND VGND VPWR VPWR pp_row73_20 sky130_fd_sc_hd__dfxtp_1
X_1285_ clknet_leaf_1_clk booth_b8_m19 VGND VGND VPWR VPWR pp_row27_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_37_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_38_0 c$2912 c$2914 c$2916 VGND VGND VPWR VPWR c$3548 s$3549 sky130_fd_sc_hd__fa_1
XFILLER_23_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0236_ clknet_leaf_151_clk booth_b44_m27 VGND VGND VPWR VPWR pp_row71_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_92_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_112_0 c$3356 c$3358 c$3360 VGND VGND VPWR VPWR c$3844 s$3845 sky130_fd_sc_hd__fa_1
XFILLER_166_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4419_1830 VGND VGND VPWR VPWR U$$4419_1830/HI net1830 sky130_fd_sc_hd__conb_1
XFILLER_30_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1209 net68 VGND VGND VPWR VPWR net1209 sky130_fd_sc_hd__buf_6
XFILLER_132_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_70_2 pp_row70_20 pp_row70_21 pp_row70_22 VGND VGND VPWR VPWR c$712 s$713
+ sky130_fd_sc_hd__fa_1
XFILLER_8_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_63_1 pp_row63_20 pp_row63_21 pp_row63_22 VGND VGND VPWR VPWR c$584 s$585
+ sky130_fd_sc_hd__fa_1
XFILLER_75_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_40_0 s$1217 c$2150 c$2152 VGND VGND VPWR VPWR c$2930 s$2931 sky130_fd_sc_hd__fa_1
XFILLER_75_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_56_0 pp_row56_8 pp_row56_9 pp_row56_10 VGND VGND VPWR VPWR c$456 s$457
+ sky130_fd_sc_hd__fa_2
XFILLER_189_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1609 net1698 net618 net1690 net891 VGND VGND VPWR VPWR t$5227 sky130_fd_sc_hd__a22o_1
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_92_3 s$1835 s$1837 s$1839 VGND VGND VPWR VPWR c$2580 s$2581 sky130_fd_sc_hd__fa_1
XFILLER_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_85_2 c$1744 s$1747 s$1749 VGND VGND VPWR VPWR c$2522 s$2523 sky130_fd_sc_hd__fa_1
XFILLER_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_78_1 c$1654 c$1656 c$1658 VGND VGND VPWR VPWR c$2464 s$2465 sky130_fd_sc_hd__fa_1
Xdadda_fa_6_55_0 c$3612 c$3614 s$3617 VGND VGND VPWR VPWR c$4006 s$4007 sky130_fd_sc_hd__fa_1
Xfanout1710 net105 VGND VGND VPWR VPWR net1710 sky130_fd_sc_hd__buf_6
XFILLER_2_496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1721 net1723 VGND VGND VPWR VPWR net1721 sky130_fd_sc_hd__clkbuf_4
Xfanout1732 net102 VGND VGND VPWR VPWR net1732 sky130_fd_sc_hd__buf_4
XFILLER_104_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1743 net1744 VGND VGND VPWR VPWR net1743 sky130_fd_sc_hd__buf_4
XU$$4202 net1743 net440 net1735 net722 VGND VGND VPWR VPWR t$6552 sky130_fd_sc_hd__a22o_1
XU$$4213 t$6557 net1267 VGND VGND VPWR VPWR booth_b60_m48 sky130_fd_sc_hd__xor2_1
XFILLER_172_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4224 net1636 net439 net1625 net721 VGND VGND VPWR VPWR t$6563 sky130_fd_sc_hd__a22o_1
XFILLER_66_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4235 t$6568 net1265 VGND VGND VPWR VPWR booth_b60_m59 sky130_fd_sc_hd__xor2_1
XFILLER_133_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3501 net984 net485 net975 net758 VGND VGND VPWR VPWR t$6194 sky130_fd_sc_hd__a22o_1
XFILLER_19_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4246 net1268 VGND VGND VPWR VPWR notsign$6574 sky130_fd_sc_hd__inv_1
XU$$4257 net1129 net422 net1037 net704 VGND VGND VPWR VPWR t$6581 sky130_fd_sc_hd__a22o_1
XFILLER_37_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3512 t$6199 net1334 VGND VGND VPWR VPWR booth_b50_m40 sky130_fd_sc_hd__xor2_1
XU$$4268 t$6586 net1259 VGND VGND VPWR VPWR booth_b62_m7 sky130_fd_sc_hd__xor2_1
XU$$3523 net1717 net490 net1708 net763 VGND VGND VPWR VPWR t$6205 sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_114_2 c$2740 s$2743 s$2745 VGND VGND VPWR VPWR c$3378 s$3379 sky130_fd_sc_hd__fa_1
X_1070_ clknet_leaf_52_clk booth_b6_m4 VGND VGND VPWR VPWR pp_row10_3 sky130_fd_sc_hd__dfxtp_1
XU$$3534 t$6210 net1335 VGND VGND VPWR VPWR booth_b50_m51 sky130_fd_sc_hd__xor2_1
XU$$4279 net1205 net418 net1196 net700 VGND VGND VPWR VPWR t$6592 sky130_fd_sc_hd__a22o_1
XFILLER_92_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2800 net1070 net539 net1062 net812 VGND VGND VPWR VPWR t$5836 sky130_fd_sc_hd__a22o_1
XU$$3545 net1608 net486 net1600 net759 VGND VGND VPWR VPWR t$6216 sky130_fd_sc_hd__a22o_1
XU$$2811 t$5841 net1376 VGND VGND VPWR VPWR booth_b40_m32 sky130_fd_sc_hd__xor2_1
XFILLER_80_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3556 t$6221 net1334 VGND VGND VPWR VPWR booth_b50_m62 sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_107_1 c$2690 c$2692 s$2695 VGND VGND VPWR VPWR c$3334 s$3335 sky130_fd_sc_hd__fa_1
XTAP_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2822 net958 net537 net951 net810 VGND VGND VPWR VPWR t$5847 sky130_fd_sc_hd__a22o_1
XFILLER_65_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3567 net48 net1332 VGND VGND VPWR VPWR sel_1$6228 sky130_fd_sc_hd__xor2_4
XTAP_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2833 t$5852 net1378 VGND VGND VPWR VPWR booth_b40_m43 sky130_fd_sc_hd__xor2_1
XU$$3578 net1677 net481 net1566 net754 VGND VGND VPWR VPWR t$6234 sky130_fd_sc_hd__a22o_1
XU$$2844 net1689 net538 net1681 net811 VGND VGND VPWR VPWR t$5858 sky130_fd_sc_hd__a22o_1
XU$$3589 t$6239 net1320 VGND VGND VPWR VPWR booth_b52_m10 sky130_fd_sc_hd__xor2_1
XTAP_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2855 t$5863 net1382 VGND VGND VPWR VPWR booth_b40_m54 sky130_fd_sc_hd__xor2_1
XTAP_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2866 net1584 net541 net1558 net814 VGND VGND VPWR VPWR t$5869 sky130_fd_sc_hd__a22o_1
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_160 net849 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2877 net1379 VGND VGND VPWR VPWR notblock$5875\[0\] sky130_fd_sc_hd__inv_1
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2888 t$5881 net1367 VGND VGND VPWR VPWR booth_b42_m2 sky130_fd_sc_hd__xor2_1
XANTENNA_171 net909 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2899 net1516 net523 net1509 net796 VGND VGND VPWR VPWR t$5887 sky130_fd_sc_hd__a22o_1
XANTENNA_182 net963 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_193 net1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1972_ clknet_leaf_138_clk booth_b50_m58 VGND VGND VPWR VPWR pp_row108_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0923_ clknet_leaf_112_clk booth_b34_m63 VGND VGND VPWR VPWR pp_row97_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_187_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0854_ clknet_leaf_142_clk booth_b58_m35 VGND VGND VPWR VPWR pp_row93_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_174_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0785_ clknet_leaf_138_clk booth_b56_m34 VGND VGND VPWR VPWR pp_row90_16 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_80_1 c$874 c$876 c$878 VGND VGND VPWR VPWR c$1688 s$1689 sky130_fd_sc_hd__fa_1
XFILLER_103_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2455_ clknet_leaf_92_clk booth_b22_m46 VGND VGND VPWR VPWR pp_row68_10 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_73_0 s$185 c$744 c$746 VGND VGND VPWR VPWR c$1602 s$1603 sky130_fd_sc_hd__fa_1
XFILLER_170_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1406_ clknet_leaf_109_clk booth_b52_m52 VGND VGND VPWR VPWR pp_row104_7 sky130_fd_sc_hd__dfxtp_1
X_2386_ clknet_leaf_77_clk booth_b30_m36 VGND VGND VPWR VPWR pp_row66_15 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$817 final_adder.p_new$832 final_adder.g_new$865 final_adder.g_new$833
+ VGND VGND VPWR VPWR final_adder.g_new$945 sky130_fd_sc_hd__a21o_2
XFILLER_68_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1337_ clknet_leaf_0_clk booth_b8_m22 VGND VGND VPWR VPWR pp_row30_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_60_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$839 final_adder.p_new$870 final_adder.g_new$935 final_adder.g_new$871
+ VGND VGND VPWR VPWR final_adder.g_new$967 sky130_fd_sc_hd__a21o_2
XFILLER_56_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4449_1845 VGND VGND VPWR VPWR U$$4449_1845/HI net1845 sky130_fd_sc_hd__conb_1
X_1268_ clknet_leaf_1_clk booth_b12_m14 VGND VGND VPWR VPWR pp_row26_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_43_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0219_ clknet_leaf_200_clk booth_b14_m57 VGND VGND VPWR VPWR pp_row71_4 sky130_fd_sc_hd__dfxtp_1
X_1199_ clknet_leaf_245_clk net170 VGND VGND VPWR VPWR pp_row21_11 sky130_fd_sc_hd__dfxtp_2
XFILLER_51_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_140_clk clknet_5_25__leaf_clk VGND VGND VPWR VPWR clknet_leaf_140_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_165_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_95_1 c$2594 c$2596 s$2599 VGND VGND VPWR VPWR c$3262 s$3263 sky130_fd_sc_hd__fa_1
XFILLER_137_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1030 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_72_0 s$3687 c$4038 s$4041 VGND VGND VPWR VPWR c$4296 s$4297 sky130_fd_sc_hd__fa_1
Xdadda_fa_4_88_0 s$1793 c$2534 c$2536 VGND VGND VPWR VPWR c$3218 s$3219 sky130_fd_sc_hd__fa_1
XFILLER_193_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_109_3 pp_row109_9 pp_row109_10 pp_row109_11 VGND VGND VPWR VPWR c$2716
+ s$2717 sky130_fd_sc_hd__fa_1
Xoutput370 net370 VGND VGND VPWR VPWR o[87] sky130_fd_sc_hd__buf_2
Xoutput381 net381 VGND VGND VPWR VPWR o[97] sky130_fd_sc_hd__buf_2
Xfanout1006 net1008 VGND VGND VPWR VPWR net1006 sky130_fd_sc_hd__buf_6
XFILLER_0_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1017 net1018 VGND VGND VPWR VPWR net1017 sky130_fd_sc_hd__buf_4
XFILLER_0_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1028 net1029 VGND VGND VPWR VPWR net1028 sky130_fd_sc_hd__buf_4
Xfanout1039 net1040 VGND VGND VPWR VPWR net1039 sky130_fd_sc_hd__clkbuf_8
XFILLER_120_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2107 net1100 net580 net1091 net853 VGND VGND VPWR VPWR t$5482 sky130_fd_sc_hd__a22o_1
XU$$2118 t$5487 net1442 VGND VGND VPWR VPWR booth_b30_m28 sky130_fd_sc_hd__xor2_1
XU$$2129 net991 net581 net983 net854 VGND VGND VPWR VPWR t$5493 sky130_fd_sc_hd__a22o_1
XU$$1406 net1179 net629 net1170 net902 VGND VGND VPWR VPWR t$5124 sky130_fd_sc_hd__a22o_1
XFILLER_28_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1417 t$5129 net1486 VGND VGND VPWR VPWR booth_b20_m20 sky130_fd_sc_hd__xor2_1
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1428 net1072 net628 net1064 net901 VGND VGND VPWR VPWR t$5135 sky130_fd_sc_hd__a22o_1
XFILLER_128_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1439 t$5140 net1489 VGND VGND VPWR VPWR booth_b20_m31 sky130_fd_sc_hd__xor2_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_131_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_131_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_156_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_90_0 s$1025 c$1794 c$1796 VGND VGND VPWR VPWR c$2558 s$2559 sky130_fd_sc_hd__fa_2
XFILLER_125_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0570_ clknet_leaf_188_clk booth_b36_m46 VGND VGND VPWR VPWR pp_row82_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2240_ clknet_leaf_227_clk booth_b32_m30 VGND VGND VPWR VPWR pp_row62_16 sky130_fd_sc_hd__dfxtp_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1540 net1542 VGND VGND VPWR VPWR net1540 sky130_fd_sc_hd__buf_4
Xfanout1551 net1552 VGND VGND VPWR VPWR net1551 sky130_fd_sc_hd__buf_4
XFILLER_111_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_198_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_198_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2171_ clknet_leaf_136_clk booth_b62_m47 VGND VGND VPWR VPWR pp_row109_9 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_52_5 s$395 s$397 s$399 VGND VGND VPWR VPWR c$1360 s$1361 sky130_fd_sc_hd__fa_2
XU$$4010 t$6454 net1282 VGND VGND VPWR VPWR booth_b58_m15 sky130_fd_sc_hd__xor2_1
Xfanout1562 net1563 VGND VGND VPWR VPWR net1562 sky130_fd_sc_hd__buf_4
XU$$4021 net1119 net454 net1112 net727 VGND VGND VPWR VPWR t$6460 sky130_fd_sc_hd__a22o_1
XFILLER_93_521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1573 net1574 VGND VGND VPWR VPWR net1573 sky130_fd_sc_hd__buf_4
Xfanout1584 net1585 VGND VGND VPWR VPWR net1584 sky130_fd_sc_hd__buf_4
XU$$4032 t$6465 net1286 VGND VGND VPWR VPWR booth_b58_m26 sky130_fd_sc_hd__xor2_1
Xfanout1595 net1598 VGND VGND VPWR VPWR net1595 sky130_fd_sc_hd__buf_4
X_1122_ clknet_leaf_248_clk net163 VGND VGND VPWR VPWR pp_row15_8 sky130_fd_sc_hd__dfxtp_2
XFILLER_76_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4043 net1021 net456 net1004 net729 VGND VGND VPWR VPWR t$6471 sky130_fd_sc_hd__a22o_1
XU$$4054 t$6476 net1290 VGND VGND VPWR VPWR booth_b58_m37 sky130_fd_sc_hd__xor2_1
XU$$3320 net1205 net493 net1196 net766 VGND VGND VPWR VPWR t$6102 sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_45_4 c$274 s$277 s$279 VGND VGND VPWR VPWR c$1274 s$1275 sky130_fd_sc_hd__fa_1
XU$$4065 net1742 net457 net1734 net730 VGND VGND VPWR VPWR t$6482 sky130_fd_sc_hd__a22o_1
XU$$3331 t$6107 net1343 VGND VGND VPWR VPWR booth_b48_m18 sky130_fd_sc_hd__xor2_1
XU$$4076 t$6487 net1288 VGND VGND VPWR VPWR booth_b58_m48 sky130_fd_sc_hd__xor2_1
XU$$3342 net1090 net493 net1082 net766 VGND VGND VPWR VPWR t$6113 sky130_fd_sc_hd__a22o_1
XU$$4087 net1634 net456 net1624 net729 VGND VGND VPWR VPWR t$6493 sky130_fd_sc_hd__a22o_1
XFILLER_19_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3353 t$6118 net1340 VGND VGND VPWR VPWR booth_b48_m29 sky130_fd_sc_hd__xor2_1
XU$$4098 t$6498 net1284 VGND VGND VPWR VPWR booth_b58_m59 sky130_fd_sc_hd__xor2_1
X_1053_ clknet_leaf_53_clk booth_b2_m6 VGND VGND VPWR VPWR pp_row8_1 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_38_3 pp_row38_17 pp_row38_18 pp_row38_19 VGND VGND VPWR VPWR c$1188 s$1189
+ sky130_fd_sc_hd__fa_1
XU$$3364 net984 net494 net975 net767 VGND VGND VPWR VPWR t$6124 sky130_fd_sc_hd__a22o_1
XFILLER_20_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2630 t$5749 net1394 VGND VGND VPWR VPWR booth_b38_m10 sky130_fd_sc_hd__xor2_1
XU$$3375 t$6129 net1342 VGND VGND VPWR VPWR booth_b48_m40 sky130_fd_sc_hd__xor2_1
XU$$3386 net1717 net498 net1708 net771 VGND VGND VPWR VPWR t$6135 sky130_fd_sc_hd__a22o_1
XU$$2641 net1171 net549 net1162 net822 VGND VGND VPWR VPWR t$5755 sky130_fd_sc_hd__a22o_1
XU$$3397 t$6140 net1344 VGND VGND VPWR VPWR booth_b48_m51 sky130_fd_sc_hd__xor2_1
XFILLER_179_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2652 t$5760 net1395 VGND VGND VPWR VPWR booth_b38_m21 sky130_fd_sc_hd__xor2_1
XU$$2663 net1067 net549 net1058 net822 VGND VGND VPWR VPWR t$5766 sky130_fd_sc_hd__a22o_1
XU$$2674 t$5771 net1397 VGND VGND VPWR VPWR booth_b38_m32 sky130_fd_sc_hd__xor2_1
XFILLER_34_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2685 net959 net545 net950 net818 VGND VGND VPWR VPWR t$5777 sky130_fd_sc_hd__a22o_1
XU$$1940 net1516 net588 net1508 net861 VGND VGND VPWR VPWR t$5397 sky130_fd_sc_hd__a22o_1
XU$$1951 t$5402 net1448 VGND VGND VPWR VPWR booth_b28_m13 sky130_fd_sc_hd__xor2_1
XU$$2696 t$5782 net1396 VGND VGND VPWR VPWR booth_b38_m43 sky130_fd_sc_hd__xor2_1
XU$$1962 net1140 net586 net1132 net859 VGND VGND VPWR VPWR t$5408 sky130_fd_sc_hd__a22o_1
XU$$1973 t$5413 net1451 VGND VGND VPWR VPWR booth_b28_m24 sky130_fd_sc_hd__xor2_1
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1984 net1042 net588 net1026 net861 VGND VGND VPWR VPWR t$5419 sky130_fd_sc_hd__a22o_1
XU$$1995 t$5424 net1450 VGND VGND VPWR VPWR booth_b28_m35 sky130_fd_sc_hd__xor2_1
X_1955_ clknet_leaf_66_clk booth_b14_m40 VGND VGND VPWR VPWR pp_row54_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_174_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0906_ clknet_leaf_103_clk booth_b40_m56 VGND VGND VPWR VPWR pp_row96_5 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_122_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_122_clk
+ sky130_fd_sc_hd__clkbuf_16
X_1886_ clknet_leaf_80_clk booth_b4_m48 VGND VGND VPWR VPWR pp_row52_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0837_ clknet_leaf_194_clk net248 VGND VGND VPWR VPWR pp_row92_20 sky130_fd_sc_hd__dfxtp_2
XFILLER_134_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0768_ clknet_leaf_194_clk net244 VGND VGND VPWR VPWR pp_row89_21 sky130_fd_sc_hd__dfxtp_2
XFILLER_143_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0699_ clknet_leaf_181_clk net148 VGND VGND VPWR VPWR pp_row117_7 sky130_fd_sc_hd__dfxtp_2
XFILLER_102_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput109 b[4] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_4
X_2438_ clknet_leaf_75_clk booth_b54_m13 VGND VGND VPWR VPWR pp_row67_27 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$603 final_adder.p_new$606 final_adder.g_new$615 final_adder.g_new$607
+ VGND VGND VPWR VPWR final_adder.g_new$731 sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_189_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_189_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_111_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_1072 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$614 final_adder.p_new$626 final_adder.p_new$618 VGND VGND VPWR VPWR
+ final_adder.p_new$742 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$625 final_adder.p_new$628 final_adder.g_new$383 final_adder.g_new$629
+ VGND VGND VPWR VPWR final_adder.g_new$753 sky130_fd_sc_hd__a21o_4
XFILLER_29_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2369_ clknet_leaf_198_clk net218 VGND VGND VPWR VPWR pp_row65_33 sky130_fd_sc_hd__dfxtp_1
XTAP_3907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$636 final_adder.p_new$660 final_adder.p_new$644 VGND VGND VPWR VPWR
+ final_adder.p_new$764 sky130_fd_sc_hd__and2_1
XFILLER_56_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$647 final_adder.p_new$654 final_adder.g_new$671 final_adder.g_new$655
+ VGND VGND VPWR VPWR final_adder.g_new$775 sky130_fd_sc_hd__a21o_1
XTAP_3929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$658 final_adder.p_new$682 final_adder.p_new$666 VGND VGND VPWR VPWR
+ final_adder.p_new$786 sky130_fd_sc_hd__and2_1
XU$$508 t$4664 net1251 VGND VGND VPWR VPWR booth_b6_m45 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$669 final_adder.p_new$676 final_adder.g_new$693 final_adder.g_new$677
+ VGND VGND VPWR VPWR final_adder.g_new$797 sky130_fd_sc_hd__a21o_1
XU$$519 net1657 net433 net1649 net715 VGND VGND VPWR VPWR t$4670 sky130_fd_sc_hd__a22o_1
XFILLER_186_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$80 net964 net442 net956 net684 VGND VGND VPWR VPWR t$4447 sky130_fd_sc_hd__a22o_1
XU$$91 t$4452 net1570 VGND VGND VPWR VPWR booth_b0_m42 sky130_fd_sc_hd__xor2_1
XFILLER_13_816 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4503_1872 VGND VGND VPWR VPWR U$$4503_1872/HI net1872 sky130_fd_sc_hd__conb_1
XFILLER_184_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_113_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_113_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_60 net400 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_71 net441 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_82 net509 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_93 net530 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_107_0 pp_row107_3 pp_row107_4 pp_row107_5 VGND VGND VPWR VPWR c$2694 s$2695
+ sky130_fd_sc_hd__fa_1
XFILLER_107_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_55_3 s$1391 s$1393 s$1395 VGND VGND VPWR VPWR c$2284 s$2285 sky130_fd_sc_hd__fa_1
XFILLER_82_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_48_2 c$1300 s$1303 s$1305 VGND VGND VPWR VPWR c$2226 s$2227 sky130_fd_sc_hd__fa_1
XFILLER_75_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_18_0 c$3464 c$3466 s$3469 VGND VGND VPWR VPWR c$3932 s$3933 sky130_fd_sc_hd__fa_2
XFILLER_62_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1203 t$5019 net1011 VGND VGND VPWR VPWR booth_b16_m50 sky130_fd_sc_hd__xor2_1
XFILLER_15_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1214 net1614 net649 net1606 net922 VGND VGND VPWR VPWR t$5025 sky130_fd_sc_hd__a22o_1
XFILLER_188_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1225 t$5030 net1012 VGND VGND VPWR VPWR booth_b16_m61 sky130_fd_sc_hd__xor2_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1236 net1668 notblock$5035\[1\] VGND VGND VPWR VPWR t$5036 sky130_fd_sc_hd__and2_1
XU$$1247 net936 net637 net1676 net910 VGND VGND VPWR VPWR t$5043 sky130_fd_sc_hd__a22o_1
XFILLER_188_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1258 t$5048 net1662 VGND VGND VPWR VPWR booth_b18_m9 sky130_fd_sc_hd__xor2_1
XU$$1269 net1179 net638 net1170 net911 VGND VGND VPWR VPWR t$5054 sky130_fd_sc_hd__a22o_1
XFILLER_148_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_104_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_104_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_15_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1740_ clknet_leaf_236_clk booth_b6_m41 VGND VGND VPWR VPWR pp_row47_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_12_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1030 final_adder.$signal$1159 final_adder.g_new$1055 VGND VGND VPWR
+ VPWR net350 sky130_fd_sc_hd__xor2_2
XFILLER_183_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1041 final_adder.$signal$1170 final_adder.g_new$1011 VGND VGND VPWR
+ VPWR net363 sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$1052 final_adder.$signal$1181 final_adder.g_new$1044 VGND VGND VPWR
+ VPWR net375 sky130_fd_sc_hd__xor2_2
X_1671_ clknet_leaf_241_clk booth_b34_m10 VGND VGND VPWR VPWR pp_row44_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_116_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1063 final_adder.$signal$1192 final_adder.g_new$989 VGND VGND VPWR
+ VPWR net260 sky130_fd_sc_hd__xor2_1
XFILLER_172_846 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1074 final_adder.$signal$1203 final_adder.g_new$1033 VGND VGND VPWR
+ VPWR net272 sky130_fd_sc_hd__xor2_2
X_0622_ clknet_leaf_164_clk notsign$6294 VGND VGND VPWR VPWR pp_row117_0 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$1085 final_adder.$signal$1214 final_adder.g_new$967 VGND VGND VPWR
+ VPWR net284 sky130_fd_sc_hd__xor2_2
XFILLER_98_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0553_ clknet_leaf_171_clk booth_b56_m25 VGND VGND VPWR VPWR pp_row81_20 sky130_fd_sc_hd__dfxtp_1
XFILLER_113_924 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0484_ clknet_leaf_156_clk booth_b36_m43 VGND VGND VPWR VPWR pp_row79_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_98_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2223_ clknet_leaf_227_clk booth_b2_m60 VGND VGND VPWR VPWR pp_row62_1 sky130_fd_sc_hd__dfxtp_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1370 net1371 VGND VGND VPWR VPWR net1370 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_50_2 c$340 c$342 c$344 VGND VGND VPWR VPWR c$1330 s$1331 sky130_fd_sc_hd__fa_1
XFILLER_22_1128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1381 net1384 VGND VGND VPWR VPWR net1381 sky130_fd_sc_hd__buf_6
X_2154_ clknet_leaf_214_clk booth_b8_m52 VGND VGND VPWR VPWR pp_row60_4 sky130_fd_sc_hd__dfxtp_1
Xfanout1392 net1393 VGND VGND VPWR VPWR net1392 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_43_1 pp_row43_17 pp_row43_18 pp_row43_19 VGND VGND VPWR VPWR c$1244 s$1245
+ sky130_fd_sc_hd__fa_1
XFILLER_66_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1105_ clknet_leaf_121_clk booth_b56_m46 VGND VGND VPWR VPWR pp_row102_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_66_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_20_0 c$2804 c$2806 c$2808 VGND VGND VPWR VPWR c$3476 s$3477 sky130_fd_sc_hd__fa_1
X_2085_ clknet_leaf_32_clk booth_b8_m50 VGND VGND VPWR VPWR pp_row58_4 sky130_fd_sc_hd__dfxtp_1
XU$$3150 net1360 VGND VGND VPWR VPWR notsign$6014 sky130_fd_sc_hd__inv_1
Xdadda_fa_2_36_0 pp_row36_5 pp_row36_6 pp_row36_7 VGND VGND VPWR VPWR c$1158 s$1159
+ sky130_fd_sc_hd__fa_1
XFILLER_4_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3161 net1125 net501 net1034 net774 VGND VGND VPWR VPWR t$6021 sky130_fd_sc_hd__a22o_1
XU$$3172 t$6026 net1353 VGND VGND VPWR VPWR booth_b46_m7 sky130_fd_sc_hd__xor2_1
X_1036_ clknet_leaf_61_clk booth_b2_m3 VGND VGND VPWR VPWR pp_row5_1 sky130_fd_sc_hd__dfxtp_1
XU$$3183 net1202 net501 net1193 net774 VGND VGND VPWR VPWR t$6032 sky130_fd_sc_hd__a22o_1
XU$$3194 t$6037 net1353 VGND VGND VPWR VPWR booth_b46_m18 sky130_fd_sc_hd__xor2_1
XU$$2460 t$5661 net1428 VGND VGND VPWR VPWR booth_b34_m62 sky130_fd_sc_hd__xor2_1
XFILLER_35_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2471 net30 net1427 VGND VGND VPWR VPWR sel_1$5668 sky130_fd_sc_hd__xor2_1
XU$$2482 net1671 net551 net1560 net824 VGND VGND VPWR VPWR t$5674 sky130_fd_sc_hd__a22o_1
XU$$2493 t$5679 net1403 VGND VGND VPWR VPWR booth_b36_m10 sky130_fd_sc_hd__xor2_1
XU$$1770 net1579 net608 net1553 net881 VGND VGND VPWR VPWR t$5309 sky130_fd_sc_hd__a22o_1
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1781 net1471 VGND VGND VPWR VPWR notblock$5315\[0\] sky130_fd_sc_hd__inv_1
XU$$1792 t$5321 net1457 VGND VGND VPWR VPWR booth_b26_m2 sky130_fd_sc_hd__xor2_1
XFILLER_50_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1938_ clknet_leaf_136_clk booth_b44_m64 VGND VGND VPWR VPWR pp_row108_1 sky130_fd_sc_hd__dfxtp_1
X_1869_ clknet_leaf_66_clk booth_b28_m23 VGND VGND VPWR VPWR pp_row51_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput80 b[23] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__buf_4
XFILLER_174_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput91 b[33] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__buf_6
XFILLER_66_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_88_3 pp_row88_9 pp_row88_10 pp_row88_11 VGND VGND VPWR VPWR c$1006 s$1007
+ sky130_fd_sc_hd__fa_1
XFILLER_131_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_65_2 s$2361 s$2363 s$2365 VGND VGND VPWR VPWR c$3084 s$3085 sky130_fd_sc_hd__fa_1
XFILLER_192_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_58_1 c$2298 c$2300 s$2303 VGND VGND VPWR VPWR c$3040 s$3041 sky130_fd_sc_hd__fa_1
XTAP_4405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$400 final_adder.p_new$406 final_adder.p_new$402 VGND VGND VPWR VPWR
+ final_adder.p_new$528 sky130_fd_sc_hd__and2_1
Xdadda_fa_7_35_0 s$3539 c$3964 s$3967 VGND VGND VPWR VPWR c$4222 s$4223 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$411 final_adder.p_new$412 final_adder.g_new$417 final_adder.g_new$413
+ VGND VGND VPWR VPWR final_adder.g_new$539 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$422 final_adder.p_new$428 final_adder.p_new$424 VGND VGND VPWR VPWR
+ final_adder.p_new$550 sky130_fd_sc_hd__and2_1
XTAP_3704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$433 final_adder.p_new$434 final_adder.g_new$439 final_adder.g_new$435
+ VGND VGND VPWR VPWR final_adder.g_new$561 sky130_fd_sc_hd__a21o_1
XTAP_3715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$444 final_adder.p_new$450 final_adder.p_new$446 VGND VGND VPWR VPWR
+ final_adder.p_new$572 sky130_fd_sc_hd__and2_1
XFILLER_57_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$455 final_adder.p_new$456 final_adder.g_new$461 final_adder.g_new$457
+ VGND VGND VPWR VPWR final_adder.g_new$583 sky130_fd_sc_hd__a21o_1
XTAP_3737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$305 t$4561 net1274 VGND VGND VPWR VPWR booth_b4_m12 sky130_fd_sc_hd__xor2_1
XFILLER_83_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$466 final_adder.p_new$472 final_adder.p_new$468 VGND VGND VPWR VPWR
+ final_adder.p_new$594 sky130_fd_sc_hd__and2_1
XTAP_3748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$316 net1149 net532 net1143 net805 VGND VGND VPWR VPWR t$4567 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$477 final_adder.p_new$478 final_adder.g_new$483 final_adder.g_new$479
+ VGND VGND VPWR VPWR final_adder.g_new$605 sky130_fd_sc_hd__a21o_1
XTAP_3759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$327 t$4572 net1273 VGND VGND VPWR VPWR booth_b4_m23 sky130_fd_sc_hd__xor2_1
XFILLER_72_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$488 final_adder.p_new$494 final_adder.p_new$490 VGND VGND VPWR VPWR
+ final_adder.p_new$616 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$499 final_adder.p_new$500 final_adder.g_new$505 final_adder.g_new$501
+ VGND VGND VPWR VPWR final_adder.g_new$627 sky130_fd_sc_hd__a21o_1
XU$$338 net1050 net531 net1042 net804 VGND VGND VPWR VPWR t$4578 sky130_fd_sc_hd__a22o_1
XU$$349 t$4583 net1276 VGND VGND VPWR VPWR booth_b4_m34 sky130_fd_sc_hd__xor2_1
XFILLER_26_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_60_1 c$1438 c$1440 c$1442 VGND VGND VPWR VPWR c$2320 s$2321 sky130_fd_sc_hd__fa_1
XFILLER_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_53_0 s$419 c$1350 c$1352 VGND VGND VPWR VPWR c$2262 s$2263 sky130_fd_sc_hd__fa_1
XFILLER_121_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_0_69_0 pp_row69_0 pp_row69_1 pp_row69_2 VGND VGND VPWR VPWR c$144 s$145
+ sky130_fd_sc_hd__fa_1
XFILLER_35_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$850 net1221 net396 net1212 net662 VGND VGND VPWR VPWR t$4840 sky130_fd_sc_hd__a22o_1
XU$$861 t$4845 net1310 VGND VGND VPWR VPWR booth_b12_m16 sky130_fd_sc_hd__xor2_1
XU$$1000 t$4916 net1183 VGND VGND VPWR VPWR booth_b14_m17 sky130_fd_sc_hd__xor2_1
XFILLER_90_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1011 net1100 net388 net1091 net654 VGND VGND VPWR VPWR t$4922 sky130_fd_sc_hd__a22o_1
XU$$872 net1108 net397 net1100 net663 VGND VGND VPWR VPWR t$4851 sky130_fd_sc_hd__a22o_1
XU$$1022 t$4927 net1184 VGND VGND VPWR VPWR booth_b14_m28 sky130_fd_sc_hd__xor2_1
XU$$883 t$4856 net1311 VGND VGND VPWR VPWR booth_b12_m27 sky130_fd_sc_hd__xor2_1
XU$$1033 net990 net386 net982 net652 VGND VGND VPWR VPWR t$4933 sky130_fd_sc_hd__a22o_1
XFILLER_44_782 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$894 net999 net396 net991 net662 VGND VGND VPWR VPWR t$4862 sky130_fd_sc_hd__a22o_1
XU$$1044 t$4938 net1186 VGND VGND VPWR VPWR booth_b14_m39 sky130_fd_sc_hd__xor2_1
XFILLER_189_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1055 net1720 net390 net1711 net656 VGND VGND VPWR VPWR t$4944 sky130_fd_sc_hd__a22o_1
XFILLER_188_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1066 t$4949 net1191 VGND VGND VPWR VPWR booth_b14_m50 sky130_fd_sc_hd__xor2_1
XFILLER_189_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1077 net1615 net392 net1607 net658 VGND VGND VPWR VPWR t$4955 sky130_fd_sc_hd__a22o_1
XU$$1088 t$4960 net1188 VGND VGND VPWR VPWR booth_b14_m61 sky130_fd_sc_hd__xor2_1
XFILLER_32_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1099 net1012 notblock$4965\[1\] VGND VGND VPWR VPWR t$4966 sky130_fd_sc_hd__and2_1
XFILLER_31_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_110_0 s$3839 c$4114 s$4117 VGND VGND VPWR VPWR c$4372 s$4373 sky130_fd_sc_hd__fa_1
XFILLER_78_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1723_ clknet_leaf_21_clk booth_b30_m16 VGND VGND VPWR VPWR pp_row46_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_172_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_98_2 pp_row98_6 pp_row98_7 pp_row98_8 VGND VGND VPWR VPWR c$1906 s$1907
+ sky130_fd_sc_hd__fa_1
XFILLER_7_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1654_ clknet_leaf_221_clk booth_b2_m42 VGND VGND VPWR VPWR pp_row44_1 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_75_1 s$3141 s$3143 s$3145 VGND VGND VPWR VPWR c$3698 s$3699 sky130_fd_sc_hd__fa_2
XFILLER_137_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0605_ clknet_leaf_188_clk booth_b50_m33 VGND VGND VPWR VPWR pp_row83_16 sky130_fd_sc_hd__dfxtp_1
X_1585_ clknet_leaf_243_clk booth_b16_m25 VGND VGND VPWR VPWR pp_row41_8 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_68_0 c$3092 c$3094 c$3096 VGND VGND VPWR VPWR c$3668 s$3669 sky130_fd_sc_hd__fa_1
Xfanout607 net609 VGND VGND VPWR VPWR net607 sky130_fd_sc_hd__buf_6
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout618 sel_0$5177 VGND VGND VPWR VPWR net618 sky130_fd_sc_hd__buf_6
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0536_ clknet_leaf_163_clk booth_b24_m57 VGND VGND VPWR VPWR pp_row81_4 sky130_fd_sc_hd__dfxtp_1
Xfanout629 net630 VGND VGND VPWR VPWR net629 sky130_fd_sc_hd__clkbuf_8
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0467_ clknet_leaf_155_clk booth_b58_m20 VGND VGND VPWR VPWR pp_row78_23 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_67_8 s$125 s$127 s$129 VGND VGND VPWR VPWR c$670 s$671 sky130_fd_sc_hd__fa_2
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2206_ clknet_leaf_29_clk booth_b34_m27 VGND VGND VPWR VPWR pp_row61_17 sky130_fd_sc_hd__dfxtp_1
X_0398_ clknet_leaf_190_clk booth_b44_m32 VGND VGND VPWR VPWR pp_row76_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2137_ clknet_leaf_26_clk booth_b40_m19 VGND VGND VPWR VPWR pp_row59_20 sky130_fd_sc_hd__dfxtp_1
XFILLER_96_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2068_ clknet_leaf_43_clk booth_b38_m19 VGND VGND VPWR VPWR pp_row57_19 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_6_7_0 c$3420 c$3422 s$3425 VGND VGND VPWR VPWR c$3910 s$3911 sky130_fd_sc_hd__fa_1
X_1019_ clknet_leaf_249_clk net129 VGND VGND VPWR VPWR pp_row0_2 sky130_fd_sc_hd__dfxtp_2
XFILLER_22_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2290 net1713 net574 net1704 net847 VGND VGND VPWR VPWR t$5575 sky130_fd_sc_hd__a22o_1
XFILLER_139_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_1057 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_93_1 pp_row93_3 pp_row93_4 pp_row93_5 VGND VGND VPWR VPWR c$1040 s$1041
+ sky130_fd_sc_hd__fa_1
XFILLER_162_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_70_0 s$1577 c$2390 c$2392 VGND VGND VPWR VPWR c$3110 s$3111 sky130_fd_sc_hd__fa_1
XFILLER_162_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_86_0 net1899 pp_row86_1 pp_row86_2 VGND VGND VPWR VPWR c$978 s$979 sky130_fd_sc_hd__fa_1
XFILLER_131_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4388_1813 VGND VGND VPWR VPWR U$$4388_1813/HI net1813 sky130_fd_sc_hd__conb_1
Xdadda_ha_2_106_1 pp_row106_3 pp_row106_4 VGND VGND VPWR VPWR c$1968 s$1969 sky130_fd_sc_hd__ha_1
XTAP_4224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3908 net1003 net462 net995 net735 VGND VGND VPWR VPWR t$6402 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$230 final_adder.$signal$1114 final_adder.$signal$1115 VGND VGND VPWR
+ VPWR final_adder.p_new$358 sky130_fd_sc_hd__and2_1
XTAP_4257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3919 t$6407 net1296 VGND VGND VPWR VPWR booth_b56_m38 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$241 final_adder.$signal$1105 final_adder.$signal$30 final_adder.$signal$32
+ VGND VGND VPWR VPWR final_adder.g_new$369 sky130_fd_sc_hd__a21o_1
XTAP_4268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$252 final_adder.$signal$1092 final_adder.$signal$1093 VGND VGND VPWR
+ VPWR final_adder.p_new$380 sky130_fd_sc_hd__and2_1
XTAP_3523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$102 net1695 net444 net1687 net686 VGND VGND VPWR VPWR t$4458 sky130_fd_sc_hd__a22o_1
XFILLER_73_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$263 final_adder.p_new$262 final_adder.g_new$265 final_adder.g_new$263
+ VGND VGND VPWR VPWR final_adder.g_new$391 sky130_fd_sc_hd__a21o_1
XU$$113 t$4463 net1576 VGND VGND VPWR VPWR booth_b0_m53 sky130_fd_sc_hd__xor2_1
XTAP_3545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$274 final_adder.p_new$276 final_adder.p_new$274 VGND VGND VPWR VPWR
+ final_adder.p_new$402 sky130_fd_sc_hd__and2_1
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$285 final_adder.p_new$284 final_adder.g_new$287 final_adder.g_new$285
+ VGND VGND VPWR VPWR final_adder.g_new$413 sky130_fd_sc_hd__a21o_1
XFILLER_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$124 net1586 net445 net1578 net687 VGND VGND VPWR VPWR t$4469 sky130_fd_sc_hd__a22o_1
XTAP_3567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$135 t$4474 net1571 VGND VGND VPWR VPWR booth_b0_m64 sky130_fd_sc_hd__xor2_1
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$296 final_adder.p_new$298 final_adder.p_new$296 VGND VGND VPWR VPWR
+ final_adder.p_new$424 sky130_fd_sc_hd__and2_1
XU$$146 t$4480 net1390 VGND VGND VPWR VPWR booth_b2_m1 sky130_fd_sc_hd__xor2_1
XTAP_3578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$157 net1523 net624 net1515 net897 VGND VGND VPWR VPWR t$4486 sky130_fd_sc_hd__a22o_1
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$168 t$4491 net1389 VGND VGND VPWR VPWR booth_b2_m12 sky130_fd_sc_hd__xor2_1
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$179 net1149 net623 net1143 net896 VGND VGND VPWR VPWR t$4497 sky130_fd_sc_hd__a22o_1
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_85_0 c$3732 c$3734 s$3737 VGND VGND VPWR VPWR c$4066 s$4067 sky130_fd_sc_hd__fa_1
XFILLER_126_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1370_ clknet_leaf_244_clk net181 VGND VGND VPWR VPWR pp_row31_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_96_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0321_ clknet_leaf_200_clk booth_b20_m54 VGND VGND VPWR VPWR pp_row74_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_96_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0252_ clknet_leaf_209_clk booth_b14_m58 VGND VGND VPWR VPWR pp_row72_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_64_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0183_ clknet_leaf_147_clk booth_b10_m60 VGND VGND VPWR VPWR pp_row70_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_24_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_888 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$680 net1535 net411 net1527 net677 VGND VGND VPWR VPWR t$4752 sky130_fd_sc_hd__a22o_1
XU$$691 net1885 net404 net1231 net670 VGND VGND VPWR VPWR t$4759 sky130_fd_sc_hd__a22o_1
XFILLER_189_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1239_1757 VGND VGND VPWR VPWR U$$1239_1757/HI net1757 sky130_fd_sc_hd__conb_1
X_1706_ clknet_leaf_236_clk net196 VGND VGND VPWR VPWR pp_row45_23 sky130_fd_sc_hd__dfxtp_1
X_1637_ clknet_leaf_240_clk booth_b18_m25 VGND VGND VPWR VPWR pp_row43_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_160_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_903 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout404 net407 VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__buf_4
XFILLER_98_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1568_ clknet_leaf_7_clk booth_b32_m8 VGND VGND VPWR VPWR pp_row40_16 sky130_fd_sc_hd__dfxtp_1
Xfanout415 net417 VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__buf_4
Xfanout426 net427 VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_72_6 pp_row72_29 pp_row72_30 c$164 VGND VGND VPWR VPWR c$756 s$757 sky130_fd_sc_hd__fa_1
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout437 net441 VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__buf_4
XFILLER_58_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout448 net449 VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__buf_4
X_0519_ clknet_leaf_166_clk booth_b46_m34 VGND VGND VPWR VPWR pp_row80_16 sky130_fd_sc_hd__dfxtp_1
Xfanout459 sel_0$6437 VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__clkbuf_4
XFILLER_58_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_65_5 pp_row65_33 c$84 c$86 VGND VGND VPWR VPWR c$628 s$629 sky130_fd_sc_hd__fa_2
XFILLER_101_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1499_ clknet_leaf_41_clk booth_b34_m3 VGND VGND VPWR VPWR pp_row37_17 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_58_4 pp_row58_23 pp_row58_24 pp_row58_25 VGND VGND VPWR VPWR c$500 s$501
+ sky130_fd_sc_hd__fa_1
XFILLER_67_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_93_clk clknet_5_25__leaf_clk VGND VGND VPWR VPWR clknet_leaf_93_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_27_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_28_2 s$2065 s$2067 s$2069 VGND VGND VPWR VPWR c$2862 s$2863 sky130_fd_sc_hd__fa_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4406 net1518 sel_0$6647 net1507 net694 VGND VGND VPWR VPWR t$6657 sky130_fd_sc_hd__a22o_1
Xfanout960 net95 VGND VGND VPWR VPWR net960 sky130_fd_sc_hd__buf_4
Xfanout971 net972 VGND VGND VPWR VPWR net971 sky130_fd_sc_hd__buf_2
XTAP_4010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4417 t$6662 net1829 VGND VGND VPWR VPWR booth_b64_m13 sky130_fd_sc_hd__xor2_1
XTAP_4021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout982 net983 VGND VGND VPWR VPWR net982 sky130_fd_sc_hd__buf_4
XU$$4428 net1141 sel_0$6647 net1135 net694 VGND VGND VPWR VPWR t$6668 sky130_fd_sc_hd__a22o_1
XTAP_4032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout993 net91 VGND VGND VPWR VPWR net993 sky130_fd_sc_hd__clkbuf_4
XTAP_4043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4439 t$6673 net1840 VGND VGND VPWR VPWR booth_b64_m24 sky130_fd_sc_hd__xor2_1
XTAP_4054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3705 net1797 net472 net1233 net745 VGND VGND VPWR VPWR t$6299 sky130_fd_sc_hd__a22o_1
XFILLER_86_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3716 t$6304 net1300 VGND VGND VPWR VPWR booth_b54_m5 sky130_fd_sc_hd__xor2_1
XTAP_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3727 net1226 net475 net1217 net748 VGND VGND VPWR VPWR t$6310 sky130_fd_sc_hd__a22o_1
XTAP_4076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3738 t$6315 net1309 VGND VGND VPWR VPWR booth_b54_m16 sky130_fd_sc_hd__xor2_1
XTAP_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3749 net1111 net468 net1102 net741 VGND VGND VPWR VPWR t$6321 sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_84_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_84_clk sky130_fd_sc_hd__clkbuf_16
XTAP_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_30_2 c$1086 c$1088 s$1091 VGND VGND VPWR VPWR c$2082 s$2083 sky130_fd_sc_hd__fa_1
XFILLER_18_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_320 net601 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_331 net707 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1778_1766 VGND VGND VPWR VPWR U$$1778_1766/HI net1766 sky130_fd_sc_hd__conb_1
XANTENNA_342 net839 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdadda_fa_3_23_1 pp_row23_5 pp_row23_6 pp_row23_7 VGND VGND VPWR VPWR c$2024 s$2025
+ sky130_fd_sc_hd__fa_1
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_353 net931 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_364 net1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_16_0 pp_row16_0 pp_row16_1 pp_row16_2 VGND VGND VPWR VPWR c$1978 s$1979
+ sky130_fd_sc_hd__fa_1
XFILLER_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_375 net1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_386 net1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_397 net1559 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0870_ clknet_leaf_104_clk booth_b48_m46 VGND VGND VPWR VPWR pp_row94_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_186_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1060 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2471_ clknet_leaf_98_clk booth_b50_m18 VGND VGND VPWR VPWR pp_row68_24 sky130_fd_sc_hd__dfxtp_1
XFILLER_5_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_82_5 s$931 s$933 s$935 VGND VGND VPWR VPWR c$1720 s$1721 sky130_fd_sc_hd__fa_1
XFILLER_141_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1422_ clknet_leaf_55_clk booth_b14_m20 VGND VGND VPWR VPWR pp_row34_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_142_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2737_1781 VGND VGND VPWR VPWR U$$2737_1781/HI net1781 sky130_fd_sc_hd__conb_1
Xdadda_fa_2_75_4 s$803 s$805 s$807 VGND VGND VPWR VPWR c$1634 s$1635 sky130_fd_sc_hd__fa_1
X_1353_ clknet_leaf_4_clk booth_b0_m31 VGND VGND VPWR VPWR pp_row31_0 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_68_3 c$670 s$673 s$675 VGND VGND VPWR VPWR c$1548 s$1549 sky130_fd_sc_hd__fa_1
XFILLER_96_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0304_ clknet_leaf_225_clk booth_b46_m27 VGND VGND VPWR VPWR pp_row73_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1284_ clknet_leaf_1_clk booth_b6_m21 VGND VGND VPWR VPWR pp_row27_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_110_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_38_1 s$2919 s$2921 s$2923 VGND VGND VPWR VPWR c$3550 s$3551 sky130_fd_sc_hd__fa_1
XFILLER_55_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0235_ clknet_leaf_151_clk booth_b42_m29 VGND VGND VPWR VPWR pp_row71_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_83_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_75_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_75_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_36_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_587 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_112_1 s$3363 s$3365 s$3367 VGND VGND VPWR VPWR c$3846 s$3847 sky130_fd_sc_hd__fa_1
XFILLER_192_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0999_ clknet_leaf_164_clk booth_b58_m64 VGND VGND VPWR VPWR pp_row122_1 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_105_0 c$3314 c$3316 c$3318 VGND VGND VPWR VPWR c$3816 s$3817 sky130_fd_sc_hd__fa_1
XFILLER_30_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_70_3 pp_row70_23 pp_row70_24 pp_row70_25 VGND VGND VPWR VPWR c$714 s$715
+ sky130_fd_sc_hd__fa_1
XFILLER_59_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_63_2 pp_row63_23 pp_row63_24 pp_row63_25 VGND VGND VPWR VPWR c$586 s$587
+ sky130_fd_sc_hd__fa_1
XFILLER_86_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_40_1 c$2154 c$2156 s$2159 VGND VGND VPWR VPWR c$2932 s$2933 sky130_fd_sc_hd__fa_1
Xdadda_fa_1_56_1 pp_row56_11 pp_row56_12 pp_row56_13 VGND VGND VPWR VPWR c$458 s$459
+ sky130_fd_sc_hd__fa_2
XFILLER_189_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_33_0 s$1133 c$2094 c$2096 VGND VGND VPWR VPWR c$2888 s$2889 sky130_fd_sc_hd__fa_1
Xclkbuf_leaf_66_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_66_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_28_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_49_0 pp_row49_0 pp_row49_1 pp_row49_2 VGND VGND VPWR VPWR c$332 s$333
+ sky130_fd_sc_hd__fa_2
XFILLER_28_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_85_3 s$1751 s$1753 s$1755 VGND VGND VPWR VPWR c$2524 s$2525 sky130_fd_sc_hd__fa_1
XFILLER_163_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_78_2 c$1660 s$1663 s$1665 VGND VGND VPWR VPWR c$2466 s$2467 sky130_fd_sc_hd__fa_1
XFILLER_111_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1700 net1702 VGND VGND VPWR VPWR net1700 sky130_fd_sc_hd__buf_4
XFILLER_85_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1711 net1714 VGND VGND VPWR VPWR net1711 sky130_fd_sc_hd__buf_4
Xfanout1722 net1723 VGND VGND VPWR VPWR net1722 sky130_fd_sc_hd__buf_4
XFILLER_104_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1733 net1736 VGND VGND VPWR VPWR net1733 sky130_fd_sc_hd__buf_6
XFILLER_78_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1744 net101 VGND VGND VPWR VPWR net1744 sky130_fd_sc_hd__buf_4
XFILLER_27_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_48_0 c$3584 c$3586 s$3589 VGND VGND VPWR VPWR c$3992 s$3993 sky130_fd_sc_hd__fa_1
XU$$4203 t$6552 net1271 VGND VGND VPWR VPWR booth_b60_m43 sky130_fd_sc_hd__xor2_1
XFILLER_78_777 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4214 net1692 net435 net1685 net717 VGND VGND VPWR VPWR t$6558 sky130_fd_sc_hd__a22o_1
XFILLER_65_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4225 t$6563 net1270 VGND VGND VPWR VPWR booth_b60_m54 sky130_fd_sc_hd__xor2_1
Xfanout790 net791 VGND VGND VPWR VPWR net790 sky130_fd_sc_hd__clkbuf_8
XU$$4236 net1580 net436 net1554 net718 VGND VGND VPWR VPWR t$6569 sky130_fd_sc_hd__a22o_1
XU$$3502 t$6194 net1331 VGND VGND VPWR VPWR booth_b50_m35 sky130_fd_sc_hd__xor2_1
XFILLER_59_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4247 net1265 VGND VGND VPWR VPWR notblock$6575\[0\] sky130_fd_sc_hd__inv_1
XFILLER_133_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4258 t$6581 net1259 VGND VGND VPWR VPWR booth_b62_m2 sky130_fd_sc_hd__xor2_1
XU$$3513 net929 net490 net1750 net763 VGND VGND VPWR VPWR t$6200 sky130_fd_sc_hd__a22o_1
XFILLER_1_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3524 t$6205 net1335 VGND VGND VPWR VPWR booth_b50_m46 sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_57_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_57_clk sky130_fd_sc_hd__clkbuf_16
XU$$4269 net1518 net421 net1507 net703 VGND VGND VPWR VPWR t$6587 sky130_fd_sc_hd__a22o_1
XU$$3535 net1653 net491 net1645 net764 VGND VGND VPWR VPWR t$6211 sky130_fd_sc_hd__a22o_1
XU$$2801 t$5836 net1384 VGND VGND VPWR VPWR booth_b40_m27 sky130_fd_sc_hd__xor2_1
XU$$3546 t$6216 net1330 VGND VGND VPWR VPWR booth_b50_m57 sky130_fd_sc_hd__xor2_1
XU$$2812 net1005 net536 net991 net809 VGND VGND VPWR VPWR t$5842 sky130_fd_sc_hd__a22o_1
XU$$3557 net1541 net489 net1533 net762 VGND VGND VPWR VPWR t$6222 sky130_fd_sc_hd__a22o_1
XTAP_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2823 t$5847 net1378 VGND VGND VPWR VPWR booth_b40_m38 sky130_fd_sc_hd__xor2_1
XU$$3568 net1795 net479 net1233 net752 VGND VGND VPWR VPWR t$6229 sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_107_2 s$2697 s$2699 s$2701 VGND VGND VPWR VPWR c$3336 s$3337 sky130_fd_sc_hd__fa_1
XTAP_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2834 net1731 net537 net1722 net810 VGND VGND VPWR VPWR t$5853 sky130_fd_sc_hd__a22o_1
XFILLER_46_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3579 t$6234 net1325 VGND VGND VPWR VPWR booth_b52_m5 sky130_fd_sc_hd__xor2_1
XTAP_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2845 t$5858 net1380 VGND VGND VPWR VPWR booth_b40_m49 sky130_fd_sc_hd__xor2_1
XU$$2856 net1627 net540 net1619 net813 VGND VGND VPWR VPWR t$5864 sky130_fd_sc_hd__a22o_1
XTAP_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2867 t$5869 net1382 VGND VGND VPWR VPWR booth_b40_m60 sky130_fd_sc_hd__xor2_1
XANTENNA_150 net794 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2878 net37 VGND VGND VPWR VPWR notblock$5875\[1\] sky130_fd_sc_hd__inv_1
XFILLER_60_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_161 net861 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2889 net1033 net520 net934 net793 VGND VGND VPWR VPWR t$5882 sky130_fd_sc_hd__a22o_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_172 net909 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_183 net968 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_194 net1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1971_ clknet_leaf_72_clk booth_b44_m10 VGND VGND VPWR VPWR pp_row54_22 sky130_fd_sc_hd__dfxtp_1
XFILLER_61_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0922_ clknet_leaf_112_clk notsign$5594 VGND VGND VPWR VPWR pp_row97_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0853_ clknet_leaf_144_clk booth_b56_m37 VGND VGND VPWR VPWR pp_row93_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_128_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0784_ clknet_leaf_138_clk booth_b54_m36 VGND VGND VPWR VPWR pp_row90_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_127_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_80_2 c$880 c$882 c$884 VGND VGND VPWR VPWR c$1690 s$1691 sky130_fd_sc_hd__fa_1
XFILLER_115_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2454_ clknet_leaf_141_clk booth_b20_m48 VGND VGND VPWR VPWR pp_row68_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_142_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_73_1 c$748 c$750 c$752 VGND VGND VPWR VPWR c$1604 s$1605 sky130_fd_sc_hd__fa_1
XFILLER_64_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1405_ clknet_leaf_51_clk booth_b20_m13 VGND VGND VPWR VPWR pp_row33_10 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_50_0 c$2984 c$2986 c$2988 VGND VGND VPWR VPWR c$3596 s$3597 sky130_fd_sc_hd__fa_1
X_2385_ clknet_leaf_83_clk booth_b28_m38 VGND VGND VPWR VPWR pp_row66_14 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_66_0 s$119 c$618 c$620 VGND VGND VPWR VPWR c$1518 s$1519 sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$807 final_adder.p_new$822 final_adder.g_new$855 final_adder.g_new$823
+ VGND VGND VPWR VPWR final_adder.g_new$935 sky130_fd_sc_hd__a21o_1
X_1336_ clknet_leaf_247_clk booth_b6_m24 VGND VGND VPWR VPWR pp_row30_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_68_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$829 final_adder.p_new$844 final_adder.g_new$633 final_adder.g_new$845
+ VGND VGND VPWR VPWR final_adder.g_new$957 sky130_fd_sc_hd__a21o_2
XFILLER_112_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput1 a[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_4
X_1267_ clknet_leaf_2_clk booth_b10_m16 VGND VGND VPWR VPWR pp_row26_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_84_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_48_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_48_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_65_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0218_ clknet_leaf_199_clk booth_b12_m59 VGND VGND VPWR VPWR pp_row71_3 sky130_fd_sc_hd__dfxtp_1
X_1198_ clknet_leaf_51_clk booth_b20_m1 VGND VGND VPWR VPWR pp_row21_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_101_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_95_2 s$2601 s$2603 s$2605 VGND VGND VPWR VPWR c$3264 s$3265 sky130_fd_sc_hd__fa_1
XFILLER_192_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1042 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_88_1 c$2538 c$2540 s$2543 VGND VGND VPWR VPWR c$3220 s$3221 sky130_fd_sc_hd__fa_1
XFILLER_145_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_65_0 s$3659 c$4024 s$4027 VGND VGND VPWR VPWR c$4282 s$4283 sky130_fd_sc_hd__fa_1
XFILLER_117_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput360 net360 VGND VGND VPWR VPWR o[78] sky130_fd_sc_hd__buf_2
XFILLER_161_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput371 net371 VGND VGND VPWR VPWR o[88] sky130_fd_sc_hd__buf_2
Xoutput382 net382 VGND VGND VPWR VPWR o[98] sky130_fd_sc_hd__buf_2
Xfanout1007 net1008 VGND VGND VPWR VPWR net1007 sky130_fd_sc_hd__buf_6
Xfanout1018 net1022 VGND VGND VPWR VPWR net1018 sky130_fd_sc_hd__buf_6
Xfanout1029 net1030 VGND VGND VPWR VPWR net1029 sky130_fd_sc_hd__buf_6
XFILLER_75_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_39_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_16
XU$$2108 t$5482 net1442 VGND VGND VPWR VPWR booth_b30_m23 sky130_fd_sc_hd__xor2_1
XFILLER_90_717 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2119 net1050 net581 net1042 net854 VGND VGND VPWR VPWR t$5488 sky130_fd_sc_hd__a22o_1
XU$$1407 t$5124 net1488 VGND VGND VPWR VPWR booth_b20_m15 sky130_fd_sc_hd__xor2_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1418 net1114 net627 net1105 net900 VGND VGND VPWR VPWR t$5130 sky130_fd_sc_hd__a22o_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1429 t$5135 net1486 VGND VGND VPWR VPWR booth_b20_m26 sky130_fd_sc_hd__xor2_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_90_1 c$1798 c$1800 c$1802 VGND VGND VPWR VPWR c$2560 s$2561 sky130_fd_sc_hd__fa_1
XFILLER_183_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_83_0 s$951 c$1710 c$1712 VGND VGND VPWR VPWR c$2502 s$2503 sky130_fd_sc_hd__fa_1
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1530 net124 VGND VGND VPWR VPWR net1530 sky130_fd_sc_hd__buf_4
Xfanout1541 net1542 VGND VGND VPWR VPWR net1541 sky130_fd_sc_hd__clkbuf_4
XU$$4000 t$6449 net1287 VGND VGND VPWR VPWR booth_b58_m10 sky130_fd_sc_hd__xor2_1
Xfanout1552 net1559 VGND VGND VPWR VPWR net1552 sky130_fd_sc_hd__clkbuf_4
X_2170_ clknet_leaf_28_clk booth_b38_m22 VGND VGND VPWR VPWR pp_row60_19 sky130_fd_sc_hd__dfxtp_1
XU$$4011 net1168 net451 net1159 net724 VGND VGND VPWR VPWR t$6455 sky130_fd_sc_hd__a22o_1
Xfanout1563 net120 VGND VGND VPWR VPWR net1563 sky130_fd_sc_hd__clkbuf_8
XU$$4022 t$6460 net1286 VGND VGND VPWR VPWR booth_b58_m21 sky130_fd_sc_hd__xor2_1
Xfanout1574 net1575 VGND VGND VPWR VPWR net1574 sky130_fd_sc_hd__buf_4
Xfanout1585 net119 VGND VGND VPWR VPWR net1585 sky130_fd_sc_hd__buf_4
XU$$4033 net1069 net454 net1061 net727 VGND VGND VPWR VPWR t$6466 sky130_fd_sc_hd__a22o_1
X_1121_ clknet_leaf_48_clk booth_b14_m1 VGND VGND VPWR VPWR pp_row15_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_93_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1596 net1598 VGND VGND VPWR VPWR net1596 sky130_fd_sc_hd__buf_2
XU$$4044 t$6471 net1288 VGND VGND VPWR VPWR booth_b58_m32 sky130_fd_sc_hd__xor2_1
XU$$4055 net962 net455 net953 net728 VGND VGND VPWR VPWR t$6477 sky130_fd_sc_hd__a22o_1
XU$$3310 net1517 net500 net1510 net773 VGND VGND VPWR VPWR t$6097 sky130_fd_sc_hd__a22o_1
XU$$4066 t$6482 net1289 VGND VGND VPWR VPWR booth_b58_m43 sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_112_0 pp_row112_8 pp_row112_9 pp_row112_10 VGND VGND VPWR VPWR c$3362
+ s$3363 sky130_fd_sc_hd__fa_2
XFILLER_20_1012 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3321 t$6102 net1338 VGND VGND VPWR VPWR booth_b48_m13 sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_45_5 s$281 s$283 s$285 VGND VGND VPWR VPWR c$1276 s$1277 sky130_fd_sc_hd__fa_1
XU$$3332 net1145 net497 net1137 net770 VGND VGND VPWR VPWR t$6108 sky130_fd_sc_hd__a22o_1
XU$$4077 net1692 net453 net1685 net726 VGND VGND VPWR VPWR t$6488 sky130_fd_sc_hd__a22o_1
XU$$3343 t$6113 net1338 VGND VGND VPWR VPWR booth_b48_m24 sky130_fd_sc_hd__xor2_1
X_1052_ clknet_leaf_53_clk booth_b0_m8 VGND VGND VPWR VPWR pp_row8_0 sky130_fd_sc_hd__dfxtp_1
XU$$4088 t$6493 net1288 VGND VGND VPWR VPWR booth_b58_m54 sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_38_4 pp_row38_20 pp_row38_21 c$212 VGND VGND VPWR VPWR c$1190 s$1191 sky130_fd_sc_hd__fa_1
XU$$3354 net1043 net494 net1027 net767 VGND VGND VPWR VPWR t$6119 sky130_fd_sc_hd__a22o_1
XU$$4099 net1584 net459 net1557 net732 VGND VGND VPWR VPWR t$6499 sky130_fd_sc_hd__a22o_1
XU$$3365 t$6124 net1341 VGND VGND VPWR VPWR booth_b48_m35 sky130_fd_sc_hd__xor2_1
XU$$2620 t$5744 net1394 VGND VGND VPWR VPWR booth_b38_m5 sky130_fd_sc_hd__xor2_1
XFILLER_62_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3376 net927 net495 net1748 net768 VGND VGND VPWR VPWR t$6130 sky130_fd_sc_hd__a22o_1
XU$$2631 net1222 net544 net1214 net817 VGND VGND VPWR VPWR t$5750 sky130_fd_sc_hd__a22o_1
XU$$2642 t$5755 net1399 VGND VGND VPWR VPWR booth_b38_m16 sky130_fd_sc_hd__xor2_1
XU$$3387 t$6135 net1344 VGND VGND VPWR VPWR booth_b48_m46 sky130_fd_sc_hd__xor2_1
XFILLER_46_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2653 net1107 net550 net1098 net823 VGND VGND VPWR VPWR t$5761 sky130_fd_sc_hd__a22o_1
XU$$3398 net1652 net498 net1644 net771 VGND VGND VPWR VPWR t$6141 sky130_fd_sc_hd__a22o_1
XU$$2664 t$5766 net1399 VGND VGND VPWR VPWR booth_b38_m27 sky130_fd_sc_hd__xor2_1
XU$$1930 net1031 net584 net932 net857 VGND VGND VPWR VPWR t$5392 sky130_fd_sc_hd__a22o_1
XFILLER_55_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2675 net1002 net546 net994 net819 VGND VGND VPWR VPWR t$5772 sky130_fd_sc_hd__a22o_1
XU$$2686 t$5777 net1396 VGND VGND VPWR VPWR booth_b38_m38 sky130_fd_sc_hd__xor2_1
XU$$1941 t$5397 net1451 VGND VGND VPWR VPWR booth_b28_m8 sky130_fd_sc_hd__xor2_1
XU$$2697 net1731 net546 net1722 net819 VGND VGND VPWR VPWR t$5783 sky130_fd_sc_hd__a22o_1
XU$$1952 net1192 net584 net1173 net857 VGND VGND VPWR VPWR t$5403 sky130_fd_sc_hd__a22o_1
XFILLER_21_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1963 t$5408 net1450 VGND VGND VPWR VPWR booth_b28_m19 sky130_fd_sc_hd__xor2_1
XU$$1974 net1083 net587 net1074 net860 VGND VGND VPWR VPWR t$5414 sky130_fd_sc_hd__a22o_1
XU$$1985 t$5419 net1452 VGND VGND VPWR VPWR booth_b28_m30 sky130_fd_sc_hd__xor2_1
XU$$1996 net977 net588 net969 net861 VGND VGND VPWR VPWR t$5425 sky130_fd_sc_hd__a22o_1
X_1954_ clknet_leaf_66_clk booth_b12_m42 VGND VGND VPWR VPWR pp_row54_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_187_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0905_ clknet_leaf_103_clk booth_b38_m58 VGND VGND VPWR VPWR pp_row96_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_147_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1885_ clknet_leaf_78_clk booth_b2_m50 VGND VGND VPWR VPWR pp_row52_1 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_98_0 c$3272 c$3274 c$3276 VGND VGND VPWR VPWR c$3788 s$3789 sky130_fd_sc_hd__fa_1
XFILLER_174_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0836_ clknet_leaf_106_clk booth_b64_m28 VGND VGND VPWR VPWR pp_row92_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0767_ clknet_leaf_152_clk booth_b64_m25 VGND VGND VPWR VPWR pp_row89_20 sky130_fd_sc_hd__dfxtp_1
XFILLER_88_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0698_ clknet_leaf_174_clk booth_b30_m57 VGND VGND VPWR VPWR pp_row87_4 sky130_fd_sc_hd__dfxtp_1
X_2437_ clknet_leaf_74_clk booth_b52_m15 VGND VGND VPWR VPWR pp_row67_26 sky130_fd_sc_hd__dfxtp_1
XFILLER_5_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$604 final_adder.p_new$616 final_adder.p_new$608 VGND VGND VPWR VPWR
+ final_adder.p_new$732 sky130_fd_sc_hd__and2_2
X_2368_ clknet_leaf_98_clk booth_b64_m1 VGND VGND VPWR VPWR pp_row65_32 sky130_fd_sc_hd__dfxtp_1
XFILLER_99_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$615 final_adder.p_new$618 final_adder.g_new$627 final_adder.g_new$619
+ VGND VGND VPWR VPWR final_adder.g_new$743 sky130_fd_sc_hd__a21o_1
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$637 final_adder.p_new$644 final_adder.g_new$661 final_adder.g_new$645
+ VGND VGND VPWR VPWR final_adder.g_new$765 sky130_fd_sc_hd__a21o_1
XTAP_3919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$648 final_adder.p_new$672 final_adder.p_new$656 VGND VGND VPWR VPWR
+ final_adder.p_new$776 sky130_fd_sc_hd__and2_1
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1319_ clknet_leaf_250_clk booth_b6_m23 VGND VGND VPWR VPWR pp_row29_3 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$659 final_adder.p_new$666 final_adder.g_new$683 final_adder.g_new$667
+ VGND VGND VPWR VPWR final_adder.g_new$787 sky130_fd_sc_hd__a21o_1
X_2299_ clknet_leaf_199_clk booth_b4_m60 VGND VGND VPWR VPWR pp_row64_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_186_1016 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$509 net1716 net430 net1707 net712 VGND VGND VPWR VPWR t$4665 sky130_fd_sc_hd__a22o_1
XFILLER_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$70 net1016 net442 net999 net684 VGND VGND VPWR VPWR t$4442 sky130_fd_sc_hd__a22o_1
XU$$81 t$4447 net1568 VGND VGND VPWR VPWR booth_b0_m37 sky130_fd_sc_hd__xor2_1
XFILLER_71_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$92 net1737 net444 net1729 net686 VGND VGND VPWR VPWR t$4453 sky130_fd_sc_hd__a22o_1
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_1090 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_50 net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_61 net402 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 net441 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_83 net509 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_94 net534 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_107_1 pp_row107_6 pp_row107_7 pp_row107_8 VGND VGND VPWR VPWR c$2696 s$2697
+ sky130_fd_sc_hd__fa_1
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_48_3 s$1307 s$1309 s$1311 VGND VGND VPWR VPWR c$2228 s$2229 sky130_fd_sc_hd__fa_1
XFILLER_101_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1204 net1657 net650 net1649 net923 VGND VGND VPWR VPWR t$5020 sky130_fd_sc_hd__a22o_1
XU$$1215 t$5025 net1012 VGND VGND VPWR VPWR booth_b16_m56 sky130_fd_sc_hd__xor2_1
XFILLER_188_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1226 net1546 net648 net1538 net921 VGND VGND VPWR VPWR t$5031 sky130_fd_sc_hd__a22o_1
XU$$1237 notblock$5035\[2\] net10 net1013 t$5036 notblock$5035\[0\] VGND VGND VPWR
+ VPWR sel_0$5037 sky130_fd_sc_hd__a32o_2
XFILLER_71_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1248 t$5043 net1664 VGND VGND VPWR VPWR booth_b18_m4 sky130_fd_sc_hd__xor2_1
Xclkbuf_5_0__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_5_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_16_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1259 net1494 net635 net1219 net908 VGND VGND VPWR VPWR t$5049 sky130_fd_sc_hd__a22o_1
XFILLER_188_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$1020 final_adder.$signal$1149 final_adder.g_new$1060 VGND VGND VPWR
+ VPWR net339 sky130_fd_sc_hd__xor2_2
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1031 final_adder.$signal$1160 final_adder.g_new$1021 VGND VGND VPWR
+ VPWR net352 sky130_fd_sc_hd__xor2_2
X_1670_ clknet_leaf_19_clk booth_b32_m12 VGND VGND VPWR VPWR pp_row44_16 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$1042 final_adder.$signal$1171 final_adder.g_new$1049 VGND VGND VPWR
+ VPWR net364 sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$1053 final_adder.$signal$1182 final_adder.g_new$999 VGND VGND VPWR
+ VPWR net376 sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$1064 final_adder.$signal$1193 final_adder.g_new$1038 VGND VGND VPWR
+ VPWR net261 sky130_fd_sc_hd__xor2_1
XFILLER_172_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$1075 final_adder.$signal$1204 final_adder.g_new$977 VGND VGND VPWR
+ VPWR net273 sky130_fd_sc_hd__xor2_2
X_0621_ clknet_leaf_187_clk booth_b30_m54 VGND VGND VPWR VPWR pp_row84_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1086 final_adder.$signal$1215 final_adder.g_new$1027 VGND VGND VPWR
+ VPWR net285 sky130_fd_sc_hd__xor2_2
X_0552_ clknet_leaf_171_clk booth_b54_m27 VGND VGND VPWR VPWR pp_row81_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_125_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0483_ clknet_leaf_156_clk booth_b34_m45 VGND VGND VPWR VPWR pp_row79_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_98_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2222_ clknet_leaf_229_clk booth_b0_m62 VGND VGND VPWR VPWR pp_row62_0 sky130_fd_sc_hd__dfxtp_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_991 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1360 net1361 VGND VGND VPWR VPWR net1360 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_50_3 c$346 s$349 s$351 VGND VGND VPWR VPWR c$1332 s$1333 sky130_fd_sc_hd__fa_2
Xfanout1371 net38 VGND VGND VPWR VPWR net1371 sky130_fd_sc_hd__buf_6
XFILLER_66_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1382 net1383 VGND VGND VPWR VPWR net1382 sky130_fd_sc_hd__buf_6
X_2153_ clknet_leaf_214_clk booth_b6_m54 VGND VGND VPWR VPWR pp_row60_3 sky130_fd_sc_hd__dfxtp_1
Xfanout1393 net34 VGND VGND VPWR VPWR net1393 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_43_2 pp_row43_20 pp_row43_21 pp_row43_22 VGND VGND VPWR VPWR c$1246 s$1247
+ sky130_fd_sc_hd__fa_1
X_1104_ clknet_leaf_13_clk booth_b4_m10 VGND VGND VPWR VPWR pp_row14_2 sky130_fd_sc_hd__dfxtp_1
XU$$3140 net1585 net515 net1558 net788 VGND VGND VPWR VPWR t$6009 sky130_fd_sc_hd__a22o_1
XFILLER_81_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2084_ clknet_leaf_31_clk booth_b6_m52 VGND VGND VPWR VPWR pp_row58_3 sky130_fd_sc_hd__dfxtp_1
XU$$3151 net1361 VGND VGND VPWR VPWR notblock$6015\[0\] sky130_fd_sc_hd__inv_1
Xdadda_fa_5_20_1 s$2811 s$2813 s$2815 VGND VGND VPWR VPWR c$3478 s$3479 sky130_fd_sc_hd__fa_1
XU$$3162 t$6021 net1348 VGND VGND VPWR VPWR booth_b46_m2 sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_36_1 pp_row36_8 pp_row36_9 pp_row36_10 VGND VGND VPWR VPWR c$1160 s$1161
+ sky130_fd_sc_hd__fa_1
XU$$3173 net1517 net505 net1510 net778 VGND VGND VPWR VPWR t$6027 sky130_fd_sc_hd__a22o_1
X_1035_ clknet_leaf_61_clk booth_b0_m5 VGND VGND VPWR VPWR pp_row5_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_81_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3184 t$6032 net1348 VGND VGND VPWR VPWR booth_b46_m13 sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_13_0 c$2762 c$2764 c$2766 VGND VGND VPWR VPWR c$3448 s$3449 sky130_fd_sc_hd__fa_1
XU$$3195 net1145 net505 net1137 net778 VGND VGND VPWR VPWR t$6038 sky130_fd_sc_hd__a22o_1
XFILLER_62_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2450 t$5656 net1428 VGND VGND VPWR VPWR booth_b34_m57 sky130_fd_sc_hd__xor2_1
XU$$2461 net1542 net567 net1534 net840 VGND VGND VPWR VPWR t$5662 sky130_fd_sc_hd__a22o_1
XU$$1504_1762 VGND VGND VPWR VPWR U$$1504_1762/HI net1762 sky130_fd_sc_hd__conb_1
Xdadda_fa_2_29_0 pp_row29_0 pp_row29_1 pp_row29_2 VGND VGND VPWR VPWR c$1082 s$1083
+ sky130_fd_sc_hd__fa_1
XU$$2472 net1777 net554 net1232 net827 VGND VGND VPWR VPWR t$5669 sky130_fd_sc_hd__a22o_1
XFILLER_34_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2483 t$5674 net1403 VGND VGND VPWR VPWR booth_b36_m5 sky130_fd_sc_hd__xor2_1
XFILLER_61_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2494 net1220 net551 net1213 net824 VGND VGND VPWR VPWR t$5680 sky130_fd_sc_hd__a22o_1
XFILLER_107_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1760 net1622 net608 net1613 net881 VGND VGND VPWR VPWR t$5304 sky130_fd_sc_hd__a22o_1
XFILLER_167_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1771 t$5309 net1471 VGND VGND VPWR VPWR booth_b24_m60 sky130_fd_sc_hd__xor2_1
XU$$1782 net19 VGND VGND VPWR VPWR notblock$5315\[1\] sky130_fd_sc_hd__inv_1
XU$$1793 net1031 net593 net932 net866 VGND VGND VPWR VPWR t$5322 sky130_fd_sc_hd__a22o_1
XFILLER_148_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1937_ clknet_leaf_70_clk booth_b40_m13 VGND VGND VPWR VPWR pp_row53_20 sky130_fd_sc_hd__dfxtp_1
XFILLER_30_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1868_ clknet_leaf_66_clk booth_b26_m25 VGND VGND VPWR VPWR pp_row51_13 sky130_fd_sc_hd__dfxtp_1
Xinput70 b[14] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_2
XFILLER_174_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0819_ clknet_leaf_111_clk booth_b36_m56 VGND VGND VPWR VPWR pp_row92_5 sky130_fd_sc_hd__dfxtp_1
Xinput81 b[24] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__buf_6
Xinput92 b[34] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_4
X_1799_ clknet_leaf_220_clk booth_b10_m39 VGND VGND VPWR VPWR pp_row49_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_58_2 s$2305 s$2307 s$2309 VGND VGND VPWR VPWR c$3042 s$3043 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$401 final_adder.p_new$402 final_adder.g_new$407 final_adder.g_new$403
+ VGND VGND VPWR VPWR final_adder.g_new$529 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$412 final_adder.p_new$418 final_adder.p_new$414 VGND VGND VPWR VPWR
+ final_adder.p_new$540 sky130_fd_sc_hd__and2_1
XFILLER_29_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$423 final_adder.p_new$424 final_adder.g_new$429 final_adder.g_new$425
+ VGND VGND VPWR VPWR final_adder.g_new$551 sky130_fd_sc_hd__a21o_1
XTAP_3705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$434 final_adder.p_new$440 final_adder.p_new$436 VGND VGND VPWR VPWR
+ final_adder.p_new$562 sky130_fd_sc_hd__and2_1
XTAP_3716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$445 final_adder.p_new$446 final_adder.g_new$451 final_adder.g_new$447
+ VGND VGND VPWR VPWR final_adder.g_new$573 sky130_fd_sc_hd__a21o_1
XFILLER_29_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_28_0 s$3511 c$3950 s$3953 VGND VGND VPWR VPWR c$4208 s$4209 sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$456 final_adder.p_new$462 final_adder.p_new$458 VGND VGND VPWR VPWR
+ final_adder.p_new$584 sky130_fd_sc_hd__and2_1
XTAP_3738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$306 net1203 net528 net1194 net801 VGND VGND VPWR VPWR t$4562 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$467 final_adder.p_new$468 final_adder.g_new$473 final_adder.g_new$469
+ VGND VGND VPWR VPWR final_adder.g_new$595 sky130_fd_sc_hd__a21o_1
XTAP_3749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$317 t$4567 net1279 VGND VGND VPWR VPWR booth_b4_m18 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$478 final_adder.p_new$484 final_adder.p_new$480 VGND VGND VPWR VPWR
+ final_adder.p_new$606 sky130_fd_sc_hd__and2_1
XFILLER_45_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$328 net1088 net527 net1080 net800 VGND VGND VPWR VPWR t$4573 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$489 final_adder.p_new$490 final_adder.g_new$495 final_adder.g_new$491
+ VGND VGND VPWR VPWR final_adder.g_new$617 sky130_fd_sc_hd__a21o_1
XU$$339 t$4578 net1277 VGND VGND VPWR VPWR booth_b4_m29 sky130_fd_sc_hd__xor2_1
XFILLER_72_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_60_2 c$1444 s$1447 s$1449 VGND VGND VPWR VPWR c$2322 s$2323 sky130_fd_sc_hd__fa_1
XFILLER_110_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_53_1 c$1354 c$1356 c$1358 VGND VGND VPWR VPWR c$2264 s$2265 sky130_fd_sc_hd__fa_1
XFILLER_88_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_0_69_1 pp_row69_3 pp_row69_4 pp_row69_5 VGND VGND VPWR VPWR c$146 s$147
+ sky130_fd_sc_hd__fa_1
Xdadda_fa_6_30_0 c$3512 c$3514 s$3517 VGND VGND VPWR VPWR c$3956 s$3957 sky130_fd_sc_hd__fa_1
XFILLER_48_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_46_0 s$301 c$1266 c$1268 VGND VGND VPWR VPWR c$2206 s$2207 sky130_fd_sc_hd__fa_1
XFILLER_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$990 final_adder.$signal$1119 final_adder.g_new$1075 VGND VGND VPWR
+ VPWR net306 sky130_fd_sc_hd__xor2_2
XU$$840 net1561 net396 net1522 net662 VGND VGND VPWR VPWR t$4835 sky130_fd_sc_hd__a22o_1
XFILLER_63_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$851 t$4840 net1312 VGND VGND VPWR VPWR booth_b12_m11 sky130_fd_sc_hd__xor2_1
XU$$862 net1155 net393 net1146 net659 VGND VGND VPWR VPWR t$4846 sky130_fd_sc_hd__a22o_1
XU$$1001 net1149 net388 net1143 net654 VGND VGND VPWR VPWR t$4917 sky130_fd_sc_hd__a22o_1
XU$$1012 t$4922 net1186 VGND VGND VPWR VPWR booth_b14_m23 sky130_fd_sc_hd__xor2_1
XU$$873 t$4851 net1313 VGND VGND VPWR VPWR booth_b12_m22 sky130_fd_sc_hd__xor2_1
XU$$1023 net1047 net386 net1039 net652 VGND VGND VPWR VPWR t$4928 sky130_fd_sc_hd__a22o_1
XU$$884 net1055 net394 net1047 net660 VGND VGND VPWR VPWR t$4857 sky130_fd_sc_hd__a22o_1
XFILLER_188_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1034 t$4933 net1184 VGND VGND VPWR VPWR booth_b14_m34 sky130_fd_sc_hd__xor2_1
XU$$895 t$4862 net1314 VGND VGND VPWR VPWR booth_b12_m33 sky130_fd_sc_hd__xor2_1
XFILLER_16_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1045 net944 net388 net928 net654 VGND VGND VPWR VPWR t$4939 sky130_fd_sc_hd__a22o_1
XU$$1056 t$4944 net1190 VGND VGND VPWR VPWR booth_b14_m45 sky130_fd_sc_hd__xor2_1
XFILLER_189_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1067 net1657 net391 net1649 net657 VGND VGND VPWR VPWR t$4950 sky130_fd_sc_hd__a22o_1
XFILLER_188_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1078 t$4955 net1191 VGND VGND VPWR VPWR booth_b14_m56 sky130_fd_sc_hd__xor2_1
XFILLER_189_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1089 net1543 net391 net1535 net657 VGND VGND VPWR VPWR t$4961 sky130_fd_sc_hd__a22o_1
XFILLER_89_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1722_ clknet_leaf_22_clk booth_b28_m18 VGND VGND VPWR VPWR pp_row46_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_117_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_103_0 s$3811 c$4100 s$4103 VGND VGND VPWR VPWR c$4358 s$4359 sky130_fd_sc_hd__fa_1
XFILLER_145_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1653_ clknet_leaf_221_clk booth_b0_m44 VGND VGND VPWR VPWR pp_row44_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_98_3 pp_row98_9 pp_row98_10 pp_row98_11 VGND VGND VPWR VPWR c$1908 s$1909
+ sky130_fd_sc_hd__fa_1
XU$$3979_1801 VGND VGND VPWR VPWR U$$3979_1801/HI net1801 sky130_fd_sc_hd__conb_1
X_0604_ clknet_leaf_174_clk booth_b48_m35 VGND VGND VPWR VPWR pp_row83_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_113_700 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1584_ clknet_leaf_243_clk booth_b14_m27 VGND VGND VPWR VPWR pp_row41_7 sky130_fd_sc_hd__dfxtp_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout608 net609 VGND VGND VPWR VPWR net608 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_5_68_1 s$3099 s$3101 s$3103 VGND VGND VPWR VPWR c$3670 s$3671 sky130_fd_sc_hd__fa_1
XFILLER_152_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0535_ clknet_leaf_166_clk booth_b22_m59 VGND VGND VPWR VPWR pp_row81_3 sky130_fd_sc_hd__dfxtp_1
Xfanout619 net622 VGND VGND VPWR VPWR net619 sky130_fd_sc_hd__buf_4
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0466_ clknet_leaf_130_clk booth_b56_m59 VGND VGND VPWR VPWR pp_row115_3 sky130_fd_sc_hd__dfxtp_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2205_ clknet_leaf_133_clk booth_b46_m64 VGND VGND VPWR VPWR pp_row110_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0397_ clknet_leaf_191_clk booth_b42_m34 VGND VGND VPWR VPWR pp_row76_16 sky130_fd_sc_hd__dfxtp_1
Xfanout1190 net1191 VGND VGND VPWR VPWR net1190 sky130_fd_sc_hd__buf_4
XFILLER_113_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2136_ clknet_leaf_27_clk booth_b38_m21 VGND VGND VPWR VPWR pp_row59_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_96_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2067_ clknet_leaf_35_clk booth_b36_m21 VGND VGND VPWR VPWR pp_row57_18 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_107_0 pp_row107_0 pp_row107_1 pp_row107_2 VGND VGND VPWR VPWR c$1970 s$1971
+ sky130_fd_sc_hd__fa_1
X_1018_ clknet_leaf_60_clk net1574 VGND VGND VPWR VPWR pp_row0_1 sky130_fd_sc_hd__dfxtp_4
XU$$2280 net925 net570 net1746 net843 VGND VGND VPWR VPWR t$5570 sky130_fd_sc_hd__a22o_1
XU$$2291 t$5575 net1435 VGND VGND VPWR VPWR booth_b32_m46 sky130_fd_sc_hd__xor2_1
XFILLER_22_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1590 t$5217 net1477 VGND VGND VPWR VPWR booth_b22_m38 sky130_fd_sc_hd__xor2_1
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_70_1 c$2394 c$2396 s$2399 VGND VGND VPWR VPWR c$3112 s$3113 sky130_fd_sc_hd__fa_1
XFILLER_150_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_86_1 pp_row86_3 pp_row86_4 pp_row86_5 VGND VGND VPWR VPWR c$980 s$981
+ sky130_fd_sc_hd__fa_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_63_0 s$1493 c$2334 c$2336 VGND VGND VPWR VPWR c$3068 s$3069 sky130_fd_sc_hd__fa_1
Xdadda_fa_1_79_0 pp_row79_0 pp_row79_1 pp_row79_2 VGND VGND VPWR VPWR c$870 s$871
+ sky130_fd_sc_hd__fa_1
XTAP_4203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$220 final_adder.$signal$1124 final_adder.$signal$1125 VGND VGND VPWR
+ VPWR final_adder.p_new$348 sky130_fd_sc_hd__and2_1
XTAP_4247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$231 final_adder.$signal$1115 final_adder.$signal$50 final_adder.$signal$52
+ VGND VGND VPWR VPWR final_adder.g_new$359 sky130_fd_sc_hd__a21o_1
XTAP_3513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3909 t$6402 net1293 VGND VGND VPWR VPWR booth_b56_m33 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$242 final_adder.$signal$1102 final_adder.$signal$1103 VGND VGND VPWR
+ VPWR final_adder.p_new$370 sky130_fd_sc_hd__and2_1
XTAP_4258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$253 final_adder.$signal$1093 final_adder.$signal$6 final_adder.$signal$8
+ VGND VGND VPWR VPWR final_adder.g_new$381 sky130_fd_sc_hd__a21o_1
XTAP_3524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$103 t$4458 net1570 VGND VGND VPWR VPWR booth_b0_m48 sky130_fd_sc_hd__xor2_1
XFILLER_40_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$264 final_adder.p_new$266 final_adder.p_new$264 VGND VGND VPWR VPWR
+ final_adder.p_new$392 sky130_fd_sc_hd__and2_1
XFILLER_175_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$114 net1633 net449 net1623 net691 VGND VGND VPWR VPWR t$4464 sky130_fd_sc_hd__a22o_1
XTAP_3546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$275 final_adder.p_new$274 final_adder.g_new$277 final_adder.g_new$275
+ VGND VGND VPWR VPWR final_adder.g_new$403 sky130_fd_sc_hd__a21o_1
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$286 final_adder.p_new$288 final_adder.p_new$286 VGND VGND VPWR VPWR
+ final_adder.p_new$414 sky130_fd_sc_hd__and2_1
XU$$125 t$4469 net1572 VGND VGND VPWR VPWR booth_b0_m59 sky130_fd_sc_hd__xor2_1
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$136 net1577 VGND VGND VPWR VPWR notsign sky130_fd_sc_hd__inv_1
Xfinal_adder.U$$297 final_adder.p_new$296 final_adder.g_new$299 final_adder.g_new$297
+ VGND VGND VPWR VPWR final_adder.g_new$425 sky130_fd_sc_hd__a21o_1
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$147 net1127 net624 net1035 net897 VGND VGND VPWR VPWR t$4481 sky130_fd_sc_hd__a22o_1
XTAP_3579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$158 t$4486 net1390 VGND VGND VPWR VPWR booth_b2_m7 sky130_fd_sc_hd__xor2_1
XU$$169 net1203 net620 net1194 net893 VGND VGND VPWR VPWR t$4492 sky130_fd_sc_hd__a22o_1
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4395_1818 VGND VGND VPWR VPWR U$$4395_1818/HI net1818 sky130_fd_sc_hd__conb_1
XFILLER_12_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_78_0 c$3704 c$3706 s$3709 VGND VGND VPWR VPWR c$4052 s$4053 sky130_fd_sc_hd__fa_1
XFILLER_57_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_243_clk clknet_5_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_243_clk
+ sky130_fd_sc_hd__clkbuf_16
X_0320_ clknet_leaf_200_clk booth_b18_m56 VGND VGND VPWR VPWR pp_row74_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_96_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0251_ clknet_leaf_210_clk booth_b12_m60 VGND VGND VPWR VPWR pp_row72_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_48_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0182_ clknet_leaf_147_clk booth_b8_m62 VGND VGND VPWR VPWR pp_row70_2 sky130_fd_sc_hd__dfxtp_1
XU$$670 net1599 net416 net1590 net682 VGND VGND VPWR VPWR t$4747 sky130_fd_sc_hd__a22o_1
XU$$681 t$4752 net1237 VGND VGND VPWR VPWR booth_b8_m63 sky130_fd_sc_hd__xor2_1
XFILLER_189_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$692 t$4759 net1414 VGND VGND VPWR VPWR booth_b10_m0 sky130_fd_sc_hd__xor2_1
XFILLER_16_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1705_ clknet_leaf_123_clk booth_b52_m54 VGND VGND VPWR VPWR pp_row106_6 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_80_0 c$3164 c$3166 c$3168 VGND VGND VPWR VPWR c$3716 s$3717 sky130_fd_sc_hd__fa_1
Xdadda_fa_2_96_0 pp_row96_2 pp_row96_3 pp_row96_4 VGND VGND VPWR VPWR c$1878 s$1879
+ sky130_fd_sc_hd__fa_1
XFILLER_172_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1636_ clknet_leaf_223_clk booth_b16_m27 VGND VGND VPWR VPWR pp_row43_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_99_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1567_ clknet_leaf_7_clk booth_b30_m10 VGND VGND VPWR VPWR pp_row40_15 sky130_fd_sc_hd__dfxtp_1
Xfanout405 net406 VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__buf_2
XFILLER_87_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout416 net417 VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_234_clk clknet_5_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_234_clk
+ sky130_fd_sc_hd__clkbuf_16
Xfanout427 net428 VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__buf_6
XFILLER_59_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_72_7 c$166 c$168 c$170 VGND VGND VPWR VPWR c$758 s$759 sky130_fd_sc_hd__fa_1
XFILLER_113_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout438 net441 VGND VGND VPWR VPWR net438 sky130_fd_sc_hd__clkbuf_4
X_0518_ clknet_leaf_166_clk booth_b44_m36 VGND VGND VPWR VPWR pp_row80_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_140_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout449 net450 VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__buf_6
XFILLER_100_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1498_ clknet_leaf_45_clk booth_b32_m5 VGND VGND VPWR VPWR pp_row37_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_58_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_65_6 c$88 c$90 c$92 VGND VGND VPWR VPWR c$630 s$631 sky130_fd_sc_hd__fa_1
X_0449_ clknet_leaf_206_clk booth_b26_m52 VGND VGND VPWR VPWR pp_row78_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_55_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_58_5 pp_row58_26 pp_row58_27 pp_row58_28 VGND VGND VPWR VPWR c$502 s$503
+ sky130_fd_sc_hd__fa_1
XFILLER_55_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2119_ clknet_leaf_218_clk booth_b6_m53 VGND VGND VPWR VPWR pp_row59_3 sky130_fd_sc_hd__dfxtp_1
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_580 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_95_0 s$3779 c$4084 s$4087 VGND VGND VPWR VPWR c$4342 s$4343 sky130_fd_sc_hd__fa_1
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_225_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_225_clk
+ sky130_fd_sc_hd__clkbuf_16
Xfanout950 net952 VGND VGND VPWR VPWR net950 sky130_fd_sc_hd__buf_6
XFILLER_131_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4407 t$6657 net1824 VGND VGND VPWR VPWR booth_b64_m8 sky130_fd_sc_hd__xor2_1
Xfanout961 net963 VGND VGND VPWR VPWR net961 sky130_fd_sc_hd__buf_4
Xfanout972 net94 VGND VGND VPWR VPWR net972 sky130_fd_sc_hd__buf_6
XTAP_4011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4418 net1196 sel_0$6647 net1177 net694 VGND VGND VPWR VPWR t$6663 sky130_fd_sc_hd__a22o_1
XU$$4429 t$6668 net1835 VGND VGND VPWR VPWR booth_b64_m19 sky130_fd_sc_hd__xor2_1
Xfanout983 net986 VGND VGND VPWR VPWR net983 sky130_fd_sc_hd__buf_6
XTAP_4033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout994 net997 VGND VGND VPWR VPWR net994 sky130_fd_sc_hd__buf_6
Xdadda_fa_6_110_0 c$3832 c$3834 s$3837 VGND VGND VPWR VPWR c$4116 s$4117 sky130_fd_sc_hd__fa_1
XTAP_4044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3706 t$6299 net1304 VGND VGND VPWR VPWR booth_b54_m0 sky130_fd_sc_hd__xor2_1
XFILLER_18_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3717 net1563 net468 net1522 net741 VGND VGND VPWR VPWR t$6305 sky130_fd_sc_hd__a22o_1
XTAP_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3728 t$6310 net1304 VGND VGND VPWR VPWR booth_b54_m11 sky130_fd_sc_hd__xor2_1
XTAP_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3739 net1160 net470 net1151 net743 VGND VGND VPWR VPWR t$6316 sky130_fd_sc_hd__a22o_1
XTAP_4088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_30_3 s$1093 s$1095 s$1097 VGND VGND VPWR VPWR c$2084 s$2085 sky130_fd_sc_hd__fa_1
XTAP_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_310 net479 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_321 net622 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_332 net712 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdadda_fa_3_23_2 pp_row23_8 pp_row23_9 pp_row23_10 VGND VGND VPWR VPWR c$2026 s$2027
+ sky130_fd_sc_hd__fa_1
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_343 net841 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_354 net931 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_365 net1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_376 net1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_387 net1507 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_398 net1627 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1072 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2470_ clknet_leaf_98_clk booth_b48_m20 VGND VGND VPWR VPWR pp_row68_23 sky130_fd_sc_hd__dfxtp_1
XFILLER_154_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1421_ clknet_leaf_54_clk booth_b12_m22 VGND VGND VPWR VPWR pp_row34_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_69_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_75_5 s$809 s$811 s$813 VGND VGND VPWR VPWR c$1636 s$1637 sky130_fd_sc_hd__fa_1
Xclkbuf_leaf_216_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_216_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_96_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1352_ clknet_leaf_244_clk net180 VGND VGND VPWR VPWR pp_row30_17 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_68_4 s$677 s$679 s$681 VGND VGND VPWR VPWR c$1550 s$1551 sky130_fd_sc_hd__fa_2
XFILLER_110_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0303_ clknet_leaf_227_clk booth_b44_m29 VGND VGND VPWR VPWR pp_row73_18 sky130_fd_sc_hd__dfxtp_1
X_1283_ clknet_leaf_181_clk net154 VGND VGND VPWR VPWR pp_row122_5 sky130_fd_sc_hd__dfxtp_2
XFILLER_37_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0234_ clknet_leaf_151_clk booth_b40_m31 VGND VGND VPWR VPWR pp_row71_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_1106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0998_ clknet_leaf_118_clk booth_b38_m63 VGND VGND VPWR VPWR pp_row101_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_146_931 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1102_1755 VGND VGND VPWR VPWR U$$1102_1755/HI net1755 sky130_fd_sc_hd__conb_1
XFILLER_192_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_105_1 s$3321 s$3323 s$3325 VGND VGND VPWR VPWR c$3818 s$3819 sky130_fd_sc_hd__fa_1
XFILLER_145_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1619_ clknet_leaf_240_clk booth_b32_m10 VGND VGND VPWR VPWR pp_row42_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_114_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_207_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_207_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_99_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_70_4 pp_row70_26 pp_row70_27 pp_row70_28 VGND VGND VPWR VPWR c$716 s$717
+ sky130_fd_sc_hd__fa_1
XFILLER_87_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_63_3 pp_row63_26 pp_row63_27 pp_row63_28 VGND VGND VPWR VPWR c$588 s$589
+ sky130_fd_sc_hd__fa_1
XFILLER_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_40_2 s$2161 s$2163 s$2165 VGND VGND VPWR VPWR c$2934 s$2935 sky130_fd_sc_hd__fa_1
XFILLER_101_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_56_2 pp_row56_14 pp_row56_15 pp_row56_16 VGND VGND VPWR VPWR c$460 s$461
+ sky130_fd_sc_hd__fa_1
XFILLER_83_940 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_33_1 c$2098 c$2100 s$2103 VGND VGND VPWR VPWR c$2890 s$2891 sky130_fd_sc_hd__fa_1
Xdadda_fa_1_49_1 pp_row49_3 pp_row49_4 pp_row49_5 VGND VGND VPWR VPWR c$334 s$335
+ sky130_fd_sc_hd__fa_1
Xdadda_fa_7_10_0 s$3439 c$3914 s$3917 VGND VGND VPWR VPWR c$4172 s$4173 sky130_fd_sc_hd__fa_1
XFILLER_131_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_26_0 s$1067 c$2038 c$2040 VGND VGND VPWR VPWR c$2846 s$2847 sky130_fd_sc_hd__fa_1
XFILLER_70_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1083 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_78_3 s$1667 s$1669 s$1671 VGND VGND VPWR VPWR c$2468 s$2469 sky130_fd_sc_hd__fa_1
XFILLER_151_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1701 net1702 VGND VGND VPWR VPWR net1701 sky130_fd_sc_hd__clkbuf_2
Xfanout1712 net1714 VGND VGND VPWR VPWR net1712 sky130_fd_sc_hd__clkbuf_4
Xfanout1723 net103 VGND VGND VPWR VPWR net1723 sky130_fd_sc_hd__buf_4
XFILLER_132_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1734 net1735 VGND VGND VPWR VPWR net1734 sky130_fd_sc_hd__buf_4
Xfanout1745 net1746 VGND VGND VPWR VPWR net1745 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4204 net1735 net440 net1727 net722 VGND VGND VPWR VPWR t$6553 sky130_fd_sc_hd__a22o_1
XFILLER_49_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4215 t$6558 net1267 VGND VGND VPWR VPWR booth_b60_m49 sky130_fd_sc_hd__xor2_1
XFILLER_172_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout780 net781 VGND VGND VPWR VPWR net780 sky130_fd_sc_hd__buf_4
XU$$4226 net1625 net439 net1617 net721 VGND VGND VPWR VPWR t$6564 sky130_fd_sc_hd__a22o_1
Xfanout791 sel_1$5948 VGND VGND VPWR VPWR net791 sky130_fd_sc_hd__buf_4
XFILLER_93_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4237 t$6569 net1265 VGND VGND VPWR VPWR booth_b60_m60 sky130_fd_sc_hd__xor2_1
XFILLER_18_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3503 net975 net485 net966 net758 VGND VGND VPWR VPWR t$6195 sky130_fd_sc_hd__a22o_1
Xdadda_ha_3_15_0 pp_row15_0 pp_row15_1 VGND VGND VPWR VPWR c$1976 s$1977 sky130_fd_sc_hd__ha_1
XU$$4248 net59 VGND VGND VPWR VPWR notblock$6575\[1\] sky130_fd_sc_hd__inv_1
XU$$4259 net1037 net422 net938 net704 VGND VGND VPWR VPWR t$6582 sky130_fd_sc_hd__a22o_1
XFILLER_168_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3514 t$6200 net1335 VGND VGND VPWR VPWR booth_b50_m41 sky130_fd_sc_hd__xor2_1
XU$$3525 net1708 net490 net1700 net763 VGND VGND VPWR VPWR t$6206 sky130_fd_sc_hd__a22o_1
XFILLER_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3536 t$6211 net1336 VGND VGND VPWR VPWR booth_b50_m52 sky130_fd_sc_hd__xor2_1
XU$$2802 net1062 net540 net1053 net813 VGND VGND VPWR VPWR t$5837 sky130_fd_sc_hd__a22o_1
XFILLER_65_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3547 net1600 net489 net1591 net762 VGND VGND VPWR VPWR t$6217 sky130_fd_sc_hd__a22o_1
XTAP_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2813 t$5842 net1377 VGND VGND VPWR VPWR booth_b40_m33 sky130_fd_sc_hd__xor2_1
XU$$1641_1764 VGND VGND VPWR VPWR U$$1641_1764/HI net1764 sky130_fd_sc_hd__conb_1
XU$$3558 t$6222 net1334 VGND VGND VPWR VPWR booth_b50_m63 sky130_fd_sc_hd__xor2_1
XTAP_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2824 net950 net537 net942 net810 VGND VGND VPWR VPWR t$5848 sky130_fd_sc_hd__a22o_1
XU$$3569 t$6229 net1319 VGND VGND VPWR VPWR booth_b52_m0 sky130_fd_sc_hd__xor2_1
XU$$2835 t$5853 net1378 VGND VGND VPWR VPWR booth_b40_m44 sky130_fd_sc_hd__xor2_1
XTAP_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2846 net1685 net541 net1659 net814 VGND VGND VPWR VPWR t$5859 sky130_fd_sc_hd__a22o_1
XTAP_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2857 t$5864 net1382 VGND VGND VPWR VPWR booth_b40_m55 sky130_fd_sc_hd__xor2_1
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_140 net760 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2868 net1558 net540 net1550 net813 VGND VGND VPWR VPWR t$5870 sky130_fd_sc_hd__a22o_1
XANTENNA_151 net799 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_162 net861 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2879 net1369 VGND VGND VPWR VPWR notblock$5875\[2\] sky130_fd_sc_hd__inv_1
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_173 net915 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_184 net968 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1970_ clknet_leaf_72_clk booth_b42_m12 VGND VGND VPWR VPWR pp_row54_21 sky130_fd_sc_hd__dfxtp_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_195 net1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0921_ clknet_leaf_181_clk net152 VGND VGND VPWR VPWR pp_row120_6 sky130_fd_sc_hd__dfxtp_2
XFILLER_147_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0852_ clknet_leaf_144_clk booth_b54_m39 VGND VGND VPWR VPWR pp_row93_13 sky130_fd_sc_hd__dfxtp_1
X_0783_ clknet_leaf_140_clk booth_b52_m38 VGND VGND VPWR VPWR pp_row90_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_170_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_80_3 c$886 s$889 s$891 VGND VGND VPWR VPWR c$1692 s$1693 sky130_fd_sc_hd__fa_1
X_2453_ clknet_leaf_92_clk booth_b18_m50 VGND VGND VPWR VPWR pp_row68_8 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_73_2 c$754 c$756 c$758 VGND VGND VPWR VPWR c$1606 s$1607 sky130_fd_sc_hd__fa_1
X_1404_ clknet_leaf_51_clk booth_b18_m15 VGND VGND VPWR VPWR pp_row33_9 sky130_fd_sc_hd__dfxtp_1
X_2384_ clknet_leaf_83_clk booth_b26_m40 VGND VGND VPWR VPWR pp_row66_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_69_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_50_1 s$2991 s$2993 s$2995 VGND VGND VPWR VPWR c$3598 s$3599 sky130_fd_sc_hd__fa_1
Xdadda_fa_2_66_1 c$622 c$624 c$626 VGND VGND VPWR VPWR c$1520 s$1521 sky130_fd_sc_hd__fa_2
XFILLER_110_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1335_ clknet_leaf_0_clk booth_b4_m26 VGND VGND VPWR VPWR pp_row30_2 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_43_0 c$2942 c$2944 c$2946 VGND VGND VPWR VPWR c$3568 s$3569 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$819 final_adder.p_new$834 final_adder.g_new$747 final_adder.g_new$835
+ VGND VGND VPWR VPWR final_adder.g_new$947 sky130_fd_sc_hd__a21o_1
Xdadda_fa_2_59_0 s$39 c$492 c$494 VGND VGND VPWR VPWR c$1434 s$1435 sky130_fd_sc_hd__fa_1
XFILLER_110_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput2 a[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_2
X_1266_ clknet_leaf_2_clk booth_b8_m18 VGND VGND VPWR VPWR pp_row26_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0217_ clknet_leaf_198_clk booth_b10_m61 VGND VGND VPWR VPWR pp_row71_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_65_973 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1197_ clknet_leaf_51_clk booth_b18_m3 VGND VGND VPWR VPWR pp_row21_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_188_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$0 pp_row0_2 s$4153 VGND VGND VPWR VPWR final_adder.$signal final_adder.$signal$1
+ sky130_fd_sc_hd__ha_1
XFILLER_192_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_88_2 s$2545 s$2547 s$2549 VGND VGND VPWR VPWR c$3222 s$3223 sky130_fd_sc_hd__fa_1
XFILLER_69_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_1024 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput350 net350 VGND VGND VPWR VPWR o[69] sky130_fd_sc_hd__buf_2
XFILLER_161_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput361 net361 VGND VGND VPWR VPWR o[79] sky130_fd_sc_hd__buf_2
Xdadda_fa_7_58_0 s$3631 c$4010 s$4013 VGND VGND VPWR VPWR c$4268 s$4269 sky130_fd_sc_hd__fa_1
XFILLER_133_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput372 net372 VGND VGND VPWR VPWR o[89] sky130_fd_sc_hd__buf_2
Xoutput383 net383 VGND VGND VPWR VPWR o[99] sky130_fd_sc_hd__buf_2
XFILLER_0_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1008 net1011 VGND VGND VPWR VPWR net1008 sky130_fd_sc_hd__buf_6
XFILLER_99_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1019 net1021 VGND VGND VPWR VPWR net1019 sky130_fd_sc_hd__buf_6
XFILLER_102_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_61_0 pp_row61_14 pp_row61_15 pp_row61_16 VGND VGND VPWR VPWR c$546 s$547
+ sky130_fd_sc_hd__fa_2
XFILLER_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2109 net1092 net580 net1083 net853 VGND VGND VPWR VPWR t$5483 sky130_fd_sc_hd__a22o_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1408 net1170 net629 net1161 net902 VGND VGND VPWR VPWR t$5125 sky130_fd_sc_hd__a22o_1
XU$$1419 t$5130 net1485 VGND VGND VPWR VPWR booth_b20_m21 sky130_fd_sc_hd__xor2_1
XFILLER_163_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_19__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_5_19__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_90_2 c$1804 s$1807 s$1809 VGND VGND VPWR VPWR c$2562 s$2563 sky130_fd_sc_hd__fa_1
XFILLER_100_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_83_1 c$1714 c$1716 c$1718 VGND VGND VPWR VPWR c$2504 s$2505 sky130_fd_sc_hd__fa_1
XFILLER_124_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_1135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_904 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_60_0 c$3632 c$3634 s$3637 VGND VGND VPWR VPWR c$4016 s$4017 sky130_fd_sc_hd__fa_1
XFILLER_183_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_76_0 s$833 c$1626 c$1628 VGND VGND VPWR VPWR c$2446 s$2447 sky130_fd_sc_hd__fa_1
XFILLER_124_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1520 net1521 VGND VGND VPWR VPWR net1520 sky130_fd_sc_hd__buf_2
Xfanout1531 net124 VGND VGND VPWR VPWR net1531 sky130_fd_sc_hd__buf_4
Xfanout1542 net123 VGND VGND VPWR VPWR net1542 sky130_fd_sc_hd__buf_4
XFILLER_39_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4001 net66 net458 net1218 net731 VGND VGND VPWR VPWR t$6450 sky130_fd_sc_hd__a22o_1
Xfanout1553 net1559 VGND VGND VPWR VPWR net1553 sky130_fd_sc_hd__buf_4
XFILLER_38_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4012 t$6455 net1282 VGND VGND VPWR VPWR booth_b58_m16 sky130_fd_sc_hd__xor2_1
Xfanout1564 net1565 VGND VGND VPWR VPWR net1564 sky130_fd_sc_hd__buf_4
XU$$4023 net1112 net453 net1103 net726 VGND VGND VPWR VPWR t$6461 sky130_fd_sc_hd__a22o_1
Xfanout1575 net1576 VGND VGND VPWR VPWR net1575 sky130_fd_sc_hd__buf_6
X_1120_ clknet_leaf_48_clk booth_b12_m3 VGND VGND VPWR VPWR pp_row15_6 sky130_fd_sc_hd__dfxtp_1
Xfanout1586 net1594 VGND VGND VPWR VPWR net1586 sky130_fd_sc_hd__buf_4
XU$$4034 t$6466 net1286 VGND VGND VPWR VPWR booth_b58_m27 sky130_fd_sc_hd__xor2_1
XFILLER_65_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4045 net1004 net455 net996 net728 VGND VGND VPWR VPWR t$6472 sky130_fd_sc_hd__a22o_1
XU$$3300 net1034 net496 net935 net769 VGND VGND VPWR VPWR t$6092 sky130_fd_sc_hd__a22o_1
Xfanout1597 net1598 VGND VGND VPWR VPWR net1597 sky130_fd_sc_hd__buf_4
XU$$3311 t$6097 net1346 VGND VGND VPWR VPWR booth_b48_m8 sky130_fd_sc_hd__xor2_1
XU$$4056 t$6477 net1290 VGND VGND VPWR VPWR booth_b58_m38 sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_112_1 c$2726 c$2728 c$2730 VGND VGND VPWR VPWR c$3364 s$3365 sky130_fd_sc_hd__fa_1
XU$$4067 net1736 net457 net1728 net730 VGND VGND VPWR VPWR t$6483 sky130_fd_sc_hd__a22o_1
XFILLER_20_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3322 net1196 net496 net1178 net769 VGND VGND VPWR VPWR t$6103 sky130_fd_sc_hd__a22o_1
XU$$3333 t$6108 net1343 VGND VGND VPWR VPWR booth_b48_m19 sky130_fd_sc_hd__xor2_1
X_1051_ clknet_leaf_248_clk net234 VGND VGND VPWR VPWR pp_row7_4 sky130_fd_sc_hd__dfxtp_2
XU$$4078 t$6488 net1285 VGND VGND VPWR VPWR booth_b58_m49 sky130_fd_sc_hd__xor2_1
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3344 net1082 net493 net1073 net766 VGND VGND VPWR VPWR t$6114 sky130_fd_sc_hd__a22o_1
XU$$4089 net1625 net456 net1616 net729 VGND VGND VPWR VPWR t$6494 sky130_fd_sc_hd__a22o_1
XU$$2610 t$5739 net1394 VGND VGND VPWR VPWR booth_b38_m0 sky130_fd_sc_hd__xor2_1
XU$$3355 t$6119 net1341 VGND VGND VPWR VPWR booth_b48_m30 sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_105_0 s$1965 c$2670 c$2672 VGND VGND VPWR VPWR c$3320 s$3321 sky130_fd_sc_hd__fa_1
XU$$2621 net1562 net543 net1520 net816 VGND VGND VPWR VPWR t$5745 sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_38_5 c$214 s$217 s$219 VGND VGND VPWR VPWR c$1192 s$1193 sky130_fd_sc_hd__fa_2
XU$$3366 net975 net494 net966 net767 VGND VGND VPWR VPWR t$6125 sky130_fd_sc_hd__a22o_1
XU$$2632 t$5750 net1395 VGND VGND VPWR VPWR booth_b38_m11 sky130_fd_sc_hd__xor2_1
XU$$3377 t$6130 net1340 VGND VGND VPWR VPWR booth_b48_m41 sky130_fd_sc_hd__xor2_1
XU$$2643 net1162 net549 net1150 net822 VGND VGND VPWR VPWR t$5756 sky130_fd_sc_hd__a22o_1
XU$$3388 net1706 net497 net1698 net770 VGND VGND VPWR VPWR t$6136 sky130_fd_sc_hd__a22o_1
XU$$3399 t$6141 net1344 VGND VGND VPWR VPWR booth_b48_m52 sky130_fd_sc_hd__xor2_1
XU$$2654 t$5761 net1395 VGND VGND VPWR VPWR booth_b38_m22 sky130_fd_sc_hd__xor2_1
XU$$2665 net1058 net549 net1054 net822 VGND VGND VPWR VPWR t$5767 sky130_fd_sc_hd__a22o_1
XU$$1920 net1453 VGND VGND VPWR VPWR notblock$5385\[2\] sky130_fd_sc_hd__inv_1
XU$$1931 t$5392 net1448 VGND VGND VPWR VPWR booth_b28_m3 sky130_fd_sc_hd__xor2_1
XU$$2676 t$5772 net1397 VGND VGND VPWR VPWR booth_b38_m33 sky130_fd_sc_hd__xor2_1
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1942 net1508 net587 net1499 net860 VGND VGND VPWR VPWR t$5398 sky130_fd_sc_hd__a22o_1
XU$$2687 net951 net545 net943 net818 VGND VGND VPWR VPWR t$5778 sky130_fd_sc_hd__a22o_1
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2698 t$5783 net1396 VGND VGND VPWR VPWR booth_b38_m44 sky130_fd_sc_hd__xor2_1
XU$$1953 t$5403 net1448 VGND VGND VPWR VPWR booth_b28_m14 sky130_fd_sc_hd__xor2_1
XFILLER_61_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1964 net1132 net584 net1116 net857 VGND VGND VPWR VPWR t$5409 sky130_fd_sc_hd__a22o_1
XU$$1975 t$5414 net1451 VGND VGND VPWR VPWR booth_b28_m25 sky130_fd_sc_hd__xor2_1
XU$$1986 net1026 net588 net1018 net861 VGND VGND VPWR VPWR t$5420 sky130_fd_sc_hd__a22o_1
XFILLER_159_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1997 t$5425 net1452 VGND VGND VPWR VPWR booth_b28_m36 sky130_fd_sc_hd__xor2_1
X_1953_ clknet_leaf_66_clk booth_b10_m44 VGND VGND VPWR VPWR pp_row54_5 sky130_fd_sc_hd__dfxtp_1
X_0904_ clknet_leaf_103_clk booth_b36_m60 VGND VGND VPWR VPWR pp_row96_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_119_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1884_ clknet_leaf_78_clk booth_b0_m52 VGND VGND VPWR VPWR pp_row52_0 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_98_1 s$3279 s$3281 s$3283 VGND VGND VPWR VPWR c$3790 s$3791 sky130_fd_sc_hd__fa_1
X_0835_ clknet_leaf_107_clk booth_b62_m30 VGND VGND VPWR VPWR pp_row92_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0766_ clknet_leaf_128_clk booth_b64_m54 VGND VGND VPWR VPWR pp_row118_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_170_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0697_ clknet_leaf_187_clk booth_b28_m59 VGND VGND VPWR VPWR pp_row87_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_9_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2436_ clknet_leaf_184_clk net142 VGND VGND VPWR VPWR pp_row111_10 sky130_fd_sc_hd__dfxtp_2
XFILLER_29_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2367_ clknet_leaf_98_clk booth_b62_m3 VGND VGND VPWR VPWR pp_row65_31 sky130_fd_sc_hd__dfxtp_1
XFILLER_99_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$605 final_adder.p_new$608 final_adder.g_new$617 final_adder.g_new$609
+ VGND VGND VPWR VPWR final_adder.g_new$733 sky130_fd_sc_hd__a21o_2
Xfinal_adder.U$$616 final_adder.p_new$628 final_adder.p_new$620 VGND VGND VPWR VPWR
+ final_adder.p_new$744 sky130_fd_sc_hd__and2_1
XFILLER_97_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1318_ clknet_leaf_247_clk booth_b4_m25 VGND VGND VPWR VPWR pp_row29_2 sky130_fd_sc_hd__dfxtp_1
XTAP_3909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$638 final_adder.p_new$662 final_adder.p_new$646 VGND VGND VPWR VPWR
+ final_adder.p_new$766 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$649 final_adder.p_new$656 final_adder.g_new$673 final_adder.g_new$657
+ VGND VGND VPWR VPWR final_adder.g_new$777 sky130_fd_sc_hd__a21o_1
X_2298_ clknet_leaf_199_clk booth_b2_m62 VGND VGND VPWR VPWR pp_row64_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_186_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1249_ clknet_leaf_111_clk booth_b52_m51 VGND VGND VPWR VPWR pp_row103_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_56_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$60 net1063 net442 net1055 net684 VGND VGND VPWR VPWR t$4437 sky130_fd_sc_hd__a22o_1
XU$$71 t$4442 net1569 VGND VGND VPWR VPWR booth_b0_m32 sky130_fd_sc_hd__xor2_1
XU$$82 net960 net443 net952 net685 VGND VGND VPWR VPWR t$4448 sky130_fd_sc_hd__a22o_1
XU$$93 t$4453 net1570 VGND VGND VPWR VPWR booth_b0_m43 sky130_fd_sc_hd__xor2_1
XFILLER_72_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_40 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_51 net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_62 net412 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_73 net441 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_84 net510 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_93_0 s$1853 c$2574 c$2576 VGND VGND VPWR VPWR c$3248 s$3249 sky130_fd_sc_hd__fa_1
XFILLER_153_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_95 net534 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_107_2 pp_row107_9 pp_row107_10 pp_row107_11 VGND VGND VPWR VPWR c$2698
+ s$2699 sky130_fd_sc_hd__fa_1
XFILLER_97_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1205 t$5020 net1014 VGND VGND VPWR VPWR booth_b16_m51 sky130_fd_sc_hd__xor2_1
XU$$1216 net1604 net648 net1595 net921 VGND VGND VPWR VPWR t$5026 sky130_fd_sc_hd__a22o_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1227 t$5031 net1012 VGND VGND VPWR VPWR booth_b16_m62 sky130_fd_sc_hd__xor2_1
XU$$1238 net10 net1013 VGND VGND VPWR VPWR sel_1$5038 sky130_fd_sc_hd__xor2_4
XU$$1249 net1672 net637 net1561 net910 VGND VGND VPWR VPWR t$5044 sky130_fd_sc_hd__a22o_1
XFILLER_70_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1010 final_adder.$signal$101 final_adder.g_new$1065 VGND VGND VPWR
+ VPWR net328 sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$1021 final_adder.$signal$1150 final_adder.g_new$935 VGND VGND VPWR
+ VPWR net341 sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$1032 final_adder.$signal$1161 final_adder.g_new$1054 VGND VGND VPWR
+ VPWR net353 sky130_fd_sc_hd__xor2_2
XFILLER_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1043 final_adder.$signal$1172 final_adder.g_new$1009 VGND VGND VPWR
+ VPWR net365 sky130_fd_sc_hd__xor2_2
XFILLER_7_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$1054 final_adder.$signal$1183 final_adder.g_new$1043 VGND VGND VPWR
+ VPWR net377 sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$1065 final_adder.$signal$1194 final_adder.g_new$987 VGND VGND VPWR
+ VPWR net262 sky130_fd_sc_hd__xor2_1
X_0620_ clknet_leaf_187_clk booth_b28_m56 VGND VGND VPWR VPWR pp_row84_5 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$1076 final_adder.$signal$1205 final_adder.g_new$1032 VGND VGND VPWR
+ VPWR net274 sky130_fd_sc_hd__xor2_2
XFILLER_137_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$1087 final_adder.$signal$1216 final_adder.g_new$965 VGND VGND VPWR
+ VPWR net286 sky130_fd_sc_hd__xor2_2
X_0551_ clknet_leaf_171_clk booth_b52_m29 VGND VGND VPWR VPWR pp_row81_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_139_1041 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0482_ clknet_leaf_157_clk booth_b32_m47 VGND VGND VPWR VPWR pp_row79_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_140_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2221_ clknet_leaf_231_clk net214 VGND VGND VPWR VPWR pp_row61_31 sky130_fd_sc_hd__dfxtp_1
XFILLER_61_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1350 net1352 VGND VGND VPWR VPWR net1350 sky130_fd_sc_hd__buf_6
Xfanout1361 net1366 VGND VGND VPWR VPWR net1361 sky130_fd_sc_hd__clkbuf_4
X_2152_ clknet_leaf_215_clk booth_b4_m56 VGND VGND VPWR VPWR pp_row60_2 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_50_4 s$353 s$355 s$357 VGND VGND VPWR VPWR c$1334 s$1335 sky130_fd_sc_hd__fa_1
Xfanout1372 net1375 VGND VGND VPWR VPWR net1372 sky130_fd_sc_hd__buf_6
XFILLER_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1383 net1384 VGND VGND VPWR VPWR net1383 sky130_fd_sc_hd__buf_4
XFILLER_66_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1394 net33 VGND VGND VPWR VPWR net1394 sky130_fd_sc_hd__buf_6
X_1103_ clknet_leaf_14_clk booth_b2_m12 VGND VGND VPWR VPWR pp_row14_1 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_43_3 c$244 c$246 c$248 VGND VGND VPWR VPWR c$1248 s$1249 sky130_fd_sc_hd__fa_1
XU$$3130 net1626 net516 net1618 net789 VGND VGND VPWR VPWR t$6004 sky130_fd_sc_hd__a22o_1
XFILLER_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2083_ clknet_leaf_143_clk booth_b46_m63 VGND VGND VPWR VPWR pp_row109_1 sky130_fd_sc_hd__dfxtp_1
XU$$3141 t$6009 net1364 VGND VGND VPWR VPWR booth_b44_m60 sky130_fd_sc_hd__xor2_1
XFILLER_4_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2335_1775 VGND VGND VPWR VPWR U$$2335_1775/HI net1775 sky130_fd_sc_hd__conb_1
XU$$3152 net41 VGND VGND VPWR VPWR notblock$6015\[1\] sky130_fd_sc_hd__inv_1
X_1034_ clknet_leaf_248_clk net201 VGND VGND VPWR VPWR pp_row4_4 sky130_fd_sc_hd__dfxtp_4
XU$$3163 net1034 net501 net935 net774 VGND VGND VPWR VPWR t$6022 sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_36_2 pp_row36_11 pp_row36_12 pp_row36_13 VGND VGND VPWR VPWR c$1162 s$1163
+ sky130_fd_sc_hd__fa_1
XU$$3174 t$6027 net1353 VGND VGND VPWR VPWR booth_b46_m8 sky130_fd_sc_hd__xor2_1
XU$$3185 net1193 net501 net1177 net774 VGND VGND VPWR VPWR t$6033 sky130_fd_sc_hd__a22o_1
XU$$2440 t$5651 net1426 VGND VGND VPWR VPWR booth_b34_m52 sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_13_1 s$2769 s$2771 s$2773 VGND VGND VPWR VPWR c$3450 s$3451 sky130_fd_sc_hd__fa_1
XU$$2451 net1602 net567 net1592 net840 VGND VGND VPWR VPWR t$5657 sky130_fd_sc_hd__a22o_1
XU$$3196 t$6038 net1353 VGND VGND VPWR VPWR booth_b46_m19 sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_29_1 pp_row29_3 pp_row29_4 pp_row29_5 VGND VGND VPWR VPWR c$1084 s$1085
+ sky130_fd_sc_hd__fa_1
XU$$2462 t$5662 net1428 VGND VGND VPWR VPWR booth_b34_m63 sky130_fd_sc_hd__xor2_1
XFILLER_62_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2473 t$5669 net1406 VGND VGND VPWR VPWR booth_b36_m0 sky130_fd_sc_hd__xor2_1
XU$$2484 net1560 net551 net1520 net824 VGND VGND VPWR VPWR t$5675 sky130_fd_sc_hd__a22o_1
XU$$2495 t$5680 net1403 VGND VGND VPWR VPWR booth_b36_m11 sky130_fd_sc_hd__xor2_1
XU$$1750 net1679 net607 net1654 net880 VGND VGND VPWR VPWR t$5299 sky130_fd_sc_hd__a22o_1
XU$$1761 t$5304 net1471 VGND VGND VPWR VPWR booth_b24_m55 sky130_fd_sc_hd__xor2_1
XFILLER_61_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_957 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1772 net1553 net607 net1544 net880 VGND VGND VPWR VPWR t$5310 sky130_fd_sc_hd__a22o_1
XFILLER_148_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1783 net1463 VGND VGND VPWR VPWR notblock$5315\[2\] sky130_fd_sc_hd__inv_1
XFILLER_188_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1794 t$5322 net1457 VGND VGND VPWR VPWR booth_b26_m3 sky130_fd_sc_hd__xor2_1
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1936_ clknet_leaf_70_clk booth_b38_m15 VGND VGND VPWR VPWR pp_row53_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_174_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1867_ clknet_leaf_66_clk booth_b24_m27 VGND VGND VPWR VPWR pp_row51_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_147_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput60 a[63] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_1
XFILLER_190_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0818_ clknet_leaf_109_clk booth_b34_m58 VGND VGND VPWR VPWR pp_row92_4 sky130_fd_sc_hd__dfxtp_1
Xinput71 b[15] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_6
X_1798_ clknet_leaf_219_clk booth_b8_m41 VGND VGND VPWR VPWR pp_row49_4 sky130_fd_sc_hd__dfxtp_1
Xinput82 b[25] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput93 b[35] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0749_ clknet_leaf_160_clk booth_b32_m57 VGND VGND VPWR VPWR pp_row89_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_143_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2419_ clknet_leaf_145_clk booth_b20_m47 VGND VGND VPWR VPWR pp_row67_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_29_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$402 final_adder.p_new$408 final_adder.p_new$404 VGND VGND VPWR VPWR
+ final_adder.p_new$530 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$413 final_adder.p_new$414 final_adder.g_new$419 final_adder.g_new$415
+ VGND VGND VPWR VPWR final_adder.g_new$541 sky130_fd_sc_hd__a21o_1
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$424 final_adder.p_new$430 final_adder.p_new$426 VGND VGND VPWR VPWR
+ final_adder.p_new$552 sky130_fd_sc_hd__and2_1
XTAP_3706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$435 final_adder.p_new$436 final_adder.g_new$441 final_adder.g_new$437
+ VGND VGND VPWR VPWR final_adder.g_new$563 sky130_fd_sc_hd__a21o_1
XTAP_3717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$446 final_adder.p_new$452 final_adder.p_new$448 VGND VGND VPWR VPWR
+ final_adder.p_new$574 sky130_fd_sc_hd__and2_1
XTAP_3728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$457 final_adder.p_new$458 final_adder.g_new$463 final_adder.g_new$459
+ VGND VGND VPWR VPWR final_adder.g_new$585 sky130_fd_sc_hd__a21o_1
XTAP_3739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$307 t$4562 net1274 VGND VGND VPWR VPWR booth_b4_m13 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$468 final_adder.p_new$474 final_adder.p_new$470 VGND VGND VPWR VPWR
+ final_adder.p_new$596 sky130_fd_sc_hd__and2_1
XFILLER_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$318 net1143 net532 net1133 net805 VGND VGND VPWR VPWR t$4568 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$479 final_adder.p_new$480 final_adder.g_new$485 final_adder.g_new$481
+ VGND VGND VPWR VPWR final_adder.g_new$607 sky130_fd_sc_hd__a21o_1
XU$$329 t$4573 net1273 VGND VGND VPWR VPWR booth_b4_m24 sky130_fd_sc_hd__xor2_1
XFILLER_38_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_112_0 net1910 pp_row112_1 pp_row112_2 VGND VGND VPWR VPWR c$2732 s$2733
+ sky130_fd_sc_hd__fa_1
XFILLER_180_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2874_1784 VGND VGND VPWR VPWR U$$2874_1784/HI net1784 sky130_fd_sc_hd__conb_1
XFILLER_180_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_60_3 s$1451 s$1453 s$1455 VGND VGND VPWR VPWR c$2324 s$2325 sky130_fd_sc_hd__fa_1
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_53_2 c$1360 s$1363 s$1365 VGND VGND VPWR VPWR c$2266 s$2267 sky130_fd_sc_hd__fa_1
XFILLER_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_0_69_2 pp_row69_6 pp_row69_7 pp_row69_8 VGND VGND VPWR VPWR c$148 s$149
+ sky130_fd_sc_hd__fa_1
XFILLER_180_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_46_1 c$1270 c$1272 c$1274 VGND VGND VPWR VPWR c$2208 s$2209 sky130_fd_sc_hd__fa_1
XFILLER_169_1023 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_23_0 c$3484 c$3486 s$3489 VGND VGND VPWR VPWR c$3942 s$3943 sky130_fd_sc_hd__fa_1
Xdadda_fa_3_39_0 s$227 c$1182 c$1184 VGND VGND VPWR VPWR c$2150 s$2151 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$980 final_adder.$signal$1109 final_adder.g_new$1080 VGND VGND VPWR
+ VPWR net295 sky130_fd_sc_hd__xor2_2
XFILLER_75_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$830 net1231 net397 net1127 net663 VGND VGND VPWR VPWR t$4830 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$991 final_adder.$signal$1120 final_adder.g_new$853 VGND VGND VPWR
+ VPWR net308 sky130_fd_sc_hd__xor2_2
XU$$841 t$4835 net1312 VGND VGND VPWR VPWR booth_b12_m6 sky130_fd_sc_hd__xor2_1
XU$$852 net1211 net394 net1203 net660 VGND VGND VPWR VPWR t$4841 sky130_fd_sc_hd__a22o_1
XU$$863 t$4846 net1310 VGND VGND VPWR VPWR booth_b12_m17 sky130_fd_sc_hd__xor2_1
XU$$1002 t$4917 net1186 VGND VGND VPWR VPWR booth_b14_m18 sky130_fd_sc_hd__xor2_1
XU$$1013 net1091 net387 net1083 net653 VGND VGND VPWR VPWR t$4923 sky130_fd_sc_hd__a22o_1
XU$$874 net1101 net397 net1092 net663 VGND VGND VPWR VPWR t$4852 sky130_fd_sc_hd__a22o_1
XU$$1024 t$4928 net1184 VGND VGND VPWR VPWR booth_b14_m29 sky130_fd_sc_hd__xor2_1
XU$$885 t$4857 net1311 VGND VGND VPWR VPWR booth_b12_m28 sky130_fd_sc_hd__xor2_1
XU$$1035 net983 net390 net974 net656 VGND VGND VPWR VPWR t$4934 sky130_fd_sc_hd__a22o_1
XU$$896 net990 net393 net982 net659 VGND VGND VPWR VPWR t$4863 sky130_fd_sc_hd__a22o_1
XFILLER_43_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1046 t$4939 net1186 VGND VGND VPWR VPWR booth_b14_m40 sky130_fd_sc_hd__xor2_1
XU$$1057 net1711 net390 net1703 net656 VGND VGND VPWR VPWR t$4945 sky130_fd_sc_hd__a22o_1
XU$$1068 t$4950 net1191 VGND VGND VPWR VPWR booth_b14_m51 sky130_fd_sc_hd__xor2_1
XU$$1079 net1604 net390 net1595 net656 VGND VGND VPWR VPWR t$4956 sky130_fd_sc_hd__a22o_1
XFILLER_188_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1721_ clknet_leaf_22_clk booth_b26_m20 VGND VGND VPWR VPWR pp_row46_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_117_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1652_ clknet_leaf_235_clk net194 VGND VGND VPWR VPWR pp_row43_22 sky130_fd_sc_hd__dfxtp_1
XFILLER_172_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_98_4 pp_row98_12 pp_row98_13 pp_row98_14 VGND VGND VPWR VPWR c$1910 s$1911
+ sky130_fd_sc_hd__fa_1
XFILLER_176_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0603_ clknet_leaf_174_clk booth_b46_m37 VGND VGND VPWR VPWR pp_row83_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_99_913 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1583_ clknet_leaf_109_clk booth_b56_m49 VGND VGND VPWR VPWR pp_row105_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_113_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0534_ clknet_leaf_159_clk booth_b20_m61 VGND VGND VPWR VPWR pp_row81_2 sky130_fd_sc_hd__dfxtp_1
Xfanout609 sel_0$5247 VGND VGND VPWR VPWR net609 sky130_fd_sc_hd__buf_6
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4413_1827 VGND VGND VPWR VPWR U$$4413_1827/HI net1827 sky130_fd_sc_hd__conb_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0465_ clknet_leaf_205_clk booth_b56_m22 VGND VGND VPWR VPWR pp_row78_22 sky130_fd_sc_hd__dfxtp_1
XFILLER_98_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2204_ clknet_leaf_88_clk booth_b32_m29 VGND VGND VPWR VPWR pp_row61_16 sky130_fd_sc_hd__dfxtp_1
X_0396_ clknet_leaf_191_clk booth_b40_m36 VGND VGND VPWR VPWR pp_row76_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1180 net1181 VGND VGND VPWR VPWR net1180 sky130_fd_sc_hd__clkbuf_4
XFILLER_152_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1191 net7 VGND VGND VPWR VPWR net1191 sky130_fd_sc_hd__buf_6
XFILLER_39_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2135_ clknet_leaf_27_clk booth_b36_m23 VGND VGND VPWR VPWR pp_row59_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_27_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_41_0 pp_row41_11 pp_row41_12 pp_row41_13 VGND VGND VPWR VPWR c$1218 s$1219
+ sky130_fd_sc_hd__fa_1
XFILLER_187_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2066_ clknet_leaf_43_clk booth_b34_m23 VGND VGND VPWR VPWR pp_row57_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_35_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1017_ clknet_leaf_60_clk booth_b0_m0 VGND VGND VPWR VPWR pp_row0_0 sky130_fd_sc_hd__dfxtp_1
XU$$2270 net979 net575 net970 net848 VGND VGND VPWR VPWR t$5565 sky130_fd_sc_hd__a22o_1
XU$$2281 t$5570 net1431 VGND VGND VPWR VPWR booth_b32_m41 sky130_fd_sc_hd__xor2_1
XU$$2292 net1704 net573 net1696 net846 VGND VGND VPWR VPWR t$5576 sky130_fd_sc_hd__a22o_1
XFILLER_22_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1580 t$5212 net1479 VGND VGND VPWR VPWR booth_b22_m33 sky130_fd_sc_hd__xor2_1
XU$$1591 net948 net612 net941 net885 VGND VGND VPWR VPWR t$5218 sky130_fd_sc_hd__a22o_1
XFILLER_120_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1919_ clknet_leaf_80_clk booth_b6_m47 VGND VGND VPWR VPWR pp_row53_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_191_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_70_2 s$2401 s$2403 s$2405 VGND VGND VPWR VPWR c$3114 s$3115 sky130_fd_sc_hd__fa_1
Xdadda_fa_1_86_2 pp_row86_6 pp_row86_7 pp_row86_8 VGND VGND VPWR VPWR c$982 s$983
+ sky130_fd_sc_hd__fa_1
Xdadda_fa_4_63_1 c$2338 c$2340 s$2343 VGND VGND VPWR VPWR c$3070 s$3071 sky130_fd_sc_hd__fa_1
Xdadda_fa_1_79_1 pp_row79_3 pp_row79_4 pp_row79_5 VGND VGND VPWR VPWR c$872 s$873
+ sky130_fd_sc_hd__fa_1
XFILLER_76_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_40_0 s$3559 c$3974 s$3977 VGND VGND VPWR VPWR c$4232 s$4233 sky130_fd_sc_hd__fa_1
Xdadda_fa_4_56_0 s$1409 c$2278 c$2280 VGND VGND VPWR VPWR c$3026 s$3027 sky130_fd_sc_hd__fa_1
XTAP_4204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$210 final_adder.$signal$1134 final_adder.$signal$1135 VGND VGND VPWR
+ VPWR final_adder.p_new$338 sky130_fd_sc_hd__and2_1
XTAP_4226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$221 final_adder.$signal$1125 final_adder.$signal$70 final_adder.$signal$72
+ VGND VGND VPWR VPWR final_adder.g_new$349 sky130_fd_sc_hd__a21o_1
XTAP_4248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$232 final_adder.$signal$1112 final_adder.$signal$1113 VGND VGND VPWR
+ VPWR final_adder.p_new$360 sky130_fd_sc_hd__and2_1
XTAP_4259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$243 final_adder.$signal$1103 final_adder.$signal$26 final_adder.$signal$28
+ VGND VGND VPWR VPWR final_adder.g_new$371 sky130_fd_sc_hd__a21o_1
XTAP_3525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$104 net1690 net449 net1682 net691 VGND VGND VPWR VPWR t$4459 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$265 final_adder.p_new$264 final_adder.g_new$267 final_adder.g_new$265
+ VGND VGND VPWR VPWR final_adder.g_new$393 sky130_fd_sc_hd__a21o_1
XFILLER_100_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$115 t$4464 net1576 VGND VGND VPWR VPWR booth_b0_m54 sky130_fd_sc_hd__xor2_1
XTAP_3547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$276 final_adder.p_new$278 final_adder.p_new$276 VGND VGND VPWR VPWR
+ final_adder.p_new$404 sky130_fd_sc_hd__and2_1
XTAP_3558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$287 final_adder.p_new$286 final_adder.g_new$289 final_adder.g_new$287
+ VGND VGND VPWR VPWR final_adder.g_new$415 sky130_fd_sc_hd__a21o_1
XU$$126 net1581 net445 net1552 net687 VGND VGND VPWR VPWR t$4470 sky130_fd_sc_hd__a22o_1
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$137 net1571 VGND VGND VPWR VPWR notblock$4475\[0\] sky130_fd_sc_hd__inv_1
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$298 final_adder.p_new$300 final_adder.p_new$298 VGND VGND VPWR VPWR
+ final_adder.p_new$426 sky130_fd_sc_hd__and2_1
XU$$148 t$4481 net1390 VGND VGND VPWR VPWR booth_b2_m2 sky130_fd_sc_hd__xor2_1
XFILLER_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_879 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$159 net1515 net623 net1508 net896 VGND VGND VPWR VPWR t$4487 sky130_fd_sc_hd__a22o_1
XFILLER_168_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_120_0_1913 VGND VGND VPWR VPWR net1913 dadda_fa_4_120_0_1913/LO sky130_fd_sc_hd__conb_1
XFILLER_127_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_74_0 net1894 pp_row74_1 pp_row74_2 VGND VGND VPWR VPWR c$186 s$187 sky130_fd_sc_hd__fa_1
XFILLER_0_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0250_ clknet_leaf_209_clk booth_b10_m62 VGND VGND VPWR VPWR pp_row72_2 sky130_fd_sc_hd__dfxtp_1
Xinput250 c[94] VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0181_ clknet_leaf_147_clk booth_b6_m64 VGND VGND VPWR VPWR pp_row70_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_64_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$660 net1638 net411 net1629 net677 VGND VGND VPWR VPWR t$4742 sky130_fd_sc_hd__a22o_1
XFILLER_90_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$671 t$4747 net1242 VGND VGND VPWR VPWR booth_b8_m58 sky130_fd_sc_hd__xor2_1
XFILLER_44_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$682 net1527 net412 net1884 net678 VGND VGND VPWR VPWR t$4753 sky130_fd_sc_hd__a22o_1
XU$$693 net1230 net404 net1126 net670 VGND VGND VPWR VPWR t$4760 sky130_fd_sc_hd__a22o_1
XFILLER_189_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_990 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1704_ clknet_leaf_23_clk booth_b44_m1 VGND VGND VPWR VPWR pp_row45_22 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_80_1 s$3171 s$3173 s$3175 VGND VGND VPWR VPWR c$3718 s$3719 sky130_fd_sc_hd__fa_1
XFILLER_144_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_96_1 pp_row96_5 pp_row96_6 pp_row96_7 VGND VGND VPWR VPWR c$1880 s$1881
+ sky130_fd_sc_hd__fa_1
XFILLER_172_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1635_ clknet_leaf_239_clk booth_b14_m29 VGND VGND VPWR VPWR pp_row43_7 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_73_0 c$3122 c$3124 c$3126 VGND VGND VPWR VPWR c$3688 s$3689 sky130_fd_sc_hd__fa_1
Xdadda_fa_2_89_0 pp_row89_12 pp_row89_13 pp_row89_14 VGND VGND VPWR VPWR c$1794 s$1795
+ sky130_fd_sc_hd__fa_1
XFILLER_63_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1566_ clknet_leaf_7_clk booth_b28_m12 VGND VGND VPWR VPWR pp_row40_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_113_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout406 net407 VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__buf_4
Xfanout417 sel_0$4687 VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__buf_6
XFILLER_98_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout428 net433 VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_72_8 s$173 s$175 s$177 VGND VGND VPWR VPWR c$760 s$761 sky130_fd_sc_hd__fa_2
XFILLER_59_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0517_ clknet_leaf_155_clk booth_b42_m38 VGND VGND VPWR VPWR pp_row80_14 sky130_fd_sc_hd__dfxtp_1
Xfanout439 net440 VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__buf_4
XFILLER_87_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1497_ clknet_leaf_45_clk booth_b30_m7 VGND VGND VPWR VPWR pp_row37_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_141_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_65_7 c$94 s$97 s$99 VGND VGND VPWR VPWR c$632 s$633 sky130_fd_sc_hd__fa_1
X_0448_ clknet_leaf_206_clk booth_b24_m54 VGND VGND VPWR VPWR pp_row78_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_104_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_58_6 pp_row58_29 pp_row58_30 pp_row58_31 VGND VGND VPWR VPWR c$504 s$505
+ sky130_fd_sc_hd__fa_1
XFILLER_67_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0379_ clknet_leaf_197_clk net229 VGND VGND VPWR VPWR pp_row75_28 sky130_fd_sc_hd__dfxtp_1
XFILLER_27_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2118_ clknet_leaf_218_clk booth_b4_m55 VGND VGND VPWR VPWR pp_row59_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_55_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2049_ clknet_leaf_136_clk booth_b64_m44 VGND VGND VPWR VPWR pp_row108_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_35_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_170_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_170_clk
+ sky130_fd_sc_hd__clkbuf_16
Xdadda_ha_1_92_2 pp_row92_6 pp_row92_7 VGND VGND VPWR VPWR c$1036 s$1037 sky130_fd_sc_hd__ha_1
XFILLER_7_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_88_0 s$3751 c$4070 s$4073 VGND VGND VPWR VPWR c$4328 s$4329 sky130_fd_sc_hd__fa_2
XFILLER_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_91_0 pp_row91_0 pp_row91_1 pp_row91_2 VGND VGND VPWR VPWR c$1026 s$1027
+ sky130_fd_sc_hd__fa_1
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout940 net941 VGND VGND VPWR VPWR net940 sky130_fd_sc_hd__buf_4
Xfanout951 net952 VGND VGND VPWR VPWR net951 sky130_fd_sc_hd__buf_4
Xfanout962 net963 VGND VGND VPWR VPWR net962 sky130_fd_sc_hd__buf_6
XTAP_4001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4408 net1507 sel_0$6647 net1502 net694 VGND VGND VPWR VPWR t$6658 sky130_fd_sc_hd__a22o_1
XTAP_4012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout973 net974 VGND VGND VPWR VPWR net973 sky130_fd_sc_hd__buf_4
XU$$4419 t$6663 net1830 VGND VGND VPWR VPWR booth_b64_m14 sky130_fd_sc_hd__xor2_1
XTAP_4023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout984 net986 VGND VGND VPWR VPWR net984 sky130_fd_sc_hd__buf_4
XTAP_4034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout995 net997 VGND VGND VPWR VPWR net995 sky130_fd_sc_hd__buf_4
XTAP_4045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_662 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3707 net1233 net475 net1129 net748 VGND VGND VPWR VPWR t$6300 sky130_fd_sc_hd__a22o_1
XFILLER_46_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3718 t$6305 net1300 VGND VGND VPWR VPWR booth_b54_m6 sky130_fd_sc_hd__xor2_1
XTAP_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3729 net1217 net472 net1208 net745 VGND VGND VPWR VPWR t$6311 sky130_fd_sc_hd__a22o_1
XTAP_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_103_0 c$3804 c$3806 s$3809 VGND VGND VPWR VPWR c$4102 s$4103 sky130_fd_sc_hd__fa_1
XFILLER_100_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_300 net392 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_311 net544 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_322 net622 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_333 net713 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_23_3 pp_row23_11 pp_row23_12 c$1050 VGND VGND VPWR VPWR c$2028 s$2029
+ sky130_fd_sc_hd__fa_1
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_344 net841 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_355 net939 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_366 net1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_377 net1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_388 net1507 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_399 net1627 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_161_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_161_clk
+ sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_3_114_0_1911 VGND VGND VPWR VPWR net1911 dadda_fa_3_114_0_1911/LO sky130_fd_sc_hd__conb_1
XFILLER_13_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_90_0 c$3752 c$3754 s$3757 VGND VGND VPWR VPWR c$4076 s$4077 sky130_fd_sc_hd__fa_2
XFILLER_103_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_997 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3568_1795 VGND VGND VPWR VPWR U$$3568_1795/HI net1795 sky130_fd_sc_hd__conb_1
XFILLER_108_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1420_ clknet_leaf_54_clk booth_b10_m24 VGND VGND VPWR VPWR pp_row34_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_170_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1351_ clknet_leaf_241_clk net1439 VGND VGND VPWR VPWR pp_row30_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_96_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_68_5 s$683 s$685 s$687 VGND VGND VPWR VPWR c$1552 s$1553 sky130_fd_sc_hd__fa_1
X_0302_ clknet_leaf_227_clk booth_b42_m31 VGND VGND VPWR VPWR pp_row73_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_96_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1282_ clknet_leaf_120_clk booth_b58_m45 VGND VGND VPWR VPWR pp_row103_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_110_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0233_ clknet_leaf_125_clk booth_b50_m63 VGND VGND VPWR VPWR pp_row113_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_110_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$490 t$4655 net1244 VGND VGND VPWR VPWR booth_b6_m36 sky130_fd_sc_hd__xor2_1
XFILLER_189_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_152_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_152_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_20_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0997_ clknet_leaf_119_clk notsign$5734 VGND VGND VPWR VPWR pp_row101_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_146_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1618_ clknet_leaf_241_clk booth_b30_m12 VGND VGND VPWR VPWR pp_row42_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_120_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1549_ clknet_leaf_236_clk net189 VGND VGND VPWR VPWR pp_row39_20 sky130_fd_sc_hd__dfxtp_2
XFILLER_86_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_70_5 pp_row70_29 pp_row70_30 pp_row70_31 VGND VGND VPWR VPWR c$718 s$719
+ sky130_fd_sc_hd__fa_1
XFILLER_59_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_63_4 pp_row63_29 pp_row63_30 pp_row63_31 VGND VGND VPWR VPWR c$590 s$591
+ sky130_fd_sc_hd__fa_1
XFILLER_28_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_56_3 pp_row56_17 pp_row56_18 pp_row56_19 VGND VGND VPWR VPWR c$462 s$463
+ sky130_fd_sc_hd__fa_1
XFILLER_41_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_846 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_33_2 s$2105 s$2107 s$2109 VGND VGND VPWR VPWR c$2892 s$2893 sky130_fd_sc_hd__fa_1
Xdadda_fa_1_49_2 pp_row49_6 pp_row49_7 pp_row49_8 VGND VGND VPWR VPWR c$336 s$337
+ sky130_fd_sc_hd__fa_1
XU$$4465_1853 VGND VGND VPWR VPWR U$$4465_1853/HI net1853 sky130_fd_sc_hd__conb_1
Xdadda_fa_4_26_1 c$2042 c$2044 s$2047 VGND VGND VPWR VPWR c$2848 s$2849 sky130_fd_sc_hd__fa_1
XFILLER_83_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_19_0 pp_row19_8 pp_row19_9 pp_row19_10 VGND VGND VPWR VPWR c$2804 s$2805
+ sky130_fd_sc_hd__fa_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_143_clk clknet_5_25__leaf_clk VGND VGND VPWR VPWR clknet_leaf_143_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_11_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1702 net106 VGND VGND VPWR VPWR net1702 sky130_fd_sc_hd__buf_6
XFILLER_105_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1713 net1714 VGND VGND VPWR VPWR net1713 sky130_fd_sc_hd__buf_4
XFILLER_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1724 net1728 VGND VGND VPWR VPWR net1724 sky130_fd_sc_hd__buf_4
Xfanout1735 net1736 VGND VGND VPWR VPWR net1735 sky130_fd_sc_hd__buf_6
XFILLER_78_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1746 net1752 VGND VGND VPWR VPWR net1746 sky130_fd_sc_hd__buf_6
XU$$4205 t$6553 net1271 VGND VGND VPWR VPWR booth_b60_m44 sky130_fd_sc_hd__xor2_1
XFILLER_120_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout770 net773 VGND VGND VPWR VPWR net770 sky130_fd_sc_hd__buf_4
XFILLER_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4216 net1685 net440 net1659 net722 VGND VGND VPWR VPWR t$6559 sky130_fd_sc_hd__a22o_1
Xfanout781 net782 VGND VGND VPWR VPWR net781 sky130_fd_sc_hd__buf_4
XU$$4227 t$6564 net1270 VGND VGND VPWR VPWR booth_b60_m55 sky130_fd_sc_hd__xor2_1
XFILLER_172_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout792 net793 VGND VGND VPWR VPWR net792 sky130_fd_sc_hd__buf_4
XU$$4238 net1554 net437 net1545 net719 VGND VGND VPWR VPWR t$6570 sky130_fd_sc_hd__a22o_1
XU$$3504 t$6195 net1331 VGND VGND VPWR VPWR booth_b50_m36 sky130_fd_sc_hd__xor2_1
XU$$2472_1777 VGND VGND VPWR VPWR U$$2472_1777/HI net1777 sky130_fd_sc_hd__conb_1
XFILLER_93_749 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4249 net1256 VGND VGND VPWR VPWR notblock$6575\[2\] sky130_fd_sc_hd__inv_1
XFILLER_86_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3515 net1750 net489 net1742 net762 VGND VGND VPWR VPWR t$6201 sky130_fd_sc_hd__a22o_1
XU$$3526 t$6206 net1335 VGND VGND VPWR VPWR booth_b50_m47 sky130_fd_sc_hd__xor2_1
XTAP_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3537 net1644 net490 net1635 net763 VGND VGND VPWR VPWR t$6212 sky130_fd_sc_hd__a22o_1
XFILLER_46_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2803 t$5837 net1382 VGND VGND VPWR VPWR booth_b40_m28 sky130_fd_sc_hd__xor2_1
XU$$3548 t$6217 net1334 VGND VGND VPWR VPWR booth_b50_m58 sky130_fd_sc_hd__xor2_1
XTAP_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2814 net91 net535 net983 net808 VGND VGND VPWR VPWR t$5843 sky130_fd_sc_hd__a22o_1
XFILLER_46_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3559 net1533 net489 net1794 net762 VGND VGND VPWR VPWR t$6223 sky130_fd_sc_hd__a22o_1
XTAP_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2825 t$5848 net1378 VGND VGND VPWR VPWR booth_b40_m39 sky130_fd_sc_hd__xor2_1
XFILLER_65_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2836 net1723 net538 net1714 net811 VGND VGND VPWR VPWR t$5854 sky130_fd_sc_hd__a22o_1
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_130 net703 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdadda_fa_3_21_0 pp_row21_0 pp_row21_1 pp_row21_2 VGND VGND VPWR VPWR c$2006 s$2007
+ sky130_fd_sc_hd__fa_1
XU$$2847 t$5859 net1383 VGND VGND VPWR VPWR booth_b40_m50 sky130_fd_sc_hd__xor2_1
XTAP_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2858 net1619 net540 net1611 net813 VGND VGND VPWR VPWR t$5865 sky130_fd_sc_hd__a22o_1
XANTENNA_141 net765 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2869 t$5870 net1383 VGND VGND VPWR VPWR booth_b40_m61 sky130_fd_sc_hd__xor2_1
XANTENNA_152 net799 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_163 net874 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_174 net917 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_185 net968 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_196 net1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0920_ clknet_leaf_185_clk net252 VGND VGND VPWR VPWR pp_row96_18 sky130_fd_sc_hd__dfxtp_4
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_134_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_134_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_187_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0851_ clknet_leaf_144_clk booth_b52_m41 VGND VGND VPWR VPWR pp_row93_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0782_ clknet_leaf_140_clk booth_b50_m40 VGND VGND VPWR VPWR pp_row90_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_80_4 s$893 s$895 s$897 VGND VGND VPWR VPWR c$1694 s$1695 sky130_fd_sc_hd__fa_1
X_2452_ clknet_leaf_92_clk booth_b16_m52 VGND VGND VPWR VPWR pp_row68_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_73_3 c$760 s$763 s$765 VGND VGND VPWR VPWR c$1608 s$1609 sky130_fd_sc_hd__fa_1
X_1403_ clknet_leaf_51_clk booth_b16_m17 VGND VGND VPWR VPWR pp_row33_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2383_ clknet_leaf_83_clk booth_b24_m42 VGND VGND VPWR VPWR pp_row66_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_25_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_66_2 c$628 c$630 c$632 VGND VGND VPWR VPWR c$1522 s$1523 sky130_fd_sc_hd__fa_1
X_1334_ clknet_leaf_0_clk booth_b2_m28 VGND VGND VPWR VPWR pp_row30_1 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$809 final_adder.p_new$824 final_adder.g_new$857 final_adder.g_new$825
+ VGND VGND VPWR VPWR final_adder.g_new$937 sky130_fd_sc_hd__a21o_1
Xdadda_fa_5_43_1 s$2949 s$2951 s$2953 VGND VGND VPWR VPWR c$3570 s$3571 sky130_fd_sc_hd__fa_1
XFILLER_111_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_59_1 c$496 c$498 c$500 VGND VGND VPWR VPWR c$1436 s$1437 sky130_fd_sc_hd__fa_1
X_1265_ clknet_leaf_2_clk booth_b6_m20 VGND VGND VPWR VPWR pp_row26_3 sky130_fd_sc_hd__dfxtp_1
Xinput3 a[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_6
Xdadda_fa_5_36_0 c$2900 c$2902 c$2904 VGND VGND VPWR VPWR c$3540 s$3541 sky130_fd_sc_hd__fa_1
XFILLER_36_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0216_ clknet_leaf_198_clk booth_b8_m63 VGND VGND VPWR VPWR pp_row71_1 sky130_fd_sc_hd__dfxtp_1
X_1196_ clknet_leaf_51_clk booth_b16_m5 VGND VGND VPWR VPWR pp_row21_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_65_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_125_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_125_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_20_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_110_0 c$3344 c$3346 c$3348 VGND VGND VPWR VPWR c$3836 s$3837 sky130_fd_sc_hd__fa_1
XFILLER_192_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4495_1868 VGND VGND VPWR VPWR U$$4495_1868/HI net1868 sky130_fd_sc_hd__conb_1
Xfinal_adder.U$$1 c$4152 s$4155 VGND VGND VPWR VPWR final_adder.$signal$4 final_adder.$signal$1091
+ sky130_fd_sc_hd__ha_1
XFILLER_146_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput340 net340 VGND VGND VPWR VPWR o[5] sky130_fd_sc_hd__buf_2
XFILLER_134_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput351 net351 VGND VGND VPWR VPWR o[6] sky130_fd_sc_hd__buf_2
Xoutput362 net362 VGND VGND VPWR VPWR o[7] sky130_fd_sc_hd__buf_2
XFILLER_160_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput373 net373 VGND VGND VPWR VPWR o[8] sky130_fd_sc_hd__buf_2
XFILLER_160_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput384 net384 VGND VGND VPWR VPWR o[9] sky130_fd_sc_hd__buf_2
Xfanout1009 net1010 VGND VGND VPWR VPWR net1009 sky130_fd_sc_hd__buf_6
XFILLER_120_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_61_1 pp_row61_17 pp_row61_18 pp_row61_19 VGND VGND VPWR VPWR c$548 s$549
+ sky130_fd_sc_hd__fa_1
Xdadda_fa_1_54_0 pp_row54_5 pp_row54_6 pp_row54_7 VGND VGND VPWR VPWR c$420 s$421
+ sky130_fd_sc_hd__fa_1
XFILLER_167_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1409 t$5125 net1487 VGND VGND VPWR VPWR booth_b20_m16 sky130_fd_sc_hd__xor2_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_116_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_116_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_30_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_90_3 s$1811 s$1813 s$1815 VGND VGND VPWR VPWR c$2564 s$2565 sky130_fd_sc_hd__fa_1
XFILLER_136_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_83_2 c$1720 s$1723 s$1725 VGND VGND VPWR VPWR c$2506 s$2507 sky130_fd_sc_hd__fa_1
XFILLER_174_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_76_1 c$1630 c$1632 c$1634 VGND VGND VPWR VPWR c$2448 s$2449 sky130_fd_sc_hd__fa_1
XFILLER_151_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_53_0 c$3604 c$3606 s$3609 VGND VGND VPWR VPWR c$4002 s$4003 sky130_fd_sc_hd__fa_1
Xfanout1510 net127 VGND VGND VPWR VPWR net1510 sky130_fd_sc_hd__buf_6
Xdadda_fa_3_69_0 s$707 c$1542 c$1544 VGND VGND VPWR VPWR c$2390 s$2391 sky130_fd_sc_hd__fa_1
Xfanout1521 net1522 VGND VGND VPWR VPWR net1521 sky130_fd_sc_hd__buf_4
Xfanout1532 net1534 VGND VGND VPWR VPWR net1532 sky130_fd_sc_hd__buf_4
Xfanout1543 net1546 VGND VGND VPWR VPWR net1543 sky130_fd_sc_hd__buf_4
XFILLER_120_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4002 t$6450 net1287 VGND VGND VPWR VPWR booth_b58_m11 sky130_fd_sc_hd__xor2_1
Xfanout1554 net1559 VGND VGND VPWR VPWR net1554 sky130_fd_sc_hd__buf_2
XU$$4013 net1159 net451 net1152 net724 VGND VGND VPWR VPWR t$6456 sky130_fd_sc_hd__a22o_1
Xfanout1565 net1567 VGND VGND VPWR VPWR net1565 sky130_fd_sc_hd__clkbuf_8
XFILLER_120_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4024 t$6461 net1285 VGND VGND VPWR VPWR booth_b58_m22 sky130_fd_sc_hd__xor2_1
Xfanout1576 net1577 VGND VGND VPWR VPWR net1576 sky130_fd_sc_hd__buf_6
XU$$4035 net1061 net454 net1052 net727 VGND VGND VPWR VPWR t$6467 sky130_fd_sc_hd__a22o_1
Xfanout1587 net1594 VGND VGND VPWR VPWR net1587 sky130_fd_sc_hd__buf_2
XU$$4046 t$6472 net1287 VGND VGND VPWR VPWR booth_b58_m33 sky130_fd_sc_hd__xor2_1
XFILLER_24_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3301 t$6092 net1339 VGND VGND VPWR VPWR booth_b48_m3 sky130_fd_sc_hd__xor2_1
Xfanout1598 net117 VGND VGND VPWR VPWR net1598 sky130_fd_sc_hd__buf_4
XU$$4057 net953 net457 net945 net730 VGND VGND VPWR VPWR t$6478 sky130_fd_sc_hd__a22o_1
XU$$3312 net1510 net500 net1501 net773 VGND VGND VPWR VPWR t$6098 sky130_fd_sc_hd__a22o_1
X_1050_ clknet_leaf_57_clk booth_b6_m1 VGND VGND VPWR VPWR pp_row7_3 sky130_fd_sc_hd__dfxtp_1
XU$$4068 t$6483 net1289 VGND VGND VPWR VPWR booth_b58_m44 sky130_fd_sc_hd__xor2_1
XU$$3323 t$6103 net1339 VGND VGND VPWR VPWR booth_b48_m14 sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_112_2 s$2733 s$2735 s$2737 VGND VGND VPWR VPWR c$3366 s$3367 sky130_fd_sc_hd__fa_1
XU$$3334 net1137 net497 net1121 net770 VGND VGND VPWR VPWR t$6109 sky130_fd_sc_hd__a22o_1
XU$$4079 net1685 net453 net1659 net726 VGND VGND VPWR VPWR t$6489 sky130_fd_sc_hd__a22o_1
XU$$2600 net1534 net557 net1778 net830 VGND VGND VPWR VPWR t$5733 sky130_fd_sc_hd__a22o_1
XU$$3345 t$6114 net1338 VGND VGND VPWR VPWR booth_b48_m25 sky130_fd_sc_hd__xor2_1
XFILLER_18_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_911 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3356 net1027 net494 net1019 net767 VGND VGND VPWR VPWR t$6120 sky130_fd_sc_hd__a22o_1
XU$$2611 net1228 net544 net1123 net817 VGND VGND VPWR VPWR t$5740 sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_105_1 c$2674 c$2676 s$2679 VGND VGND VPWR VPWR c$3322 s$3323 sky130_fd_sc_hd__fa_1
XU$$3367 t$6125 net1341 VGND VGND VPWR VPWR booth_b48_m36 sky130_fd_sc_hd__xor2_1
XU$$2622 t$5745 net1394 VGND VGND VPWR VPWR booth_b38_m6 sky130_fd_sc_hd__xor2_1
XFILLER_20_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2633 net1217 net549 net1206 net822 VGND VGND VPWR VPWR t$5751 sky130_fd_sc_hd__a22o_1
XFILLER_18_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3378 net1751 net499 net1743 net772 VGND VGND VPWR VPWR t$6131 sky130_fd_sc_hd__a22o_1
XU$$2644 t$5756 net1399 VGND VGND VPWR VPWR booth_b38_m17 sky130_fd_sc_hd__xor2_1
XU$$3389 t$6136 net1346 VGND VGND VPWR VPWR booth_b48_m47 sky130_fd_sc_hd__xor2_1
XU$$1910 t$5380 net1463 VGND VGND VPWR VPWR booth_b26_m61 sky130_fd_sc_hd__xor2_1
XFILLER_62_955 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2655 net1099 net544 net1093 net817 VGND VGND VPWR VPWR t$5762 sky130_fd_sc_hd__a22o_1
XU$$2666 t$5767 net1399 VGND VGND VPWR VPWR booth_b38_m28 sky130_fd_sc_hd__xor2_1
XU$$1921 net1453 notblock$5385\[1\] VGND VGND VPWR VPWR t$5386 sky130_fd_sc_hd__and2_1
XU$$2677 net994 net546 net984 net819 VGND VGND VPWR VPWR t$5773 sky130_fd_sc_hd__a22o_1
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1932 net936 net587 net1676 net860 VGND VGND VPWR VPWR t$5393 sky130_fd_sc_hd__a22o_1
XU$$2688 t$5778 net1396 VGND VGND VPWR VPWR booth_b38_m39 sky130_fd_sc_hd__xor2_1
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1943 t$5398 net1451 VGND VGND VPWR VPWR booth_b28_m9 sky130_fd_sc_hd__xor2_1
XU$$2699 net1722 net545 net1713 net818 VGND VGND VPWR VPWR t$5784 sky130_fd_sc_hd__a22o_1
XU$$1954 net1173 net584 net1164 net857 VGND VGND VPWR VPWR t$5404 sky130_fd_sc_hd__a22o_1
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1965 t$5409 net1448 VGND VGND VPWR VPWR booth_b28_m20 sky130_fd_sc_hd__xor2_1
XFILLER_178_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1976 net1074 net587 net1066 net860 VGND VGND VPWR VPWR t$5415 sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_107_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_107_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_15_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1952_ clknet_leaf_66_clk booth_b8_m46 VGND VGND VPWR VPWR pp_row54_4 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_7_126_0 s$3899 c$4146 s$4149 VGND VGND VPWR VPWR c$4404 s$4405 sky130_fd_sc_hd__fa_2
XU$$1987 t$5420 net1452 VGND VGND VPWR VPWR booth_b28_m31 sky130_fd_sc_hd__xor2_1
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1998 net969 net588 net961 net861 VGND VGND VPWR VPWR t$5426 sky130_fd_sc_hd__a22o_1
XFILLER_187_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0903_ clknet_leaf_103_clk booth_b34_m62 VGND VGND VPWR VPWR pp_row96_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_147_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1883_ clknet_leaf_134_clk booth_b58_m49 VGND VGND VPWR VPWR pp_row107_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_147_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0834_ clknet_leaf_106_clk booth_b60_m32 VGND VGND VPWR VPWR pp_row92_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_128_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0765_ clknet_leaf_152_clk booth_b62_m27 VGND VGND VPWR VPWR pp_row89_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_115_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0696_ clknet_leaf_175_clk booth_b26_m61 VGND VGND VPWR VPWR pp_row87_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_143_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2435_ clknet_leaf_75_clk booth_b50_m17 VGND VGND VPWR VPWR pp_row67_25 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_71_0 s$171 c$708 c$710 VGND VGND VPWR VPWR c$1578 s$1579 sky130_fd_sc_hd__fa_1
XFILLER_9_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2366_ clknet_leaf_98_clk booth_b60_m5 VGND VGND VPWR VPWR pp_row65_30 sky130_fd_sc_hd__dfxtp_1
XFILLER_111_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$606 final_adder.p_new$618 final_adder.p_new$610 VGND VGND VPWR VPWR
+ final_adder.p_new$734 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$617 final_adder.p_new$620 final_adder.g_new$629 final_adder.g_new$621
+ VGND VGND VPWR VPWR final_adder.g_new$745 sky130_fd_sc_hd__a21o_1
XFILLER_111_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1317_ clknet_leaf_247_clk booth_b2_m27 VGND VGND VPWR VPWR pp_row29_1 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$628 final_adder.p_new$652 final_adder.p_new$636 VGND VGND VPWR VPWR
+ final_adder.p_new$756 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$639 final_adder.p_new$646 final_adder.g_new$663 final_adder.g_new$647
+ VGND VGND VPWR VPWR final_adder.g_new$767 sky130_fd_sc_hd__a21o_1
X_2297_ clknet_leaf_199_clk booth_b0_m64 VGND VGND VPWR VPWR pp_row64_0 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_5_25__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_5_25__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_38_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1248_ clknet_leaf_10_clk booth_b4_m21 VGND VGND VPWR VPWR pp_row25_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_65_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$50 net1108 net448 net1100 net690 VGND VGND VPWR VPWR t$4432 sky130_fd_sc_hd__a22o_1
XU$$61 t$4437 net1568 VGND VGND VPWR VPWR booth_b0_m27 sky130_fd_sc_hd__xor2_1
XFILLER_65_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$72 net1000 net447 net992 net689 VGND VGND VPWR VPWR t$4443 sky130_fd_sc_hd__a22o_1
XU$$83 t$4448 net1569 VGND VGND VPWR VPWR booth_b0_m38 sky130_fd_sc_hd__xor2_1
X_1179_ clknet_leaf_49_clk booth_b12_m8 VGND VGND VPWR VPWR pp_row20_6 sky130_fd_sc_hd__dfxtp_1
XU$$94 net1729 net445 net1720 net687 VGND VGND VPWR VPWR t$4454 sky130_fd_sc_hd__a22o_1
XFILLER_80_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3890 net1094 net462 net1085 net735 VGND VGND VPWR VPWR t$6393 sky130_fd_sc_hd__a22o_1
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_30 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_41 net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_52 net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_63 net412 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_74 net458 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_85 net517 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_96 net534 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdadda_fa_4_93_1 c$2578 c$2580 s$2583 VGND VGND VPWR VPWR c$3250 s$3251 sky130_fd_sc_hd__fa_1
XFILLER_193_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_7_70_0 s$3679 c$4034 s$4037 VGND VGND VPWR VPWR c$4292 s$4293 sky130_fd_sc_hd__fa_1
XFILLER_192_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_86_0 s$1769 c$2518 c$2520 VGND VGND VPWR VPWR c$3206 s$3207 sky130_fd_sc_hd__fa_1
Xdadda_fa_3_107_3 pp_row107_12 c$1966 c$1968 VGND VGND VPWR VPWR c$2700 s$2701 sky130_fd_sc_hd__fa_1
XFILLER_97_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1206 net1649 net650 net1641 net923 VGND VGND VPWR VPWR t$5021 sky130_fd_sc_hd__a22o_1
XU$$1217 t$5026 net1012 VGND VGND VPWR VPWR booth_b16_m57 sky130_fd_sc_hd__xor2_1
XU$$1228 net1535 net649 net1527 net922 VGND VGND VPWR VPWR t$5032 sky130_fd_sc_hd__a22o_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1239 net1757 net637 net1228 net910 VGND VGND VPWR VPWR t$5039 sky130_fd_sc_hd__a22o_1
XFILLER_43_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_857 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1000 final_adder.$signal$1129 final_adder.g_new$1070 VGND VGND VPWR
+ VPWR net317 sky130_fd_sc_hd__xor2_2
XFILLER_156_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$1011 final_adder.$signal$103 final_adder.g_new$945 VGND VGND VPWR
+ VPWR net330 sky130_fd_sc_hd__xor2_2
XFILLER_8_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1022 final_adder.$signal$1151 final_adder.g_new$1059 VGND VGND VPWR
+ VPWR net342 sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$1033 final_adder.$signal$1162 final_adder.g_new$1019 VGND VGND VPWR
+ VPWR net354 sky130_fd_sc_hd__xor2_2
XFILLER_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$1044 final_adder.$signal$1173 final_adder.g_new$1048 VGND VGND VPWR
+ VPWR net366 sky130_fd_sc_hd__xor2_2
XFILLER_184_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$1055 final_adder.$signal$1184 final_adder.g_new$997 VGND VGND VPWR
+ VPWR net378 sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$1066 final_adder.$signal$1195 final_adder.g_new$1037 VGND VGND VPWR
+ VPWR net263 sky130_fd_sc_hd__xor2_1
XFILLER_171_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$1077 final_adder.$signal$1206 final_adder.g_new$975 VGND VGND VPWR
+ VPWR net275 sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$1088 final_adder.$signal$1217 final_adder.g_new$1026 VGND VGND VPWR
+ VPWR net287 sky130_fd_sc_hd__xor2_2
X_0550_ clknet_leaf_172_clk booth_b50_m31 VGND VGND VPWR VPWR pp_row81_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0481_ clknet_leaf_205_clk booth_b30_m49 VGND VGND VPWR VPWR pp_row79_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_79_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2220_ clknet_leaf_215_clk booth_b60_m1 VGND VGND VPWR VPWR pp_row61_30 sky130_fd_sc_hd__dfxtp_1
XFILLER_97_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1340 net1342 VGND VGND VPWR VPWR net1340 sky130_fd_sc_hd__buf_6
XFILLER_39_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1351 net1352 VGND VGND VPWR VPWR net1351 sky130_fd_sc_hd__buf_6
Xfanout1362 net1363 VGND VGND VPWR VPWR net1362 sky130_fd_sc_hd__buf_6
X_2151_ clknet_leaf_215_clk booth_b2_m58 VGND VGND VPWR VPWR pp_row60_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_120_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_50_5 s$359 s$361 s$363 VGND VGND VPWR VPWR c$1336 s$1337 sky130_fd_sc_hd__fa_2
Xfanout1373 net1374 VGND VGND VPWR VPWR net1373 sky130_fd_sc_hd__buf_6
Xfanout1384 net36 VGND VGND VPWR VPWR net1384 sky130_fd_sc_hd__clkbuf_16
Xfanout1395 net33 VGND VGND VPWR VPWR net1395 sky130_fd_sc_hd__buf_6
X_1102_ clknet_leaf_14_clk booth_b0_m14 VGND VGND VPWR VPWR pp_row14_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_93_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_43_4 c$250 c$252 s$255 VGND VGND VPWR VPWR c$1250 s$1251 sky130_fd_sc_hd__fa_1
XU$$3120 net1684 net515 net1660 net788 VGND VGND VPWR VPWR t$5999 sky130_fd_sc_hd__a22o_1
X_2082_ clknet_leaf_86_clk booth_b4_m54 VGND VGND VPWR VPWR pp_row58_2 sky130_fd_sc_hd__dfxtp_1
XU$$3131 t$6004 net1364 VGND VGND VPWR VPWR booth_b44_m55 sky130_fd_sc_hd__xor2_1
Xdadda_ha_6_2_0 pp_row2_0 pp_row2_1 VGND VGND VPWR VPWR c$3900 s$3901 sky130_fd_sc_hd__ha_1
XU$$3142 net1558 net515 net1550 net788 VGND VGND VPWR VPWR t$6010 sky130_fd_sc_hd__a22o_1
XU$$3153 net1350 VGND VGND VPWR VPWR notblock$6015\[2\] sky130_fd_sc_hd__inv_1
X_1033_ clknet_leaf_60_clk net1278 VGND VGND VPWR VPWR pp_row4_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_36_3 pp_row36_14 pp_row36_15 pp_row36_16 VGND VGND VPWR VPWR c$1164 s$1165
+ sky130_fd_sc_hd__fa_1
XU$$3164 t$6022 net1348 VGND VGND VPWR VPWR booth_b46_m3 sky130_fd_sc_hd__xor2_1
XU$$3175 net1510 net505 net1501 net778 VGND VGND VPWR VPWR t$6028 sky130_fd_sc_hd__a22o_1
XU$$2430 t$5646 net1426 VGND VGND VPWR VPWR booth_b34_m47 sky130_fd_sc_hd__xor2_1
XU$$3186 t$6033 net1348 VGND VGND VPWR VPWR booth_b46_m14 sky130_fd_sc_hd__xor2_1
XU$$2441 net1639 net566 net1631 net839 VGND VGND VPWR VPWR t$5652 sky130_fd_sc_hd__a22o_1
XU$$2452 t$5657 net1428 VGND VGND VPWR VPWR booth_b34_m58 sky130_fd_sc_hd__xor2_1
XU$$3197 net1137 net505 net1121 net778 VGND VGND VPWR VPWR t$6039 sky130_fd_sc_hd__a22o_1
XU$$2463 net1534 net567 net1776 net840 VGND VGND VPWR VPWR t$5663 sky130_fd_sc_hd__a22o_1
XFILLER_34_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_29_2 pp_row29_6 pp_row29_7 pp_row29_8 VGND VGND VPWR VPWR c$1086 s$1087
+ sky130_fd_sc_hd__fa_1
XFILLER_22_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2474 net1232 net552 net1128 net825 VGND VGND VPWR VPWR t$5670 sky130_fd_sc_hd__a22o_1
XU$$2485 t$5675 net1403 VGND VGND VPWR VPWR booth_b36_m6 sky130_fd_sc_hd__xor2_1
XU$$1740 net1724 net609 net1715 net882 VGND VGND VPWR VPWR t$5294 sky130_fd_sc_hd__a22o_1
XU$$1751 t$5299 net1473 VGND VGND VPWR VPWR booth_b24_m50 sky130_fd_sc_hd__xor2_1
XU$$2496 net1213 net551 net1202 net824 VGND VGND VPWR VPWR t$5681 sky130_fd_sc_hd__a22o_1
XU$$1762 net1613 net608 net1605 net881 VGND VGND VPWR VPWR t$5305 sky130_fd_sc_hd__a22o_1
XFILLER_22_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1773 t$5310 net1471 VGND VGND VPWR VPWR booth_b24_m61 sky130_fd_sc_hd__xor2_1
XU$$1784 net1463 notblock$5315\[1\] VGND VGND VPWR VPWR t$5316 sky130_fd_sc_hd__and2_1
XFILLER_50_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1795 net932 net593 net1671 net866 VGND VGND VPWR VPWR t$5323 sky130_fd_sc_hd__a22o_1
XFILLER_188_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1935_ clknet_leaf_70_clk booth_b36_m17 VGND VGND VPWR VPWR pp_row53_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_159_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1866_ clknet_leaf_67_clk booth_b22_m29 VGND VGND VPWR VPWR pp_row51_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_174_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput50 a[54] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_2
XFILLER_135_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0817_ clknet_leaf_111_clk booth_b32_m60 VGND VGND VPWR VPWR pp_row92_3 sky130_fd_sc_hd__dfxtp_1
Xinput61 a[6] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_2
XFILLER_128_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput72 b[16] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_8
XFILLER_174_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_0_76_0_1895 VGND VGND VPWR VPWR net1895 dadda_fa_0_76_0_1895/LO sky130_fd_sc_hd__conb_1
X_1797_ clknet_leaf_218_clk booth_b6_m43 VGND VGND VPWR VPWR pp_row49_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput83 b[26] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__buf_6
Xinput94 b[36] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_4
XFILLER_104_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_860 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0748_ clknet_leaf_160_clk booth_b30_m59 VGND VGND VPWR VPWR pp_row89_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_89_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0679_ clknet_leaf_179_clk booth_b40_m46 VGND VGND VPWR VPWR pp_row86_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_130_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4_1802 VGND VGND VPWR VPWR U$$4_1802/HI net1802 sky130_fd_sc_hd__conb_1
X_2418_ clknet_leaf_145_clk booth_b18_m49 VGND VGND VPWR VPWR pp_row67_9 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$403 final_adder.p_new$404 final_adder.g_new$409 final_adder.g_new$405
+ VGND VGND VPWR VPWR final_adder.g_new$531 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$414 final_adder.p_new$420 final_adder.p_new$416 VGND VGND VPWR VPWR
+ final_adder.p_new$542 sky130_fd_sc_hd__and2_1
X_2349_ clknet_leaf_88_clk booth_b28_m37 VGND VGND VPWR VPWR pp_row65_14 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$425 final_adder.p_new$426 final_adder.g_new$431 final_adder.g_new$427
+ VGND VGND VPWR VPWR final_adder.g_new$553 sky130_fd_sc_hd__a21o_1
XTAP_3707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$436 final_adder.p_new$442 final_adder.p_new$438 VGND VGND VPWR VPWR
+ final_adder.p_new$564 sky130_fd_sc_hd__and2_1
XTAP_3718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$447 final_adder.p_new$448 final_adder.g_new$453 final_adder.g_new$449
+ VGND VGND VPWR VPWR final_adder.g_new$575 sky130_fd_sc_hd__a21o_1
XTAP_3729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$458 final_adder.p_new$464 final_adder.p_new$460 VGND VGND VPWR VPWR
+ final_adder.p_new$586 sky130_fd_sc_hd__and2_1
XU$$308 net1194 net528 net1175 net801 VGND VGND VPWR VPWR t$4563 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$469 final_adder.p_new$470 final_adder.g_new$475 final_adder.g_new$471
+ VGND VGND VPWR VPWR final_adder.g_new$597 sky130_fd_sc_hd__a21o_1
XFILLER_42_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$319 t$4568 net1279 VGND VGND VPWR VPWR booth_b4_m19 sky130_fd_sc_hd__xor2_1
XFILLER_38_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_857 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_112_1 pp_row112_3 pp_row112_4 pp_row112_5 VGND VGND VPWR VPWR c$2734 s$2735
+ sky130_fd_sc_hd__fa_1
XFILLER_153_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_105_0 pp_row105_6 pp_row105_7 pp_row105_8 VGND VGND VPWR VPWR c$2678 s$2679
+ sky130_fd_sc_hd__fa_1
XFILLER_181_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_53_3 s$1367 s$1369 s$1371 VGND VGND VPWR VPWR c$2268 s$2269 sky130_fd_sc_hd__fa_1
XFILLER_94_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_0_69_3 pp_row69_9 pp_row69_10 pp_row69_11 VGND VGND VPWR VPWR c$150 s$151
+ sky130_fd_sc_hd__fa_1
XFILLER_169_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_46_2 c$1276 s$1279 s$1281 VGND VGND VPWR VPWR c$2210 s$2211 sky130_fd_sc_hd__fa_1
XFILLER_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$970 final_adder.$signal$1099 final_adder.g_new$1085 VGND VGND VPWR
+ VPWR net384 sky130_fd_sc_hd__xor2_2
XFILLER_180_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$820 t$4823 net1417 VGND VGND VPWR VPWR booth_b10_m64 sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_39_1 c$1186 c$1188 c$1190 VGND VGND VPWR VPWR c$2152 s$2153 sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$981 final_adder.$signal$1110 final_adder.g_new$863 VGND VGND VPWR
+ VPWR net297 sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$992 final_adder.$signal$1121 final_adder.g_new$1074 VGND VGND VPWR
+ VPWR net309 sky130_fd_sc_hd__xor2_2
XU$$831 t$4830 net1312 VGND VGND VPWR VPWR booth_b12_m1 sky130_fd_sc_hd__xor2_1
XFILLER_28_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_730 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$842 net1523 net396 net1515 net662 VGND VGND VPWR VPWR t$4836 sky130_fd_sc_hd__a22o_1
XU$$853 t$4841 net1310 VGND VGND VPWR VPWR booth_b12_m12 sky130_fd_sc_hd__xor2_1
Xdadda_fa_6_16_0 c$3456 c$3458 s$3461 VGND VGND VPWR VPWR c$3928 s$3929 sky130_fd_sc_hd__fa_1
XU$$1003 net1143 net387 net1133 net653 VGND VGND VPWR VPWR t$4918 sky130_fd_sc_hd__a22o_1
XU$$864 net1146 net393 net1138 net659 VGND VGND VPWR VPWR t$4847 sky130_fd_sc_hd__a22o_1
XU$$1014 t$4923 net1185 VGND VGND VPWR VPWR booth_b14_m24 sky130_fd_sc_hd__xor2_1
XU$$875 t$4852 net1313 VGND VGND VPWR VPWR booth_b12_m23 sky130_fd_sc_hd__xor2_1
XU$$886 net1047 net394 net1039 net660 VGND VGND VPWR VPWR t$4858 sky130_fd_sc_hd__a22o_1
XU$$1025 net1039 net386 net1023 net652 VGND VGND VPWR VPWR t$4929 sky130_fd_sc_hd__a22o_1
XFILLER_32_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$897 t$4863 net1311 VGND VGND VPWR VPWR booth_b12_m34 sky130_fd_sc_hd__xor2_1
XU$$1036 t$4934 net1184 VGND VGND VPWR VPWR booth_b14_m35 sky130_fd_sc_hd__xor2_1
XFILLER_189_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1047 net928 net388 net1749 net654 VGND VGND VPWR VPWR t$4940 sky130_fd_sc_hd__a22o_1
XFILLER_32_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1058 t$4945 net1190 VGND VGND VPWR VPWR booth_b14_m46 sky130_fd_sc_hd__xor2_1
XFILLER_188_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1069 net1649 net391 net1641 net657 VGND VGND VPWR VPWR t$4951 sky130_fd_sc_hd__a22o_1
XFILLER_176_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1720_ clknet_leaf_22_clk booth_b24_m22 VGND VGND VPWR VPWR pp_row46_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_11_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1651_ clknet_leaf_239_clk booth_b42_m1 VGND VGND VPWR VPWR pp_row43_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0602_ clknet_leaf_174_clk booth_b44_m39 VGND VGND VPWR VPWR pp_row83_13 sky130_fd_sc_hd__dfxtp_1
X_1582_ clknet_leaf_242_clk booth_b12_m29 VGND VGND VPWR VPWR pp_row41_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_171_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0533_ clknet_leaf_131_clk booth_b52_m64 VGND VGND VPWR VPWR pp_row116_1 sky130_fd_sc_hd__dfxtp_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0464_ clknet_leaf_206_clk booth_b54_m24 VGND VGND VPWR VPWR pp_row78_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_79_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2203_ clknet_leaf_88_clk booth_b30_m31 VGND VGND VPWR VPWR pp_row61_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_67_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0395_ clknet_leaf_192_clk booth_b38_m38 VGND VGND VPWR VPWR pp_row76_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1170 net1172 VGND VGND VPWR VPWR net1170 sky130_fd_sc_hd__buf_6
Xfanout1181 net1182 VGND VGND VPWR VPWR net1181 sky130_fd_sc_hd__buf_4
XFILLER_187_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1192 net1193 VGND VGND VPWR VPWR net1192 sky130_fd_sc_hd__buf_4
X_2134_ clknet_leaf_27_clk booth_b34_m25 VGND VGND VPWR VPWR pp_row59_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_82_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_41_1 pp_row41_14 pp_row41_15 pp_row41_16 VGND VGND VPWR VPWR c$1220 s$1221
+ sky130_fd_sc_hd__fa_1
XFILLER_187_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2065_ clknet_leaf_34_clk booth_b32_m25 VGND VGND VPWR VPWR pp_row57_16 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_34_0 pp_row34_2 pp_row34_3 pp_row34_4 VGND VGND VPWR VPWR c$1134 s$1135
+ sky130_fd_sc_hd__fa_1
X_1016_ clknet_leaf_120_clk booth_b40_m62 VGND VGND VPWR VPWR pp_row102_2 sky130_fd_sc_hd__dfxtp_1
XU$$2260 net1024 sel_0$5527 net1016 sel_1$5528 VGND VGND VPWR VPWR t$5560 sky130_fd_sc_hd__a22o_1
XFILLER_179_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2271 t$5565 net1437 VGND VGND VPWR VPWR booth_b32_m36 sky130_fd_sc_hd__xor2_1
XFILLER_35_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2282 net1746 net570 net1738 net843 VGND VGND VPWR VPWR t$5571 sky130_fd_sc_hd__a22o_1
XFILLER_90_891 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2293 t$5576 net1434 VGND VGND VPWR VPWR booth_b32_m47 sky130_fd_sc_hd__xor2_1
XU$$1570 t$5207 net1478 VGND VGND VPWR VPWR booth_b22_m28 sky130_fd_sc_hd__xor2_1
XFILLER_22_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1581 net992 net613 net987 net886 VGND VGND VPWR VPWR t$5213 sky130_fd_sc_hd__a22o_1
XU$$1592 t$5218 net1477 VGND VGND VPWR VPWR booth_b22_m39 sky130_fd_sc_hd__xor2_1
XFILLER_50_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1918_ clknet_leaf_81_clk booth_b4_m49 VGND VGND VPWR VPWR pp_row53_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_136_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1849_ clknet_leaf_25_clk booth_b48_m2 VGND VGND VPWR VPWR pp_row50_24 sky130_fd_sc_hd__dfxtp_1
XFILLER_191_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_86_3 pp_row86_9 pp_row86_10 pp_row86_11 VGND VGND VPWR VPWR c$984 s$985
+ sky130_fd_sc_hd__fa_1
XFILLER_89_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_63_2 s$2345 s$2347 s$2349 VGND VGND VPWR VPWR c$3072 s$3073 sky130_fd_sc_hd__fa_1
Xdadda_fa_1_79_2 pp_row79_6 pp_row79_7 pp_row79_8 VGND VGND VPWR VPWR c$874 s$875
+ sky130_fd_sc_hd__fa_1
XFILLER_58_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_56_1 c$2282 c$2284 s$2287 VGND VGND VPWR VPWR c$3028 s$3029 sky130_fd_sc_hd__fa_1
XTAP_4205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$200 final_adder.$signal$111 final_adder.$signal$113 VGND VGND VPWR
+ VPWR final_adder.p_new$328 sky130_fd_sc_hd__and2_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_96_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_96_clk sky130_fd_sc_hd__clkbuf_16
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_33_0 s$3531 c$3960 s$3963 VGND VGND VPWR VPWR c$4218 s$4219 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$211 final_adder.$signal$1135 final_adder.$signal$90 final_adder.$signal$92
+ VGND VGND VPWR VPWR final_adder.g_new$339 sky130_fd_sc_hd__a21o_1
XTAP_4238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_49_0 s$1325 c$2222 c$2224 VGND VGND VPWR VPWR c$2984 s$2985 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$222 final_adder.$signal$1122 final_adder.$signal$1123 VGND VGND VPWR
+ VPWR final_adder.p_new$350 sky130_fd_sc_hd__and2_1
XTAP_3504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$233 final_adder.$signal$1113 final_adder.$signal$46 final_adder.$signal$48
+ VGND VGND VPWR VPWR final_adder.g_new$361 sky130_fd_sc_hd__a21o_1
XTAP_4249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$244 final_adder.$signal$1100 final_adder.$signal$1101 VGND VGND VPWR
+ VPWR final_adder.p_new$372 sky130_fd_sc_hd__and2_1
XFILLER_18_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$255 final_adder.$signal$1091 final_adder.$signal final_adder.$signal$4
+ VGND VGND VPWR VPWR final_adder.g_new$383 sky130_fd_sc_hd__a21o_4
XTAP_3526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$105 t$4459 net1576 VGND VGND VPWR VPWR booth_b0_m49 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$266 final_adder.p_new$268 final_adder.p_new$266 VGND VGND VPWR VPWR
+ final_adder.p_new$394 sky130_fd_sc_hd__and2_1
XTAP_3548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$116 net1623 net449 net1619 net691 VGND VGND VPWR VPWR t$4465 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$277 final_adder.p_new$276 final_adder.g_new$279 final_adder.g_new$277
+ VGND VGND VPWR VPWR final_adder.g_new$405 sky130_fd_sc_hd__a21o_1
XFILLER_57_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4429_1835 VGND VGND VPWR VPWR U$$4429_1835/HI net1835 sky130_fd_sc_hd__conb_1
XU$$127 t$4470 net1572 VGND VGND VPWR VPWR booth_b0_m60 sky130_fd_sc_hd__xor2_1
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$288 final_adder.p_new$290 final_adder.p_new$288 VGND VGND VPWR VPWR
+ final_adder.p_new$416 sky130_fd_sc_hd__and2_1
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$138 net23 VGND VGND VPWR VPWR notblock$4475\[1\] sky130_fd_sc_hd__inv_1
Xfinal_adder.U$$299 final_adder.p_new$298 final_adder.g_new$301 final_adder.g_new$299
+ VGND VGND VPWR VPWR final_adder.g_new$427 sky130_fd_sc_hd__a21o_1
XU$$149 net1035 net624 net937 net897 VGND VGND VPWR VPWR t$4482 sky130_fd_sc_hd__a22o_1
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_20_clk clknet_5_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_193_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_74_1 pp_row74_3 pp_row74_4 pp_row74_5 VGND VGND VPWR VPWR c$188 s$189
+ sky130_fd_sc_hd__fa_1
XFILLER_95_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput240 c[85] VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_3_51_0 s$383 c$1326 c$1328 VGND VGND VPWR VPWR c$2246 s$2247 sky130_fd_sc_hd__fa_2
Xinput251 c[95] VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_87_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_87_clk sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_0_67_0 pp_row67_0 pp_row67_1 pp_row67_2 VGND VGND VPWR VPWR c$120 s$121
+ sky130_fd_sc_hd__fa_1
X_0180_ clknet_leaf_197_clk net222 VGND VGND VPWR VPWR pp_row69_31 sky130_fd_sc_hd__dfxtp_2
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_1040 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$650 net1698 net416 net1690 net682 VGND VGND VPWR VPWR t$4737 sky130_fd_sc_hd__a22o_1
XU$$661 t$4742 net1237 VGND VGND VPWR VPWR booth_b8_m53 sky130_fd_sc_hd__xor2_1
XFILLER_63_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$672 net1590 net416 net1582 net682 VGND VGND VPWR VPWR t$4748 sky130_fd_sc_hd__a22o_1
XFILLER_17_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$683 t$4753 net1238 VGND VGND VPWR VPWR booth_b8_m64 sky130_fd_sc_hd__xor2_1
XFILLER_44_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$694 t$4760 net1414 VGND VGND VPWR VPWR booth_b10_m1 sky130_fd_sc_hd__xor2_1
XFILLER_56_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_11_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1703_ clknet_leaf_23_clk booth_b42_m3 VGND VGND VPWR VPWR pp_row45_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_117_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_96_2 pp_row96_8 pp_row96_9 pp_row96_10 VGND VGND VPWR VPWR c$1882 s$1883
+ sky130_fd_sc_hd__fa_1
X_1634_ clknet_leaf_239_clk booth_b12_m31 VGND VGND VPWR VPWR pp_row43_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_126_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_73_1 s$3129 s$3131 s$3133 VGND VGND VPWR VPWR c$3690 s$3691 sky130_fd_sc_hd__fa_2
Xdadda_fa_2_89_1 pp_row89_15 pp_row89_16 pp_row89_17 VGND VGND VPWR VPWR c$1796 s$1797
+ sky130_fd_sc_hd__fa_1
XFILLER_193_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1565_ clknet_leaf_8_clk booth_b26_m14 VGND VGND VPWR VPWR pp_row40_13 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_66_0 c$3080 c$3082 c$3084 VGND VGND VPWR VPWR c$3660 s$3661 sky130_fd_sc_hd__fa_1
Xfanout407 net408 VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__buf_6
XFILLER_59_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout418 net421 VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__clkbuf_8
XFILLER_113_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0516_ clknet_leaf_160_clk booth_b40_m40 VGND VGND VPWR VPWR pp_row80_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_98_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout429 net430 VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__buf_4
XFILLER_154_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1496_ clknet_leaf_45_clk booth_b28_m9 VGND VGND VPWR VPWR pp_row37_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_86_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0447_ clknet_leaf_206_clk booth_b22_m56 VGND VGND VPWR VPWR pp_row78_5 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_65_8 s$101 s$103 s$105 VGND VGND VPWR VPWR c$634 s$635 sky130_fd_sc_hd__fa_1
Xclkbuf_leaf_78_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_78_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_95_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_58_7 c$18 c$20 c$22 VGND VGND VPWR VPWR c$506 s$507 sky130_fd_sc_hd__fa_1
XFILLER_27_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0378_ clknet_leaf_200_clk booth_b64_m11 VGND VGND VPWR VPWR pp_row75_27 sky130_fd_sc_hd__dfxtp_1
X_2117_ clknet_leaf_224_clk booth_b2_m57 VGND VGND VPWR VPWR pp_row59_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2048_ clknet_leaf_38_clk booth_b4_m53 VGND VGND VPWR VPWR pp_row57_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_82_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_5_0 pp_row5_2 pp_row5_3 c$3416 VGND VGND VPWR VPWR c$3906 s$3907 sky130_fd_sc_hd__fa_1
XFILLER_120_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2090 t$5473 net1440 VGND VGND VPWR VPWR booth_b30_m14 sky130_fd_sc_hd__xor2_1
XFILLER_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_91_1 pp_row91_3 pp_row91_4 pp_row91_5 VGND VGND VPWR VPWR c$1028 s$1029
+ sky130_fd_sc_hd__fa_1
XFILLER_151_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_84_0 net1898 pp_row84_1 pp_row84_2 VGND VGND VPWR VPWR c$952 s$953 sky130_fd_sc_hd__fa_1
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout930 net931 VGND VGND VPWR VPWR net930 sky130_fd_sc_hd__buf_4
XFILLER_104_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout941 net947 VGND VGND VPWR VPWR net941 sky130_fd_sc_hd__buf_6
Xfanout952 net96 VGND VGND VPWR VPWR net952 sky130_fd_sc_hd__buf_6
XTAP_4002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout963 net95 VGND VGND VPWR VPWR net963 sky130_fd_sc_hd__buf_4
XTAP_4013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_69_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_69_clk sky130_fd_sc_hd__clkbuf_16
XU$$4409 t$6658 net1825 VGND VGND VPWR VPWR booth_b64_m9 sky130_fd_sc_hd__xor2_1
Xfanout974 net981 VGND VGND VPWR VPWR net974 sky130_fd_sc_hd__buf_6
XTAP_4024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout985 net986 VGND VGND VPWR VPWR net985 sky130_fd_sc_hd__buf_4
XTAP_4035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout996 net997 VGND VGND VPWR VPWR net996 sky130_fd_sc_hd__buf_4
XFILLER_46_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3708 t$6300 net1304 VGND VGND VPWR VPWR booth_b54_m1 sky130_fd_sc_hd__xor2_1
XFILLER_57_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3719 net1522 net471 net1514 net744 VGND VGND VPWR VPWR t$6306 sky130_fd_sc_hd__a22o_1
XTAP_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_301 net414 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_312 net558 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_323 net629 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_334 net715 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_345 net841 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_356 net947 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_891 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_367 net1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_378 net1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_389 net1507 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_83_0 c$3724 c$3726 s$3729 VGND VGND VPWR VPWR c$4062 s$4063 sky130_fd_sc_hd__fa_1
XFILLER_186_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_99_0 pp_row99_15 pp_row99_16 c$1902 VGND VGND VPWR VPWR c$2630 s$2631
+ sky130_fd_sc_hd__fa_1
XFILLER_177_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1350_ clknet_leaf_246_clk booth_b30_m0 VGND VGND VPWR VPWR pp_row30_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_150_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0301_ clknet_leaf_227_clk booth_b40_m33 VGND VGND VPWR VPWR pp_row73_16 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_5_6__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_5_6__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_122_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1281_ clknet_leaf_250_clk booth_b4_m23 VGND VGND VPWR VPWR pp_row27_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0232_ clknet_leaf_151_clk booth_b38_m33 VGND VGND VPWR VPWR pp_row71_16 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_0_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_184_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$480 t$4650 net1250 VGND VGND VPWR VPWR booth_b6_m31 sky130_fd_sc_hd__xor2_1
XU$$491 net964 net426 net956 net708 VGND VGND VPWR VPWR t$4656 sky130_fd_sc_hd__a22o_1
XFILLER_51_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0996_ clknet_leaf_184_clk net130 VGND VGND VPWR VPWR pp_row100_16 sky130_fd_sc_hd__dfxtp_4
XFILLER_157_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1617_ clknet_leaf_164_clk booth_b62_m61 VGND VGND VPWR VPWR pp_row123_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_8_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1548_ clknet_leaf_19_clk booth_b38_m1 VGND VGND VPWR VPWR pp_row39_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_141_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_70_6 c$144 c$146 c$148 VGND VGND VPWR VPWR c$720 s$721 sky130_fd_sc_hd__fa_1
XFILLER_59_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_63_5 pp_row63_32 c$60 c$62 VGND VGND VPWR VPWR c$592 s$593 sky130_fd_sc_hd__fa_1
X_1479_ clknet_leaf_236_clk net186 VGND VGND VPWR VPWR pp_row36_20 sky130_fd_sc_hd__dfxtp_2
XFILLER_68_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_56_4 pp_row56_20 pp_row56_21 pp_row56_22 VGND VGND VPWR VPWR c$464 s$465
+ sky130_fd_sc_hd__fa_1
XFILLER_28_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_49_3 pp_row49_9 pp_row49_10 pp_row49_11 VGND VGND VPWR VPWR c$338 s$339
+ sky130_fd_sc_hd__fa_1
Xdadda_fa_4_26_2 s$2049 s$2051 s$2053 VGND VGND VPWR VPWR c$2850 s$2851 sky130_fd_sc_hd__fa_1
XFILLER_55_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_19_1 c$1986 c$1988 c$1990 VGND VGND VPWR VPWR c$2806 s$2807 sky130_fd_sc_hd__fa_1
XFILLER_42_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1703 net1705 VGND VGND VPWR VPWR net1703 sky130_fd_sc_hd__buf_4
Xfanout1714 net104 VGND VGND VPWR VPWR net1714 sky130_fd_sc_hd__buf_4
XFILLER_133_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1725 net1728 VGND VGND VPWR VPWR net1725 sky130_fd_sc_hd__clkbuf_4
XU$$4513_1877 VGND VGND VPWR VPWR U$$4513_1877/HI net1877 sky130_fd_sc_hd__conb_1
Xfanout1736 net102 VGND VGND VPWR VPWR net1736 sky130_fd_sc_hd__buf_6
Xfanout1747 net1752 VGND VGND VPWR VPWR net1747 sky130_fd_sc_hd__buf_6
XFILLER_172_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4206 net1726 net440 net1717 net722 VGND VGND VPWR VPWR t$6554 sky130_fd_sc_hd__a22o_1
Xfanout760 sel_1$6158 VGND VGND VPWR VPWR net760 sky130_fd_sc_hd__clkbuf_8
Xfanout771 net772 VGND VGND VPWR VPWR net771 sky130_fd_sc_hd__buf_4
XU$$4217 t$6559 net1270 VGND VGND VPWR VPWR booth_b60_m50 sky130_fd_sc_hd__xor2_1
Xfanout782 sel_1$6018 VGND VGND VPWR VPWR net782 sky130_fd_sc_hd__clkbuf_8
XFILLER_93_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4228 net1619 net439 net1610 net721 VGND VGND VPWR VPWR t$6565 sky130_fd_sc_hd__a22o_1
Xfanout793 sel_1$5878 VGND VGND VPWR VPWR net793 sky130_fd_sc_hd__buf_4
XU$$4239 t$6570 net1265 VGND VGND VPWR VPWR booth_b60_m61 sky130_fd_sc_hd__xor2_1
XU$$3505 net967 net485 net958 net758 VGND VGND VPWR VPWR t$6196 sky130_fd_sc_hd__a22o_1
XU$$3516 t$6201 net1334 VGND VGND VPWR VPWR booth_b50_m42 sky130_fd_sc_hd__xor2_1
XU$$3527 net1700 net490 net1693 net763 VGND VGND VPWR VPWR t$6207 sky130_fd_sc_hd__a22o_1
XTAP_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3538 t$6212 net1335 VGND VGND VPWR VPWR booth_b50_m53 sky130_fd_sc_hd__xor2_1
XFILLER_45_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2804 net1053 net538 net1045 net811 VGND VGND VPWR VPWR t$5838 sky130_fd_sc_hd__a22o_1
XU$$3549 net1591 net489 net1583 net762 VGND VGND VPWR VPWR t$6218 sky130_fd_sc_hd__a22o_1
XU$$2815 t$5843 net1377 VGND VGND VPWR VPWR booth_b40_m34 sky130_fd_sc_hd__xor2_1
XTAP_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2826 net943 net538 net927 net811 VGND VGND VPWR VPWR t$5849 sky130_fd_sc_hd__a22o_1
XTAP_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2837 t$5854 net1379 VGND VGND VPWR VPWR booth_b40_m45 sky130_fd_sc_hd__xor2_1
XFILLER_74_997 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_120 net655 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2848 net1659 net541 net1651 net814 VGND VGND VPWR VPWR t$5860 sky130_fd_sc_hd__a22o_1
XANTENNA_131 net710 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_21_1 pp_row21_3 pp_row21_4 pp_row21_5 VGND VGND VPWR VPWR c$2008 s$2009
+ sky130_fd_sc_hd__fa_1
XTAP_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2859 t$5865 net1382 VGND VGND VPWR VPWR booth_b40_m56 sky130_fd_sc_hd__xor2_1
XANTENNA_142 net765 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_153 net799 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_164 net879 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_175 net917 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_186 net972 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$545_1881 VGND VGND VPWR VPWR U$$545_1881/HI net1881 sky130_fd_sc_hd__conb_1
XFILLER_187_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_197 net1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0850_ clknet_leaf_109_clk booth_b50_m43 VGND VGND VPWR VPWR pp_row93_11 sky130_fd_sc_hd__dfxtp_1
X_0781_ clknet_leaf_140_clk booth_b48_m42 VGND VGND VPWR VPWR pp_row90_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_128_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3431_1793 VGND VGND VPWR VPWR U$$3431_1793/HI net1793 sky130_fd_sc_hd__conb_1
XFILLER_142_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2451_ clknet_leaf_92_clk booth_b14_m54 VGND VGND VPWR VPWR pp_row68_6 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_80_5 s$899 s$901 s$903 VGND VGND VPWR VPWR c$1696 s$1697 sky130_fd_sc_hd__fa_2
X_1402_ clknet_leaf_51_clk booth_b14_m19 VGND VGND VPWR VPWR pp_row33_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_64_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_73_4 s$767 s$769 s$771 VGND VGND VPWR VPWR c$1610 s$1611 sky130_fd_sc_hd__fa_1
X_2382_ clknet_leaf_83_clk booth_b22_m44 VGND VGND VPWR VPWR pp_row66_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1333_ clknet_leaf_0_clk booth_b0_m30 VGND VGND VPWR VPWR pp_row30_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_111_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_66_3 c$634 s$637 s$639 VGND VGND VPWR VPWR c$1524 s$1525 sky130_fd_sc_hd__fa_1
XFILLER_122_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_59_2 c$502 c$504 c$506 VGND VGND VPWR VPWR c$1438 s$1439 sky130_fd_sc_hd__fa_1
X_1264_ clknet_leaf_2_clk booth_b4_m22 VGND VGND VPWR VPWR pp_row26_2 sky130_fd_sc_hd__dfxtp_1
Xinput4 a[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_2
Xdadda_fa_5_36_1 s$2907 s$2909 s$2911 VGND VGND VPWR VPWR c$3542 s$3543 sky130_fd_sc_hd__fa_1
X_0215_ clknet_leaf_198_clk notsign$4684 VGND VGND VPWR VPWR pp_row71_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_37_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1195_ clknet_leaf_51_clk booth_b14_m7 VGND VGND VPWR VPWR pp_row21_7 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_29_0 c$2858 c$2860 c$2862 VGND VGND VPWR VPWR c$3512 s$3513 sky130_fd_sc_hd__fa_1
XFILLER_188_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_110_1 s$3351 s$3353 s$3355 VGND VGND VPWR VPWR c$3838 s$3839 sky130_fd_sc_hd__fa_1
X_0979_ clknet_leaf_184_clk net255 VGND VGND VPWR VPWR pp_row99_16 sky130_fd_sc_hd__dfxtp_4
XFILLER_192_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$2 c$4154 s$4157 VGND VGND VPWR VPWR final_adder.$signal$6 final_adder.$signal$1092
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_5_103_0 c$3302 c$3304 c$3306 VGND VGND VPWR VPWR c$3808 s$3809 sky130_fd_sc_hd__fa_1
XFILLER_119_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput330 net330 VGND VGND VPWR VPWR o[50] sky130_fd_sc_hd__buf_2
Xoutput341 net341 VGND VGND VPWR VPWR o[60] sky130_fd_sc_hd__buf_2
XFILLER_156_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput352 net352 VGND VGND VPWR VPWR o[70] sky130_fd_sc_hd__buf_2
XFILLER_121_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput363 net363 VGND VGND VPWR VPWR o[80] sky130_fd_sc_hd__buf_2
Xoutput374 net374 VGND VGND VPWR VPWR o[90] sky130_fd_sc_hd__buf_2
XFILLER_99_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_61_2 pp_row61_20 pp_row61_21 pp_row61_22 VGND VGND VPWR VPWR c$550 s$551
+ sky130_fd_sc_hd__fa_1
XFILLER_87_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_54_1 pp_row54_8 pp_row54_9 pp_row54_10 VGND VGND VPWR VPWR c$422 s$423
+ sky130_fd_sc_hd__fa_1
Xdadda_fa_4_31_0 s$1109 c$2078 c$2080 VGND VGND VPWR VPWR c$2876 s$2877 sky130_fd_sc_hd__fa_1
XFILLER_16_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_47_0 pp_row47_0 pp_row47_1 pp_row47_2 VGND VGND VPWR VPWR c$302 s$303
+ sky130_fd_sc_hd__fa_1
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_590 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_83_3 s$1727 s$1729 s$1731 VGND VGND VPWR VPWR c$2508 s$2509 sky130_fd_sc_hd__fa_1
XFILLER_124_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_76_2 c$1636 s$1639 s$1641 VGND VGND VPWR VPWR c$2450 s$2451 sky130_fd_sc_hd__fa_1
XFILLER_151_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1500 net1501 VGND VGND VPWR VPWR net1500 sky130_fd_sc_hd__clkbuf_4
Xfanout1511 net1514 VGND VGND VPWR VPWR net1511 sky130_fd_sc_hd__buf_4
XFILLER_78_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_69_1 c$1546 c$1548 c$1550 VGND VGND VPWR VPWR c$2392 s$2393 sky130_fd_sc_hd__fa_1
Xfanout1522 net125 VGND VGND VPWR VPWR net1522 sky130_fd_sc_hd__buf_6
Xfanout1533 net1534 VGND VGND VPWR VPWR net1533 sky130_fd_sc_hd__buf_2
Xdadda_fa_6_46_0 c$3576 c$3578 s$3581 VGND VGND VPWR VPWR c$3988 s$3989 sky130_fd_sc_hd__fa_1
Xfanout1544 net1546 VGND VGND VPWR VPWR net1544 sky130_fd_sc_hd__buf_4
Xfanout1555 net1559 VGND VGND VPWR VPWR net1555 sky130_fd_sc_hd__buf_6
XU$$4003 net1215 net452 net1205 net725 VGND VGND VPWR VPWR t$6451 sky130_fd_sc_hd__a22o_1
XU$$4014 t$6456 net1282 VGND VGND VPWR VPWR booth_b58_m17 sky130_fd_sc_hd__xor2_1
Xfanout1566 net1567 VGND VGND VPWR VPWR net1566 sky130_fd_sc_hd__buf_6
Xfanout1577 net12 VGND VGND VPWR VPWR net1577 sky130_fd_sc_hd__buf_6
XU$$4025 net1103 net454 net1094 net727 VGND VGND VPWR VPWR t$6462 sky130_fd_sc_hd__a22o_1
Xfanout590 net592 VGND VGND VPWR VPWR net590 sky130_fd_sc_hd__clkbuf_4
XU$$4036 t$6467 net1286 VGND VGND VPWR VPWR booth_b58_m28 sky130_fd_sc_hd__xor2_1
Xfanout1588 net1594 VGND VGND VPWR VPWR net1588 sky130_fd_sc_hd__buf_4
XU$$3302 net938 net497 net1678 net770 VGND VGND VPWR VPWR t$6093 sky130_fd_sc_hd__a22o_1
Xfanout1599 net1603 VGND VGND VPWR VPWR net1599 sky130_fd_sc_hd__clkbuf_8
XU$$4047 net996 net455 net988 net728 VGND VGND VPWR VPWR t$6473 sky130_fd_sc_hd__a22o_1
XU$$4058 t$6478 net1289 VGND VGND VPWR VPWR booth_b58_m39 sky130_fd_sc_hd__xor2_1
XFILLER_65_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3313 t$6098 net1346 VGND VGND VPWR VPWR booth_b48_m9 sky130_fd_sc_hd__xor2_1
XU$$4069 net1728 net457 net1718 net730 VGND VGND VPWR VPWR t$6484 sky130_fd_sc_hd__a22o_1
XU$$3324 net1177 net493 net1168 net766 VGND VGND VPWR VPWR t$6104 sky130_fd_sc_hd__a22o_1
XU$$3335 t$6109 net1343 VGND VGND VPWR VPWR booth_b48_m20 sky130_fd_sc_hd__xor2_1
XFILLER_111_1143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2601 t$5733 net1411 VGND VGND VPWR VPWR booth_b36_m64 sky130_fd_sc_hd__xor2_1
XFILLER_20_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3346 net1073 net493 net1065 net766 VGND VGND VPWR VPWR t$6115 sky130_fd_sc_hd__a22o_1
XU$$2612 t$5740 net1395 VGND VGND VPWR VPWR booth_b38_m1 sky130_fd_sc_hd__xor2_1
XFILLER_94_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_105_2 s$2681 s$2683 s$2685 VGND VGND VPWR VPWR c$3324 s$3325 sky130_fd_sc_hd__fa_1
XFILLER_62_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3357 t$6120 net1340 VGND VGND VPWR VPWR booth_b48_m31 sky130_fd_sc_hd__xor2_1
XFILLER_18_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3368 net966 net495 net959 net768 VGND VGND VPWR VPWR t$6126 sky130_fd_sc_hd__a22o_1
XU$$2623 net1520 net543 net1512 net816 VGND VGND VPWR VPWR t$5746 sky130_fd_sc_hd__a22o_1
XU$$2634 t$5751 net1399 VGND VGND VPWR VPWR booth_b38_m12 sky130_fd_sc_hd__xor2_1
XFILLER_34_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3379 t$6131 net1345 VGND VGND VPWR VPWR booth_b48_m42 sky130_fd_sc_hd__xor2_1
XU$$2645 net1150 net549 net1144 net822 VGND VGND VPWR VPWR t$5757 sky130_fd_sc_hd__a22o_1
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1900 t$5375 net1463 VGND VGND VPWR VPWR booth_b26_m56 sky130_fd_sc_hd__xor2_1
XU$$2656 t$5762 net1395 VGND VGND VPWR VPWR booth_b38_m23 sky130_fd_sc_hd__xor2_1
XU$$1911 net1545 net600 net1537 net873 VGND VGND VPWR VPWR t$5381 sky130_fd_sc_hd__a22o_1
XU$$2667 net1053 net547 net1045 net820 VGND VGND VPWR VPWR t$5768 sky130_fd_sc_hd__a22o_1
XU$$1922 notblock$5385\[2\] net21 net1463 t$5386 notblock$5385\[0\] VGND VGND VPWR
+ VPWR sel_0$5387 sky130_fd_sc_hd__a32o_1
XFILLER_62_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1933 t$5393 net1451 VGND VGND VPWR VPWR booth_b28_m4 sky130_fd_sc_hd__xor2_1
XU$$2678 t$5773 net1397 VGND VGND VPWR VPWR booth_b38_m34 sky130_fd_sc_hd__xor2_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1944 net1494 net584 net1219 net857 VGND VGND VPWR VPWR t$5399 sky130_fd_sc_hd__a22o_1
XU$$2689 net943 net546 net927 net819 VGND VGND VPWR VPWR t$5779 sky130_fd_sc_hd__a22o_1
XU$$1955 t$5404 net1448 VGND VGND VPWR VPWR booth_b28_m15 sky130_fd_sc_hd__xor2_1
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1966 net1116 net584 net1107 net857 VGND VGND VPWR VPWR t$5410 sky130_fd_sc_hd__a22o_1
XU$$1977 t$5415 net1452 VGND VGND VPWR VPWR booth_b28_m26 sky130_fd_sc_hd__xor2_1
X_1951_ clknet_leaf_66_clk booth_b6_m48 VGND VGND VPWR VPWR pp_row54_3 sky130_fd_sc_hd__dfxtp_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1988 net1016 net586 net999 net859 VGND VGND VPWR VPWR t$5421 sky130_fd_sc_hd__a22o_1
XFILLER_109_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1999 t$5426 net1452 VGND VGND VPWR VPWR booth_b28_m37 sky130_fd_sc_hd__xor2_1
X_0902_ clknet_leaf_102_clk booth_b32_m64 VGND VGND VPWR VPWR pp_row96_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_147_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1882_ clknet_leaf_232_clk net203 VGND VGND VPWR VPWR pp_row51_26 sky130_fd_sc_hd__dfxtp_1
XFILLER_147_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_119_0 s$3875 c$4132 s$4135 VGND VGND VPWR VPWR c$4390 s$4391 sky130_fd_sc_hd__fa_1
XFILLER_31_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0833_ clknet_leaf_180_clk notsign$6644 VGND VGND VPWR VPWR pp_row127_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0764_ clknet_leaf_152_clk booth_b60_m29 VGND VGND VPWR VPWR pp_row89_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_116_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2503_ clknet_leaf_179_clk booth_b62_m63 VGND VGND VPWR VPWR pp_row125_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_116_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0695_ clknet_leaf_174_clk booth_b24_m63 VGND VGND VPWR VPWR pp_row87_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_115_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2434_ clknet_leaf_74_clk booth_b48_m19 VGND VGND VPWR VPWR pp_row67_24 sky130_fd_sc_hd__dfxtp_1
XFILLER_9_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_71_1 c$712 c$714 c$716 VGND VGND VPWR VPWR c$1580 s$1581 sky130_fd_sc_hd__fa_1
XFILLER_69_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2365_ clknet_leaf_74_clk booth_b58_m7 VGND VGND VPWR VPWR pp_row65_29 sky130_fd_sc_hd__dfxtp_1
XFILLER_97_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_64_0 s$95 c$582 c$584 VGND VGND VPWR VPWR c$1494 s$1495 sky130_fd_sc_hd__fa_1
XFILLER_111_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$607 final_adder.p_new$610 final_adder.g_new$619 final_adder.g_new$611
+ VGND VGND VPWR VPWR final_adder.g_new$735 sky130_fd_sc_hd__a21o_1
X_1316_ clknet_leaf_122_clk booth_b64_m39 VGND VGND VPWR VPWR pp_row103_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2296_ clknet_leaf_231_clk net216 VGND VGND VPWR VPWR pp_row63_32 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$629 final_adder.p_new$636 final_adder.g_new$653 final_adder.g_new$637
+ VGND VGND VPWR VPWR final_adder.g_new$757 sky130_fd_sc_hd__a21o_1
X_1247_ clknet_leaf_10_clk booth_b2_m23 VGND VGND VPWR VPWR pp_row25_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_25_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$40 net1157 net443 net1147 net685 VGND VGND VPWR VPWR t$4427 sky130_fd_sc_hd__a22o_1
XU$$51 t$4432 net1575 VGND VGND VPWR VPWR booth_b0_m22 sky130_fd_sc_hd__xor2_1
XU$$62 net1055 net442 net1047 net684 VGND VGND VPWR VPWR t$4438 sky130_fd_sc_hd__a22o_1
XFILLER_53_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1178_ clknet_leaf_50_clk booth_b10_m10 VGND VGND VPWR VPWR pp_row20_5 sky130_fd_sc_hd__dfxtp_1
XU$$73 t$4443 net1574 VGND VGND VPWR VPWR booth_b0_m33 sky130_fd_sc_hd__xor2_1
XU$$84 net952 net448 net947 net690 VGND VGND VPWR VPWR t$4449 sky130_fd_sc_hd__a22o_1
XU$$3880 net1141 net460 net1136 net733 VGND VGND VPWR VPWR t$6388 sky130_fd_sc_hd__a22o_1
XU$$95 t$4454 net1572 VGND VGND VPWR VPWR booth_b0_m44 sky130_fd_sc_hd__xor2_1
XU$$3891 t$6393 net1292 VGND VGND VPWR VPWR booth_b56_m24 sky130_fd_sc_hd__xor2_1
XFILLER_80_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_20 sel_0$6227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_31 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1025 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_42 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_53 net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_64 net414 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_75 net458 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_86 net518 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdadda_fa_4_93_2 s$2585 s$2587 s$2589 VGND VGND VPWR VPWR c$3252 s$3253 sky130_fd_sc_hd__fa_1
XANTENNA_97 net534 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_86_1 c$2522 c$2524 s$2527 VGND VGND VPWR VPWR c$3208 s$3209 sky130_fd_sc_hd__fa_1
XFILLER_137_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_63_0 s$3651 c$4020 s$4023 VGND VGND VPWR VPWR c$4278 s$4279 sky130_fd_sc_hd__fa_2
XFILLER_106_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_79_0 s$1685 c$2462 c$2464 VGND VGND VPWR VPWR c$3164 s$3165 sky130_fd_sc_hd__fa_1
XFILLER_97_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1207 t$5021 net1014 VGND VGND VPWR VPWR booth_b16_m52 sky130_fd_sc_hd__xor2_1
XU$$1218 net1595 net649 net1586 net922 VGND VGND VPWR VPWR t$5027 sky130_fd_sc_hd__a22o_1
XFILLER_43_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1229 t$5032 net1013 VGND VGND VPWR VPWR booth_b16_m63 sky130_fd_sc_hd__xor2_1
XFILLER_31_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1001 final_adder.$signal$1130 final_adder.g_new$955 VGND VGND VPWR
+ VPWR net319 sky130_fd_sc_hd__xor2_2
XFILLER_178_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1012 final_adder.$signal$105 final_adder.g_new$1064 VGND VGND VPWR
+ VPWR net331 sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$1023 final_adder.$signal$1152 final_adder.g_new$933 VGND VGND VPWR
+ VPWR net343 sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$1034 final_adder.$signal$1163 final_adder.g_new$1053 VGND VGND VPWR
+ VPWR net355 sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$1045 final_adder.$signal$1174 final_adder.g_new$1007 VGND VGND VPWR
+ VPWR net367 sky130_fd_sc_hd__xor2_2
XFILLER_109_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$1056 final_adder.$signal$1185 final_adder.g_new$1042 VGND VGND VPWR
+ VPWR net379 sky130_fd_sc_hd__xor2_1
XFILLER_171_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$1067 final_adder.$signal$1196 final_adder.g_new$985 VGND VGND VPWR
+ VPWR net264 sky130_fd_sc_hd__xor2_2
Xclkbuf_5_31__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_5_31__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xfinal_adder.U$$1078 final_adder.$signal$1207 final_adder.g_new$1031 VGND VGND VPWR
+ VPWR net276 sky130_fd_sc_hd__xor2_2
Xdadda_fa_3_81_0 s$921 c$1686 c$1688 VGND VGND VPWR VPWR c$2486 s$2487 sky130_fd_sc_hd__fa_1
XFILLER_125_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0480_ clknet_leaf_205_clk booth_b28_m51 VGND VGND VPWR VPWR pp_row79_7 sky130_fd_sc_hd__dfxtp_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1330 net1332 VGND VGND VPWR VPWR net1330 sky130_fd_sc_hd__buf_6
Xfanout1341 net1347 VGND VGND VPWR VPWR net1341 sky130_fd_sc_hd__buf_6
XFILLER_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2150_ clknet_leaf_215_clk booth_b0_m60 VGND VGND VPWR VPWR pp_row60_0 sky130_fd_sc_hd__dfxtp_1
Xfanout1352 net42 VGND VGND VPWR VPWR net1352 sky130_fd_sc_hd__buf_4
XFILLER_79_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1363 net1366 VGND VGND VPWR VPWR net1363 sky130_fd_sc_hd__buf_4
XFILLER_78_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1374 net1375 VGND VGND VPWR VPWR net1374 sky130_fd_sc_hd__buf_4
X_1101_ clknet_leaf_248_clk net161 VGND VGND VPWR VPWR pp_row13_7 sky130_fd_sc_hd__dfxtp_2
Xfanout1385 net1386 VGND VGND VPWR VPWR net1385 sky130_fd_sc_hd__buf_6
Xfanout1396 net1398 VGND VGND VPWR VPWR net1396 sky130_fd_sc_hd__buf_8
XFILLER_94_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3110 net1723 net513 net1714 net786 VGND VGND VPWR VPWR t$5994 sky130_fd_sc_hd__a22o_1
X_2081_ clknet_leaf_86_clk booth_b2_m56 VGND VGND VPWR VPWR pp_row58_1 sky130_fd_sc_hd__dfxtp_1
XU$$3121 t$5999 net1364 VGND VGND VPWR VPWR booth_b44_m50 sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_43_5 s$257 s$259 s$261 VGND VGND VPWR VPWR c$1252 s$1253 sky130_fd_sc_hd__fa_1
XFILLER_93_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_110_0 pp_row110_11 c$2710 c$2712 VGND VGND VPWR VPWR c$3350 s$3351 sky130_fd_sc_hd__fa_1
XU$$3132 net1618 net515 net1609 net788 VGND VGND VPWR VPWR t$6005 sky130_fd_sc_hd__a22o_1
XFILLER_53_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1032_ clknet_leaf_60_clk booth_b4_m0 VGND VGND VPWR VPWR pp_row4_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_53_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3143 t$6010 net1365 VGND VGND VPWR VPWR booth_b44_m61 sky130_fd_sc_hd__xor2_1
XU$$3154 net1350 notblock$6015\[1\] VGND VGND VPWR VPWR t$6016 sky130_fd_sc_hd__and2_1
XU$$3165 net938 net505 net1677 net778 VGND VGND VPWR VPWR t$6023 sky130_fd_sc_hd__a22o_1
XU$$2420 t$5641 net1425 VGND VGND VPWR VPWR booth_b34_m42 sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_36_4 pp_row36_17 pp_row36_18 pp_row36_19 VGND VGND VPWR VPWR c$1166 s$1167
+ sky130_fd_sc_hd__fa_1
XU$$2431 net1696 net566 net1688 net839 VGND VGND VPWR VPWR t$5647 sky130_fd_sc_hd__a22o_1
XFILLER_19_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3176 t$6028 net1353 VGND VGND VPWR VPWR booth_b46_m9 sky130_fd_sc_hd__xor2_1
XU$$2442 t$5652 net1426 VGND VGND VPWR VPWR booth_b34_m53 sky130_fd_sc_hd__xor2_1
XU$$3187 net1177 net501 net1168 net774 VGND VGND VPWR VPWR t$6034 sky130_fd_sc_hd__a22o_1
XFILLER_185_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2453 net1590 net567 net1582 net840 VGND VGND VPWR VPWR t$5658 sky130_fd_sc_hd__a22o_1
XU$$3198 t$6039 net1353 VGND VGND VPWR VPWR booth_b46_m20 sky130_fd_sc_hd__xor2_1
XU$$2464 t$5663 net1428 VGND VGND VPWR VPWR booth_b34_m64 sky130_fd_sc_hd__xor2_1
XFILLER_34_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2475 t$5670 net1403 VGND VGND VPWR VPWR booth_b36_m1 sky130_fd_sc_hd__xor2_1
XU$$1730 net944 net606 net928 net879 VGND VGND VPWR VPWR t$5289 sky130_fd_sc_hd__a22o_1
XFILLER_34_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2486 net1520 net551 net1512 net824 VGND VGND VPWR VPWR t$5676 sky130_fd_sc_hd__a22o_1
XU$$1741 t$5294 net1474 VGND VGND VPWR VPWR booth_b24_m45 sky130_fd_sc_hd__xor2_1
XU$$1752 net1654 net607 net1646 net880 VGND VGND VPWR VPWR t$5300 sky130_fd_sc_hd__a22o_1
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2497 t$5681 net1403 VGND VGND VPWR VPWR booth_b36_m12 sky130_fd_sc_hd__xor2_1
XFILLER_107_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1763 t$5305 net1472 VGND VGND VPWR VPWR booth_b24_m56 sky130_fd_sc_hd__xor2_1
XFILLER_188_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1774 net1544 net608 net1536 net881 VGND VGND VPWR VPWR t$5311 sky130_fd_sc_hd__a22o_1
XU$$1785 notblock$5315\[2\] net19 net1472 t$5316 notblock$5315\[0\] VGND VGND VPWR
+ VPWR sel_0$5317 sky130_fd_sc_hd__a32o_1
XU$$1796 t$5323 net1457 VGND VGND VPWR VPWR booth_b26_m4 sky130_fd_sc_hd__xor2_1
X_1934_ clknet_leaf_69_clk booth_b34_m19 VGND VGND VPWR VPWR pp_row53_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_30_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1865_ clknet_leaf_66_clk booth_b20_m31 VGND VGND VPWR VPWR pp_row51_10 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_96_0 c$3260 c$3262 c$3264 VGND VGND VPWR VPWR c$3780 s$3781 sky130_fd_sc_hd__fa_1
Xinput40 a[45] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
XFILLER_174_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0816_ clknet_leaf_93_clk booth_b30_m62 VGND VGND VPWR VPWR pp_row92_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput51 a[55] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_1
Xinput62 a[7] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_2
X_1796_ clknet_leaf_37_clk booth_b4_m45 VGND VGND VPWR VPWR pp_row49_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_156_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput73 b[17] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_2
XFILLER_128_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput84 b[27] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_4
XFILLER_157_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput95 b[37] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__buf_2
XFILLER_190_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0747_ clknet_leaf_143_clk booth_b28_m61 VGND VGND VPWR VPWR pp_row89_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_171_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0678_ clknet_leaf_179_clk booth_b38_m48 VGND VGND VPWR VPWR pp_row86_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_130_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2417_ clknet_leaf_92_clk booth_b16_m51 VGND VGND VPWR VPWR pp_row67_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_112_950 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$404 final_adder.p_new$410 final_adder.p_new$406 VGND VGND VPWR VPWR
+ final_adder.p_new$532 sky130_fd_sc_hd__and2_1
X_2348_ clknet_leaf_127_clk booth_b50_m61 VGND VGND VPWR VPWR pp_row111_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_123_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$415 final_adder.p_new$416 final_adder.g_new$421 final_adder.g_new$417
+ VGND VGND VPWR VPWR final_adder.g_new$543 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$426 final_adder.p_new$432 final_adder.p_new$428 VGND VGND VPWR VPWR
+ final_adder.p_new$554 sky130_fd_sc_hd__and2_1
XTAP_3708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$437 final_adder.p_new$438 final_adder.g_new$443 final_adder.g_new$439
+ VGND VGND VPWR VPWR final_adder.g_new$565 sky130_fd_sc_hd__a21o_1
XTAP_3719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$448 final_adder.p_new$454 final_adder.p_new$450 VGND VGND VPWR VPWR
+ final_adder.p_new$576 sky130_fd_sc_hd__and2_1
X_2279_ clknet_leaf_212_clk booth_b36_m27 VGND VGND VPWR VPWR pp_row63_18 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$459 final_adder.p_new$460 final_adder.g_new$465 final_adder.g_new$461
+ VGND VGND VPWR VPWR final_adder.g_new$587 sky130_fd_sc_hd__a21o_1
XU$$309 t$4563 net1274 VGND VGND VPWR VPWR booth_b4_m14 sky130_fd_sc_hd__xor2_1
XFILLER_38_1128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_105_1 pp_row105_9 pp_row105_10 pp_row105_11 VGND VGND VPWR VPWR c$2680
+ s$2681 sky130_fd_sc_hd__fa_1
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_126_0 pp_row126_2 pp_row126_3 c$3896 VGND VGND VPWR VPWR c$4148 s$4149
+ sky130_fd_sc_hd__fa_1
XFILLER_0_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_0_69_4 pp_row69_12 pp_row69_13 pp_row69_14 VGND VGND VPWR VPWR c$152 s$153
+ sky130_fd_sc_hd__fa_1
XFILLER_48_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_46_3 s$1283 s$1285 s$1287 VGND VGND VPWR VPWR c$2212 s$2213 sky130_fd_sc_hd__fa_1
XFILLER_180_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$960 final_adder.$signal$1092 final_adder.g_new$383 final_adder.$signal$6
+ VGND VGND VPWR VPWR final_adder.g_new$1088 sky130_fd_sc_hd__a21o_1
XFILLER_17_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$971 final_adder.$signal$1100 final_adder.g_new$753 VGND VGND VPWR
+ VPWR net268 sky130_fd_sc_hd__xor2_2
XU$$810 t$4818 net1419 VGND VGND VPWR VPWR booth_b10_m59 sky130_fd_sc_hd__xor2_1
XU$$821 net1417 VGND VGND VPWR VPWR notsign$4824 sky130_fd_sc_hd__inv_1
XFILLER_29_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_39_2 c$1192 s$1195 s$1197 VGND VGND VPWR VPWR c$2154 s$2155 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$982 final_adder.$signal$1111 final_adder.g_new$1079 VGND VGND VPWR
+ VPWR net298 sky130_fd_sc_hd__xor2_2
XU$$832 net1123 net396 net1032 net662 VGND VGND VPWR VPWR t$4831 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$993 final_adder.$signal$1122 final_adder.g_new$851 VGND VGND VPWR
+ VPWR net310 sky130_fd_sc_hd__xor2_2
XU$$843 t$4836 net1312 VGND VGND VPWR VPWR booth_b12_m7 sky130_fd_sc_hd__xor2_1
XFILLER_44_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$854 net1202 net394 net1193 net660 VGND VGND VPWR VPWR t$4842 sky130_fd_sc_hd__a22o_1
XU$$865 t$4847 net1310 VGND VGND VPWR VPWR booth_b12_m18 sky130_fd_sc_hd__xor2_1
XU$$1004 t$4918 net1185 VGND VGND VPWR VPWR booth_b14_m19 sky130_fd_sc_hd__xor2_1
XFILLER_16_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1015 net1081 net387 net1072 net653 VGND VGND VPWR VPWR t$4924 sky130_fd_sc_hd__a22o_1
XU$$876 net1091 net397 net1083 net663 VGND VGND VPWR VPWR t$4853 sky130_fd_sc_hd__a22o_1
XFILLER_32_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1026 t$4929 net1184 VGND VGND VPWR VPWR booth_b14_m30 sky130_fd_sc_hd__xor2_1
XU$$887 t$4858 net1311 VGND VGND VPWR VPWR booth_b12_m29 sky130_fd_sc_hd__xor2_1
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$898 net982 net393 net973 net659 VGND VGND VPWR VPWR t$4864 sky130_fd_sc_hd__a22o_1
XU$$1037 net977 net388 net969 net654 VGND VGND VPWR VPWR t$4935 sky130_fd_sc_hd__a22o_1
XFILLER_32_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1048 t$4940 net1186 VGND VGND VPWR VPWR booth_b14_m41 sky130_fd_sc_hd__xor2_1
XU$$1059 net1703 net390 net1695 net656 VGND VGND VPWR VPWR t$4946 sky130_fd_sc_hd__a22o_1
XFILLER_43_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1650_ clknet_leaf_124_clk booth_b42_m64 VGND VGND VPWR VPWR pp_row106_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_171_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0601_ clknet_leaf_188_clk booth_b42_m41 VGND VGND VPWR VPWR pp_row83_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_160_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1581_ clknet_leaf_243_clk booth_b10_m31 VGND VGND VPWR VPWR pp_row41_5 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_246_clk clknet_5_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_246_clk
+ sky130_fd_sc_hd__clkbuf_16
X_0532_ clknet_leaf_159_clk booth_b18_m63 VGND VGND VPWR VPWR pp_row81_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_99_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0463_ clknet_leaf_206_clk booth_b52_m26 VGND VGND VPWR VPWR pp_row78_20 sky130_fd_sc_hd__dfxtp_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2202_ clknet_leaf_88_clk booth_b28_m33 VGND VGND VPWR VPWR pp_row61_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0394_ clknet_leaf_191_clk booth_b36_m40 VGND VGND VPWR VPWR pp_row76_13 sky130_fd_sc_hd__dfxtp_1
Xfanout1160 net72 VGND VGND VPWR VPWR net1160 sky130_fd_sc_hd__buf_2
Xfanout1171 net1172 VGND VGND VPWR VPWR net1171 sky130_fd_sc_hd__clkbuf_4
XFILLER_39_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1182 net70 VGND VGND VPWR VPWR net1182 sky130_fd_sc_hd__clkbuf_8
X_2133_ clknet_leaf_32_clk booth_b32_m27 VGND VGND VPWR VPWR pp_row59_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_120_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1193 net1195 VGND VGND VPWR VPWR net1193 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_41_2 pp_row41_17 pp_row41_18 pp_row41_19 VGND VGND VPWR VPWR c$1222 s$1223
+ sky130_fd_sc_hd__fa_1
XFILLER_54_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2064_ clknet_leaf_35_clk booth_b30_m27 VGND VGND VPWR VPWR pp_row57_15 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_34_1 pp_row34_5 pp_row34_6 pp_row34_7 VGND VGND VPWR VPWR c$1136 s$1137
+ sky130_fd_sc_hd__fa_1
X_1015_ clknet_leaf_120_clk booth_b38_m64 VGND VGND VPWR VPWR pp_row102_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_62_550 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2250 net1075 net572 net1067 net845 VGND VGND VPWR VPWR t$5555 sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_11_0 pp_row11_5 pp_row11_6 c$2754 VGND VGND VPWR VPWR c$3440 s$3441 sky130_fd_sc_hd__fa_1
Xdadda_fa_2_27_0 pp_row27_0 pp_row27_1 pp_row27_2 VGND VGND VPWR VPWR c$1068 s$1069
+ sky130_fd_sc_hd__fa_1
XU$$2261 t$5560 net1431 VGND VGND VPWR VPWR booth_b32_m31 sky130_fd_sc_hd__xor2_1
XFILLER_35_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2272 net970 net575 net962 net848 VGND VGND VPWR VPWR t$5566 sky130_fd_sc_hd__a22o_1
XU$$2283 t$5571 net1438 VGND VGND VPWR VPWR booth_b32_m42 sky130_fd_sc_hd__xor2_1
XU$$2294 net1696 net573 net1688 net846 VGND VGND VPWR VPWR t$5577 sky130_fd_sc_hd__a22o_1
XU$$1560 t$5202 net1476 VGND VGND VPWR VPWR booth_b22_m23 sky130_fd_sc_hd__xor2_1
XU$$1571 net1049 net615 net1041 net888 VGND VGND VPWR VPWR t$5208 sky130_fd_sc_hd__a22o_1
XFILLER_179_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1582 t$5213 net1478 VGND VGND VPWR VPWR booth_b22_m34 sky130_fd_sc_hd__xor2_1
XFILLER_148_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1593 net940 net612 net924 net885 VGND VGND VPWR VPWR t$5219 sky130_fd_sc_hd__a22o_1
XFILLER_31_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1917_ clknet_leaf_68_clk booth_b2_m51 VGND VGND VPWR VPWR pp_row53_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_191_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1848_ clknet_leaf_73_clk booth_b46_m4 VGND VGND VPWR VPWR pp_row50_23 sky130_fd_sc_hd__dfxtp_1
XFILLER_129_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1779_ clknet_leaf_220_clk booth_b28_m20 VGND VGND VPWR VPWR pp_row48_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_162_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_237_clk clknet_5_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_237_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_190_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_86_4 pp_row86_12 pp_row86_13 pp_row86_14 VGND VGND VPWR VPWR c$986 s$987
+ sky130_fd_sc_hd__fa_1
XFILLER_143_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_79_3 pp_row79_9 pp_row79_10 pp_row79_11 VGND VGND VPWR VPWR c$876 s$877
+ sky130_fd_sc_hd__fa_1
XFILLER_98_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_56_2 s$2289 s$2291 s$2293 VGND VGND VPWR VPWR c$3030 s$3031 sky130_fd_sc_hd__fa_1
XTAP_4206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$201 final_adder.$signal$113 final_adder.$signal$110 final_adder.$signal$112
+ VGND VGND VPWR VPWR final_adder.g_new$329 sky130_fd_sc_hd__a21o_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$212 final_adder.$signal$1132 final_adder.$signal$1133 VGND VGND VPWR
+ VPWR final_adder.p_new$340 sky130_fd_sc_hd__and2_1
XTAP_4239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_49_1 c$2226 c$2228 s$2231 VGND VGND VPWR VPWR c$2986 s$2987 sky130_fd_sc_hd__fa_1
XFILLER_58_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$223 final_adder.$signal$1123 final_adder.$signal$66 final_adder.$signal$68
+ VGND VGND VPWR VPWR final_adder.g_new$351 sky130_fd_sc_hd__a21o_1
XTAP_3505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$234 final_adder.$signal$1110 final_adder.$signal$1111 VGND VGND VPWR
+ VPWR final_adder.p_new$362 sky130_fd_sc_hd__and2_1
XTAP_3516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$245 final_adder.$signal$1101 final_adder.$signal$22 final_adder.$signal$24
+ VGND VGND VPWR VPWR final_adder.g_new$373 sky130_fd_sc_hd__a21o_1
XTAP_3527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_26_0 s$3503 c$3946 s$3949 VGND VGND VPWR VPWR c$4204 s$4205 sky130_fd_sc_hd__fa_1
XFILLER_45_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$106 net1679 net445 net1654 net687 VGND VGND VPWR VPWR t$4460 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$267 final_adder.p_new$266 final_adder.g_new$269 final_adder.g_new$267
+ VGND VGND VPWR VPWR final_adder.g_new$395 sky130_fd_sc_hd__a21o_1
XU$$117 t$4465 net1576 VGND VGND VPWR VPWR booth_b0_m55 sky130_fd_sc_hd__xor2_1
XTAP_3549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$278 final_adder.p_new$280 final_adder.p_new$278 VGND VGND VPWR VPWR
+ final_adder.p_new$406 sky130_fd_sc_hd__and2_1
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$128 net1551 net444 net1543 net686 VGND VGND VPWR VPWR t$4471 sky130_fd_sc_hd__a22o_1
XFILLER_73_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$289 final_adder.p_new$288 final_adder.g_new$291 final_adder.g_new$289
+ VGND VGND VPWR VPWR final_adder.g_new$417 sky130_fd_sc_hd__a21o_1
XU$$139 net1387 VGND VGND VPWR VPWR notblock$4475\[2\] sky130_fd_sc_hd__inv_1
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_228_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_228_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput230 c[76] VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_3_51_1 c$1330 c$1332 c$1334 VGND VGND VPWR VPWR c$2248 s$2249 sky130_fd_sc_hd__fa_2
Xinput241 c[86] VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput252 c[96] VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_0_67_1 pp_row67_3 pp_row67_4 pp_row67_5 VGND VGND VPWR VPWR c$122 s$123
+ sky130_fd_sc_hd__fa_1
XFILLER_48_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_44_0 s$275 c$1242 c$1244 VGND VGND VPWR VPWR c$2190 s$2191 sky130_fd_sc_hd__fa_1
XFILLER_91_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$790 final_adder.p_new$838 final_adder.p_new$806 VGND VGND VPWR VPWR
+ final_adder.p_new$918 sky130_fd_sc_hd__and2_1
XU$$640 net1744 net416 net1736 net682 VGND VGND VPWR VPWR t$4732 sky130_fd_sc_hd__a22o_1
XU$$651 t$4737 net1242 VGND VGND VPWR VPWR booth_b8_m48 sky130_fd_sc_hd__xor2_1
XU$$662 net1629 net411 net1620 net677 VGND VGND VPWR VPWR t$4743 sky130_fd_sc_hd__a22o_1
XFILLER_95_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$673 t$4748 net1243 VGND VGND VPWR VPWR booth_b8_m59 sky130_fd_sc_hd__xor2_1
XU$$684 net1237 VGND VGND VPWR VPWR notsign$4754 sky130_fd_sc_hd__inv_1
XU$$695 net1127 net404 net1035 net670 VGND VGND VPWR VPWR t$4761 sky130_fd_sc_hd__a22o_1
XFILLER_108_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_101_0 s$3803 c$4096 s$4099 VGND VGND VPWR VPWR c$4354 s$4355 sky130_fd_sc_hd__fa_1
XFILLER_172_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1702_ clknet_leaf_23_clk booth_b40_m5 VGND VGND VPWR VPWR pp_row45_20 sky130_fd_sc_hd__dfxtp_1
XFILLER_118_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1633_ clknet_leaf_242_clk booth_b10_m33 VGND VGND VPWR VPWR pp_row43_5 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_96_3 pp_row96_11 pp_row96_12 pp_row96_13 VGND VGND VPWR VPWR c$1884 s$1885
+ sky130_fd_sc_hd__fa_1
XFILLER_172_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_219_clk clknet_5_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_219_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_67_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1564_ clknet_leaf_8_clk booth_b24_m16 VGND VGND VPWR VPWR pp_row40_12 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_89_2 pp_row89_18 pp_row89_19 pp_row89_20 VGND VGND VPWR VPWR c$1798 s$1799
+ sky130_fd_sc_hd__fa_1
XFILLER_99_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_66_1 s$3087 s$3089 s$3091 VGND VGND VPWR VPWR c$3662 s$3663 sky130_fd_sc_hd__fa_1
Xfanout408 sel_0$4757 VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__buf_6
X_0515_ clknet_leaf_156_clk booth_b38_m42 VGND VGND VPWR VPWR pp_row80_12 sky130_fd_sc_hd__dfxtp_1
Xfanout419 net421 VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__buf_4
X_1495_ clknet_leaf_45_clk booth_b26_m11 VGND VGND VPWR VPWR pp_row37_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_115_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_59_0 c$3038 c$3040 c$3042 VGND VGND VPWR VPWR c$3632 s$3633 sky130_fd_sc_hd__fa_1
XFILLER_141_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0446_ clknet_leaf_207_clk booth_b20_m58 VGND VGND VPWR VPWR pp_row78_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_86_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_58_8 s$25 s$27 s$29 VGND VGND VPWR VPWR c$508 s$509 sky130_fd_sc_hd__fa_1
X_0377_ clknet_leaf_126_clk booth_b58_m56 VGND VGND VPWR VPWR pp_row114_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_82_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2116_ clknet_leaf_137_clk booth_b52_m57 VGND VGND VPWR VPWR pp_row109_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_55_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2047_ clknet_leaf_82_clk booth_b2_m55 VGND VGND VPWR VPWR pp_row57_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_105_0 pp_row105_0 pp_row105_1 pp_row105_2 VGND VGND VPWR VPWR c$1962 s$1963
+ sky130_fd_sc_hd__fa_1
XU$$2080 t$5468 net1439 VGND VGND VPWR VPWR booth_b30_m9 sky130_fd_sc_hd__xor2_1
XFILLER_23_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2091 net1176 net577 net1167 net850 VGND VGND VPWR VPWR t$5474 sky130_fd_sc_hd__a22o_1
XFILLER_167_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1390 net1519 net627 net1511 net900 VGND VGND VPWR VPWR t$5116 sky130_fd_sc_hd__a22o_1
XFILLER_10_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_91_2 pp_row91_6 pp_row91_7 pp_row91_8 VGND VGND VPWR VPWR c$1030 s$1031
+ sky130_fd_sc_hd__fa_1
XFILLER_191_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_84_1 pp_row84_3 pp_row84_4 pp_row84_5 VGND VGND VPWR VPWR c$954 s$955
+ sky130_fd_sc_hd__fa_1
XFILLER_145_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_61_0 s$1469 c$2318 c$2320 VGND VGND VPWR VPWR c$3056 s$3057 sky130_fd_sc_hd__fa_1
XFILLER_131_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout920 sel_1$4968 VGND VGND VPWR VPWR net920 sky130_fd_sc_hd__buf_4
Xfanout931 net99 VGND VGND VPWR VPWR net931 sky130_fd_sc_hd__buf_12
Xdadda_fa_1_77_0 pp_row77_3 pp_row77_4 pp_row77_5 VGND VGND VPWR VPWR c$834 s$835
+ sky130_fd_sc_hd__fa_1
Xfanout942 net947 VGND VGND VPWR VPWR net942 sky130_fd_sc_hd__clkbuf_8
Xfanout953 net954 VGND VGND VPWR VPWR net953 sky130_fd_sc_hd__buf_6
XTAP_4003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout964 net965 VGND VGND VPWR VPWR net964 sky130_fd_sc_hd__buf_4
XFILLER_58_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_ha_2_104_2 pp_row104_6 pp_row104_7 VGND VGND VPWR VPWR c$1960 s$1961 sky130_fd_sc_hd__ha_1
Xfanout975 net981 VGND VGND VPWR VPWR net975 sky130_fd_sc_hd__buf_4
XTAP_4025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout986 net92 VGND VGND VPWR VPWR net986 sky130_fd_sc_hd__buf_6
XTAP_4036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout997 net91 VGND VGND VPWR VPWR net997 sky130_fd_sc_hd__clkbuf_8
XTAP_4047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3709 net1129 net472 net1037 net745 VGND VGND VPWR VPWR t$6301 sky130_fd_sc_hd__a22o_1
XTAP_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_302 net417 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_313 net564 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_324 net658 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_335 net715 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_346 net856 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_357 net958 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_368 net1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_379 net1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_99_1 c$1904 c$1906 c$1908 VGND VGND VPWR VPWR c$2632 s$2633 sky130_fd_sc_hd__fa_1
XFILLER_155_967 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_76_0 c$3696 c$3698 s$3701 VGND VGND VPWR VPWR c$4048 s$4049 sky130_fd_sc_hd__fa_1
XFILLER_126_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0300_ clknet_leaf_128_clk booth_b62_m51 VGND VGND VPWR VPWR pp_row113_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_123_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1280_ clknet_leaf_250_clk booth_b2_m25 VGND VGND VPWR VPWR pp_row27_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_68_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0231_ clknet_leaf_151_clk booth_b36_m35 VGND VGND VPWR VPWR pp_row71_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_83_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$470 t$4645 net1245 VGND VGND VPWR VPWR booth_b6_m26 sky130_fd_sc_hd__xor2_1
XU$$481 net1016 net427 net998 net709 VGND VGND VPWR VPWR t$4651 sky130_fd_sc_hd__a22o_1
XU$$492 t$4656 net1244 VGND VGND VPWR VPWR booth_b6_m37 sky130_fd_sc_hd__xor2_1
XFILLER_189_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0995_ clknet_leaf_110_clk booth_b64_m36 VGND VGND VPWR VPWR pp_row100_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_164_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_94_0 pp_row94_5 pp_row94_6 pp_row94_7 VGND VGND VPWR VPWR c$1854 s$1855
+ sky130_fd_sc_hd__fa_1
XFILLER_161_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1616_ clknet_leaf_110_clk booth_b62_m43 VGND VGND VPWR VPWR pp_row105_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_160_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1547_ clknet_leaf_19_clk booth_b36_m3 VGND VGND VPWR VPWR pp_row39_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_8_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_70_7 c$150 c$152 s$155 VGND VGND VPWR VPWR c$722 s$723 sky130_fd_sc_hd__fa_1
XFILLER_113_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1478_ clknet_leaf_38_clk net1406 VGND VGND VPWR VPWR pp_row36_19 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_63_6 c$64 c$66 c$68 VGND VGND VPWR VPWR c$594 s$595 sky130_fd_sc_hd__fa_1
X_0429_ clknet_leaf_207_clk booth_b44_m33 VGND VGND VPWR VPWR pp_row77_16 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_56_5 pp_row56_23 pp_row56_24 pp_row56_25 VGND VGND VPWR VPWR c$466 s$467
+ sky130_fd_sc_hd__fa_1
XFILLER_83_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_49_4 pp_row49_12 pp_row49_13 pp_row49_14 VGND VGND VPWR VPWR c$340 s$341
+ sky130_fd_sc_hd__fa_1
XFILLER_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_19_2 s$1993 s$1995 s$1997 VGND VGND VPWR VPWR c$2808 s$2809 sky130_fd_sc_hd__fa_1
XFILLER_165_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_93_0 s$3771 c$4080 s$4083 VGND VGND VPWR VPWR c$4338 s$4339 sky130_fd_sc_hd__fa_1
XFILLER_149_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1704 net1705 VGND VGND VPWR VPWR net1704 sky130_fd_sc_hd__buf_4
XFILLER_137_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1715 net104 VGND VGND VPWR VPWR net1715 sky130_fd_sc_hd__buf_6
XFILLER_160_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1726 net1727 VGND VGND VPWR VPWR net1726 sky130_fd_sc_hd__buf_4
Xfanout1737 net1738 VGND VGND VPWR VPWR net1737 sky130_fd_sc_hd__buf_4
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout750 net752 VGND VGND VPWR VPWR net750 sky130_fd_sc_hd__buf_4
Xfanout1748 net1752 VGND VGND VPWR VPWR net1748 sky130_fd_sc_hd__clkbuf_4
XFILLER_172_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4207 t$6554 net1271 VGND VGND VPWR VPWR booth_b60_m45 sky130_fd_sc_hd__xor2_1
Xfanout761 net765 VGND VGND VPWR VPWR net761 sky130_fd_sc_hd__buf_4
XFILLER_133_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4218 net1659 net439 net1651 net721 VGND VGND VPWR VPWR t$6560 sky130_fd_sc_hd__a22o_1
Xfanout772 net773 VGND VGND VPWR VPWR net772 sky130_fd_sc_hd__buf_6
Xfanout783 net791 VGND VGND VPWR VPWR net783 sky130_fd_sc_hd__buf_4
XU$$4229 t$6565 net1270 VGND VGND VPWR VPWR booth_b60_m56 sky130_fd_sc_hd__xor2_1
XFILLER_46_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout794 net795 VGND VGND VPWR VPWR net794 sky130_fd_sc_hd__buf_4
XFILLER_93_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3506 t$6196 net1331 VGND VGND VPWR VPWR booth_b50_m37 sky130_fd_sc_hd__xor2_1
XTAP_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3517 net1742 net490 net1734 net763 VGND VGND VPWR VPWR t$6202 sky130_fd_sc_hd__a22o_1
XFILLER_19_848 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3528 t$6207 net1335 VGND VGND VPWR VPWR booth_b50_m48 sky130_fd_sc_hd__xor2_1
XFILLER_18_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3539 net1635 net490 net1626 net763 VGND VGND VPWR VPWR t$6213 sky130_fd_sc_hd__a22o_1
XFILLER_46_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2805 t$5838 net1380 VGND VGND VPWR VPWR booth_b40_m29 sky130_fd_sc_hd__xor2_1
XTAP_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2816 net984 net537 net975 net810 VGND VGND VPWR VPWR t$5844 sky130_fd_sc_hd__a22o_1
XFILLER_73_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_110 net618 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2827 t$5849 net1380 VGND VGND VPWR VPWR booth_b40_m40 sky130_fd_sc_hd__xor2_1
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_121 net656 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2838 net1713 net537 net1704 net810 VGND VGND VPWR VPWR t$5855 sky130_fd_sc_hd__a22o_1
XFILLER_22_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_132 net710 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2849 t$5860 net1383 VGND VGND VPWR VPWR booth_b40_m51 sky130_fd_sc_hd__xor2_1
XFILLER_27_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_143 net769 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_21_2 pp_row21_6 pp_row21_7 pp_row21_8 VGND VGND VPWR VPWR c$2010 s$2011
+ sky130_fd_sc_hd__fa_1
XTAP_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_154 net803 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_165 net885 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_176 net931 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_187 net972 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_198 net1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0780_ clknet_leaf_140_clk booth_b46_m44 VGND VGND VPWR VPWR pp_row90_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_10_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2450_ clknet_leaf_91_clk booth_b12_m56 VGND VGND VPWR VPWR pp_row68_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1401_ clknet_leaf_51_clk booth_b12_m21 VGND VGND VPWR VPWR pp_row33_6 sky130_fd_sc_hd__dfxtp_1
X_2381_ clknet_leaf_83_clk booth_b20_m46 VGND VGND VPWR VPWR pp_row66_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_123_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_73_5 s$773 s$775 s$777 VGND VGND VPWR VPWR c$1612 s$1613 sky130_fd_sc_hd__fa_2
X_1332_ clknet_leaf_244_clk net178 VGND VGND VPWR VPWR pp_row29_15 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_66_4 s$641 s$643 s$645 VGND VGND VPWR VPWR c$1526 s$1527 sky130_fd_sc_hd__fa_2
XFILLER_96_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1263_ clknet_leaf_2_clk booth_b2_m24 VGND VGND VPWR VPWR pp_row26_1 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_59_3 c$508 s$511 s$513 VGND VGND VPWR VPWR c$1440 s$1441 sky130_fd_sc_hd__fa_1
XFILLER_49_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput5 a[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_4
XFILLER_65_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0214_ clknet_leaf_198_clk net224 VGND VGND VPWR VPWR pp_row70_31 sky130_fd_sc_hd__dfxtp_2
X_1194_ clknet_leaf_124_clk booth_b42_m61 VGND VGND VPWR VPWR pp_row103_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_188_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_29_1 s$2865 s$2867 s$2869 VGND VGND VPWR VPWR c$3514 s$3515 sky130_fd_sc_hd__fa_1
XFILLER_80_968 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0978_ clknet_leaf_113_clk booth_b64_m35 VGND VGND VPWR VPWR pp_row99_15 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$3 c$4156 s$4159 VGND VGND VPWR VPWR final_adder.$signal$8 final_adder.$signal$1093
+ sky130_fd_sc_hd__ha_1
XFILLER_173_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_103_1 s$3309 s$3311 s$3313 VGND VGND VPWR VPWR c$3810 s$3811 sky130_fd_sc_hd__fa_1
XFILLER_106_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput320 net320 VGND VGND VPWR VPWR o[41] sky130_fd_sc_hd__buf_2
Xoutput331 net331 VGND VGND VPWR VPWR o[51] sky130_fd_sc_hd__buf_2
XFILLER_126_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput342 net342 VGND VGND VPWR VPWR o[61] sky130_fd_sc_hd__buf_2
Xoutput353 net353 VGND VGND VPWR VPWR o[71] sky130_fd_sc_hd__buf_2
Xoutput364 net364 VGND VGND VPWR VPWR o[81] sky130_fd_sc_hd__buf_2
Xoutput375 net375 VGND VGND VPWR VPWR o[91] sky130_fd_sc_hd__buf_2
XFILLER_0_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_61_3 pp_row61_23 pp_row61_24 pp_row61_25 VGND VGND VPWR VPWR c$552 s$553
+ sky130_fd_sc_hd__fa_1
XFILLER_75_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_54_2 pp_row54_11 pp_row54_12 pp_row54_13 VGND VGND VPWR VPWR c$424 s$425
+ sky130_fd_sc_hd__fa_1
Xdadda_fa_4_31_1 c$2082 c$2084 s$2087 VGND VGND VPWR VPWR c$2878 s$2879 sky130_fd_sc_hd__fa_1
XFILLER_28_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_47_1 pp_row47_3 pp_row47_4 pp_row47_5 VGND VGND VPWR VPWR c$304 s$305
+ sky130_fd_sc_hd__fa_1
XFILLER_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_24_0 s$1057 c$2022 c$2024 VGND VGND VPWR VPWR c$2834 s$2835 sky130_fd_sc_hd__fa_1
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_578 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_76_3 s$1643 s$1645 s$1647 VGND VGND VPWR VPWR c$2452 s$2453 sky130_fd_sc_hd__fa_1
XFILLER_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1501 net1502 VGND VGND VPWR VPWR net1501 sky130_fd_sc_hd__clkbuf_8
XFILLER_133_992 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1512 net1514 VGND VGND VPWR VPWR net1512 sky130_fd_sc_hd__clkbuf_2
Xdadda_fa_3_69_2 c$1552 s$1555 s$1557 VGND VGND VPWR VPWR c$2394 s$2395 sky130_fd_sc_hd__fa_1
Xfanout1523 net1524 VGND VGND VPWR VPWR net1523 sky130_fd_sc_hd__buf_4
Xfanout1534 net124 VGND VGND VPWR VPWR net1534 sky130_fd_sc_hd__buf_4
XFILLER_120_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1545 net1546 VGND VGND VPWR VPWR net1545 sky130_fd_sc_hd__buf_2
XU$$4004 t$6451 net1283 VGND VGND VPWR VPWR booth_b58_m12 sky130_fd_sc_hd__xor2_1
Xfanout1556 net1557 VGND VGND VPWR VPWR net1556 sky130_fd_sc_hd__buf_4
XFILLER_24_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4015 net1152 net451 net1141 net724 VGND VGND VPWR VPWR t$6457 sky130_fd_sc_hd__a22o_1
XFILLER_65_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1567 net120 VGND VGND VPWR VPWR net1567 sky130_fd_sc_hd__buf_6
Xfanout580 net581 VGND VGND VPWR VPWR net580 sky130_fd_sc_hd__clkbuf_4
Xfanout1578 net1581 VGND VGND VPWR VPWR net1578 sky130_fd_sc_hd__buf_4
XU$$4026 t$6462 net1286 VGND VGND VPWR VPWR booth_b58_m23 sky130_fd_sc_hd__xor2_1
XU$$4037 net1052 net454 net1044 net727 VGND VGND VPWR VPWR t$6468 sky130_fd_sc_hd__a22o_1
Xfanout591 net592 VGND VGND VPWR VPWR net591 sky130_fd_sc_hd__buf_4
Xfanout1589 net1594 VGND VGND VPWR VPWR net1589 sky130_fd_sc_hd__buf_2
Xdadda_fa_6_39_0 c$3548 c$3550 s$3553 VGND VGND VPWR VPWR c$3974 s$3975 sky130_fd_sc_hd__fa_1
XU$$3303 t$6093 net1343 VGND VGND VPWR VPWR booth_b48_m4 sky130_fd_sc_hd__xor2_1
XU$$4048 t$6473 net1289 VGND VGND VPWR VPWR booth_b58_m34 sky130_fd_sc_hd__xor2_1
XFILLER_76_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4059 net945 net457 net929 net730 VGND VGND VPWR VPWR t$6479 sky130_fd_sc_hd__a22o_1
XU$$3314 net1497 net496 net1223 net769 VGND VGND VPWR VPWR t$6099 sky130_fd_sc_hd__a22o_1
XFILLER_46_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3325 t$6104 net1338 VGND VGND VPWR VPWR booth_b48_m15 sky130_fd_sc_hd__xor2_1
XU$$3336 net1121 net500 net1113 net773 VGND VGND VPWR VPWR t$6110 sky130_fd_sc_hd__a22o_1
XU$$2602 net1411 VGND VGND VPWR VPWR notsign$5734 sky130_fd_sc_hd__inv_1
XU$$3347 t$6115 net1338 VGND VGND VPWR VPWR booth_b48_m26 sky130_fd_sc_hd__xor2_1
XFILLER_111_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2613 net1123 net544 net1033 net817 VGND VGND VPWR VPWR t$5741 sky130_fd_sc_hd__a22o_1
XU$$3358 net1019 net495 net1002 net768 VGND VGND VPWR VPWR t$6121 sky130_fd_sc_hd__a22o_1
XU$$3369 t$6126 net1341 VGND VGND VPWR VPWR booth_b48_m37 sky130_fd_sc_hd__xor2_1
XFILLER_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2624 t$5746 net1395 VGND VGND VPWR VPWR booth_b38_m7 sky130_fd_sc_hd__xor2_1
XU$$2635 net1206 net549 net1199 net822 VGND VGND VPWR VPWR t$5752 sky130_fd_sc_hd__a22o_1
XFILLER_74_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1901 net1605 net599 net1597 net872 VGND VGND VPWR VPWR t$5376 sky130_fd_sc_hd__a22o_1
XU$$2646 t$5757 net1399 VGND VGND VPWR VPWR booth_b38_m18 sky130_fd_sc_hd__xor2_1
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1912 t$5381 net1465 VGND VGND VPWR VPWR booth_b26_m62 sky130_fd_sc_hd__xor2_1
XU$$2657 net1096 net546 net1087 net819 VGND VGND VPWR VPWR t$5763 sky130_fd_sc_hd__a22o_1
XU$$2668 t$5768 net1402 VGND VGND VPWR VPWR booth_b38_m29 sky130_fd_sc_hd__xor2_1
XU$$1923 net21 net1464 VGND VGND VPWR VPWR sel_1$5388 sky130_fd_sc_hd__xor2_2
XFILLER_61_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1934 net1675 net588 net1565 net861 VGND VGND VPWR VPWR t$5394 sky130_fd_sc_hd__a22o_1
XU$$2679 net983 net544 net974 net817 VGND VGND VPWR VPWR t$5774 sky130_fd_sc_hd__a22o_1
XFILLER_62_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1945 t$5399 net1448 VGND VGND VPWR VPWR booth_b28_m10 sky130_fd_sc_hd__xor2_1
XFILLER_15_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1956 net1166 net585 net1157 net858 VGND VGND VPWR VPWR t$5405 sky130_fd_sc_hd__a22o_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1967 t$5410 net1449 VGND VGND VPWR VPWR booth_b28_m21 sky130_fd_sc_hd__xor2_1
X_1950_ clknet_leaf_164_clk booth_b60_m64 VGND VGND VPWR VPWR pp_row124_1 sky130_fd_sc_hd__dfxtp_1
XU$$1978 net1067 net587 net1057 net860 VGND VGND VPWR VPWR t$5416 sky130_fd_sc_hd__a22o_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1989 t$5421 net1450 VGND VGND VPWR VPWR booth_b28_m32 sky130_fd_sc_hd__xor2_1
XFILLER_187_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0901_ clknet_leaf_194_clk net251 VGND VGND VPWR VPWR pp_row95_18 sky130_fd_sc_hd__dfxtp_4
X_1881_ clknet_leaf_25_clk booth_b50_m1 VGND VGND VPWR VPWR pp_row51_25 sky130_fd_sc_hd__dfxtp_1
XFILLER_119_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0832_ clknet_leaf_132_clk booth_b62_m57 VGND VGND VPWR VPWR pp_row119_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0763_ clknet_leaf_161_clk booth_b58_m31 VGND VGND VPWR VPWR pp_row89_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_115_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2502_ clknet_leaf_125_clk booth_b58_m54 VGND VGND VPWR VPWR pp_row112_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0694_ clknet_leaf_175_clk notsign$5244 VGND VGND VPWR VPWR pp_row87_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2433_ clknet_leaf_96_clk booth_b46_m21 VGND VGND VPWR VPWR pp_row67_23 sky130_fd_sc_hd__dfxtp_1
XFILLER_97_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_71_2 c$718 c$720 c$722 VGND VGND VPWR VPWR c$1582 s$1583 sky130_fd_sc_hd__fa_1
X_2364_ clknet_leaf_74_clk booth_b56_m9 VGND VGND VPWR VPWR pp_row65_28 sky130_fd_sc_hd__dfxtp_1
XFILLER_9_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_64_1 c$586 c$588 c$590 VGND VGND VPWR VPWR c$1496 s$1497 sky130_fd_sc_hd__fa_1
XFILLER_111_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$608 final_adder.p_new$620 final_adder.p_new$612 VGND VGND VPWR VPWR
+ final_adder.p_new$736 sky130_fd_sc_hd__and2_1
X_1315_ clknet_leaf_246_clk booth_b0_m29 VGND VGND VPWR VPWR pp_row29_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_56_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2295_ clknet_leaf_209_clk booth_b62_m1 VGND VGND VPWR VPWR pp_row63_31 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_41_0 c$2930 c$2932 c$2934 VGND VGND VPWR VPWR c$3560 s$3561 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$619 final_adder.p_new$622 final_adder.g_new$631 final_adder.g_new$623
+ VGND VGND VPWR VPWR final_adder.g_new$747 sky130_fd_sc_hd__a21o_2
XFILLER_116_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_57_0 s$23 c$456 c$458 VGND VGND VPWR VPWR c$1410 s$1411 sky130_fd_sc_hd__fa_1
X_1246_ clknet_leaf_10_clk booth_b0_m25 VGND VGND VPWR VPWR pp_row25_0 sky130_fd_sc_hd__dfxtp_1
XU$$30 net1218 net446 net1207 net688 VGND VGND VPWR VPWR t$4422 sky130_fd_sc_hd__a22o_1
XFILLER_37_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$41 t$4427 net1569 VGND VGND VPWR VPWR booth_b0_m17 sky130_fd_sc_hd__xor2_1
XU$$52 net1100 net448 net1091 net690 VGND VGND VPWR VPWR t$4433 sky130_fd_sc_hd__a22o_1
XFILLER_25_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1177_ clknet_leaf_50_clk booth_b8_m12 VGND VGND VPWR VPWR pp_row20_4 sky130_fd_sc_hd__dfxtp_1
XU$$63 t$4438 net1568 VGND VGND VPWR VPWR booth_b0_m28 sky130_fd_sc_hd__xor2_1
XU$$74 net992 net448 net987 net690 VGND VGND VPWR VPWR t$4444 sky130_fd_sc_hd__a22o_1
XU$$3870 net1197 net460 net1178 net733 VGND VGND VPWR VPWR t$6383 sky130_fd_sc_hd__a22o_1
XU$$85 t$4449 net1575 VGND VGND VPWR VPWR booth_b0_m39 sky130_fd_sc_hd__xor2_1
XU$$3881 t$6388 net1291 VGND VGND VPWR VPWR booth_b56_m19 sky130_fd_sc_hd__xor2_1
XU$$96 net1721 net445 net1712 net687 VGND VGND VPWR VPWR t$4455 sky130_fd_sc_hd__a22o_1
XU$$3892 net1085 net463 net1077 net736 VGND VGND VPWR VPWR t$6394 sky130_fd_sc_hd__a22o_1
XFILLER_24_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_10 final_adder.g_new$987 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 sel_1$4478 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_32 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_43 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_54 net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_65 net414 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_76 net467 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_87 net518 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_98 net542 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_86_2 s$2529 s$2531 s$2533 VGND VGND VPWR VPWR c$3210 s$3211 sky130_fd_sc_hd__fa_1
XFILLER_134_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_79_1 c$2466 c$2468 s$2471 VGND VGND VPWR VPWR c$3166 s$3167 sky130_fd_sc_hd__fa_1
Xdadda_fa_7_56_0 s$3623 c$4006 s$4009 VGND VGND VPWR VPWR c$4264 s$4265 sky130_fd_sc_hd__fa_1
XFILLER_0_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1208 net1641 net650 net1633 net923 VGND VGND VPWR VPWR t$5022 sky130_fd_sc_hd__a22o_1
XU$$1219 t$5027 net1012 VGND VGND VPWR VPWR booth_b16_m58 sky130_fd_sc_hd__xor2_1
XFILLER_44_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_798 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1002 final_adder.$signal$1131 final_adder.g_new$1069 VGND VGND VPWR
+ VPWR net320 sky130_fd_sc_hd__xor2_2
XFILLER_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1013 final_adder.$signal$107 final_adder.g_new$943 VGND VGND VPWR
+ VPWR net332 sky130_fd_sc_hd__xor2_2
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1024 final_adder.$signal$1153 final_adder.g_new$1058 VGND VGND VPWR
+ VPWR net344 sky130_fd_sc_hd__xor2_2
XFILLER_156_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1035 final_adder.$signal$1164 final_adder.g_new$1017 VGND VGND VPWR
+ VPWR net356 sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$1046 final_adder.$signal$1175 final_adder.g_new$1047 VGND VGND VPWR
+ VPWR net368 sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$1057 final_adder.$signal$1186 final_adder.g_new$995 VGND VGND VPWR
+ VPWR net380 sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$1068 final_adder.$signal$1197 final_adder.g_new$1036 VGND VGND VPWR
+ VPWR net265 sky130_fd_sc_hd__xor2_2
XFILLER_125_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1079 final_adder.$signal$1208 final_adder.g_new$973 VGND VGND VPWR
+ VPWR net277 sky130_fd_sc_hd__xor2_2
Xdadda_fa_3_81_1 c$1690 c$1692 c$1694 VGND VGND VPWR VPWR c$2488 s$2489 sky130_fd_sc_hd__fa_1
XFILLER_178_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_74_0 s$797 c$1602 c$1604 VGND VGND VPWR VPWR c$2430 s$2431 sky130_fd_sc_hd__fa_1
XFILLER_106_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1320 net1328 VGND VGND VPWR VPWR net1320 sky130_fd_sc_hd__clkbuf_4
Xfanout1331 net1332 VGND VGND VPWR VPWR net1331 sky130_fd_sc_hd__buf_6
Xfanout1342 net1347 VGND VGND VPWR VPWR net1342 sky130_fd_sc_hd__clkbuf_4
XFILLER_94_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1353 net1354 VGND VGND VPWR VPWR net1353 sky130_fd_sc_hd__buf_6
Xfanout1364 net1365 VGND VGND VPWR VPWR net1364 sky130_fd_sc_hd__buf_6
Xfanout1375 net38 VGND VGND VPWR VPWR net1375 sky130_fd_sc_hd__buf_6
X_1100_ clknet_leaf_52_clk booth_b12_m1 VGND VGND VPWR VPWR pp_row13_6 sky130_fd_sc_hd__dfxtp_1
Xfanout1386 net1393 VGND VGND VPWR VPWR net1386 sky130_fd_sc_hd__buf_6
X_2080_ clknet_leaf_86_clk booth_b0_m58 VGND VGND VPWR VPWR pp_row58_0 sky130_fd_sc_hd__dfxtp_1
XU$$3100 net942 net512 net926 net785 VGND VGND VPWR VPWR t$5989 sky130_fd_sc_hd__a22o_1
XFILLER_4_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1397 net1398 VGND VGND VPWR VPWR net1397 sky130_fd_sc_hd__buf_6
XU$$3111 t$5994 net1360 VGND VGND VPWR VPWR booth_b44_m45 sky130_fd_sc_hd__xor2_1
XU$$3122 net1658 net514 net1650 net787 VGND VGND VPWR VPWR t$6000 sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_110_1 c$2714 c$2716 s$2719 VGND VGND VPWR VPWR c$3352 s$3353 sky130_fd_sc_hd__fa_1
XU$$3133 t$6005 net1364 VGND VGND VPWR VPWR booth_b44_m56 sky130_fd_sc_hd__xor2_1
X_1031_ clknet_leaf_61_clk booth_b2_m2 VGND VGND VPWR VPWR pp_row4_1 sky130_fd_sc_hd__dfxtp_1
XU$$3144 net1548 net516 net1540 net789 VGND VGND VPWR VPWR t$6011 sky130_fd_sc_hd__a22o_1
XFILLER_19_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3155 notblock$6015\[2\] net41 net1361 t$6016 notblock$6015\[0\] VGND VGND VPWR
+ VPWR sel_0$6017 sky130_fd_sc_hd__a32o_1
XU$$2410 t$5636 net1425 VGND VGND VPWR VPWR booth_b34_m37 sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_36_5 pp_row36_20 c$206 s$209 VGND VGND VPWR VPWR c$1168 s$1169 sky130_fd_sc_hd__fa_1
XU$$3166 t$6023 net1353 VGND VGND VPWR VPWR booth_b46_m4 sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_103_0 s$1955 c$2654 c$2656 VGND VGND VPWR VPWR c$3308 s$3309 sky130_fd_sc_hd__fa_1
XU$$2421 net1738 net565 net1730 net838 VGND VGND VPWR VPWR t$5642 sky130_fd_sc_hd__a22o_1
XU$$2432 t$5647 net1426 VGND VGND VPWR VPWR booth_b34_m48 sky130_fd_sc_hd__xor2_1
XFILLER_59_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3177 net1501 net506 net1226 net779 VGND VGND VPWR VPWR t$6029 sky130_fd_sc_hd__a22o_1
XFILLER_146_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3188 t$6034 net1348 VGND VGND VPWR VPWR booth_b46_m15 sky130_fd_sc_hd__xor2_1
XU$$2443 net1632 net566 net1622 net839 VGND VGND VPWR VPWR t$5653 sky130_fd_sc_hd__a22o_1
XFILLER_179_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2454 t$5658 net1428 VGND VGND VPWR VPWR booth_b34_m59 sky130_fd_sc_hd__xor2_1
XU$$3199 net1121 net506 net1113 net779 VGND VGND VPWR VPWR t$6040 sky130_fd_sc_hd__a22o_1
XU$$1720 net983 net604 net974 net877 VGND VGND VPWR VPWR t$5284 sky130_fd_sc_hd__a22o_1
XU$$2465 net1429 VGND VGND VPWR VPWR notsign$5664 sky130_fd_sc_hd__inv_1
XFILLER_146_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2476 net1122 net551 net1031 net824 VGND VGND VPWR VPWR t$5671 sky130_fd_sc_hd__a22o_1
XU$$1731 t$5289 net1470 VGND VGND VPWR VPWR booth_b24_m40 sky130_fd_sc_hd__xor2_1
XU$$2487 t$5676 net1403 VGND VGND VPWR VPWR booth_b36_m7 sky130_fd_sc_hd__xor2_1
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1742 net1715 net609 net1706 net882 VGND VGND VPWR VPWR t$5295 sky130_fd_sc_hd__a22o_1
XFILLER_34_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1753 t$5300 net1473 VGND VGND VPWR VPWR booth_b24_m51 sky130_fd_sc_hd__xor2_1
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2498 net1204 net552 net1195 net825 VGND VGND VPWR VPWR t$5682 sky130_fd_sc_hd__a22o_1
XU$$1764 net1605 net608 net1597 net881 VGND VGND VPWR VPWR t$5306 sky130_fd_sc_hd__a22o_1
XU$$1775 t$5311 net1471 VGND VGND VPWR VPWR booth_b24_m62 sky130_fd_sc_hd__xor2_1
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1786 net19 net1472 VGND VGND VPWR VPWR sel_1$5318 sky130_fd_sc_hd__xor2_1
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1933_ clknet_leaf_62_clk booth_b32_m21 VGND VGND VPWR VPWR pp_row53_16 sky130_fd_sc_hd__dfxtp_1
XU$$1797 net1671 net593 net1560 net866 VGND VGND VPWR VPWR t$5324 sky130_fd_sc_hd__a22o_1
XFILLER_187_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1864_ clknet_leaf_67_clk booth_b18_m33 VGND VGND VPWR VPWR pp_row51_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_174_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_96_1 s$3267 s$3269 s$3271 VGND VGND VPWR VPWR c$3782 s$3783 sky130_fd_sc_hd__fa_1
Xinput30 a[36] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput41 a[46] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_1
X_0815_ clknet_leaf_139_clk booth_b28_m64 VGND VGND VPWR VPWR pp_row92_1 sky130_fd_sc_hd__dfxtp_1
Xinput52 a[56] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_2
XFILLER_174_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput63 a[8] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_2
X_1795_ clknet_leaf_32_clk booth_b2_m47 VGND VGND VPWR VPWR pp_row49_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_89_0 c$3218 c$3220 c$3222 VGND VGND VPWR VPWR c$3752 s$3753 sky130_fd_sc_hd__fa_1
Xinput74 b[18] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__buf_8
XFILLER_157_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput85 b[28] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_2
Xinput96 b[38] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__buf_4
X_0746_ clknet_leaf_142_clk booth_b26_m63 VGND VGND VPWR VPWR pp_row89_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_192_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0677_ clknet_leaf_131_clk booth_b62_m55 VGND VGND VPWR VPWR pp_row117_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_153_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2416_ clknet_leaf_92_clk booth_b14_m53 VGND VGND VPWR VPWR pp_row67_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_112_962 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$405 final_adder.p_new$406 final_adder.g_new$411 final_adder.g_new$407
+ VGND VGND VPWR VPWR final_adder.g_new$533 sky130_fd_sc_hd__a21o_1
XFILLER_69_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2347_ clknet_leaf_88_clk booth_b26_m39 VGND VGND VPWR VPWR pp_row65_13 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$416 final_adder.p_new$422 final_adder.p_new$418 VGND VGND VPWR VPWR
+ final_adder.p_new$544 sky130_fd_sc_hd__and2_1
XFILLER_123_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$427 final_adder.p_new$428 final_adder.g_new$433 final_adder.g_new$429
+ VGND VGND VPWR VPWR final_adder.g_new$555 sky130_fd_sc_hd__a21o_1
XTAP_3709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$438 final_adder.p_new$444 final_adder.p_new$440 VGND VGND VPWR VPWR
+ final_adder.p_new$566 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$449 final_adder.p_new$450 final_adder.g_new$455 final_adder.g_new$451
+ VGND VGND VPWR VPWR final_adder.g_new$577 sky130_fd_sc_hd__a21o_1
X_2278_ clknet_leaf_212_clk booth_b34_m29 VGND VGND VPWR VPWR pp_row63_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_72_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1229_ clknet_leaf_244_clk net172 VGND VGND VPWR VPWR pp_row23_12 sky130_fd_sc_hd__dfxtp_2
XU$$4390 net1815 sel_0$6647 net1233 net698 VGND VGND VPWR VPWR t$6649 sky130_fd_sc_hd__a22o_1
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_91_0 s$1829 c$2558 c$2560 VGND VGND VPWR VPWR c$3236 s$3237 sky130_fd_sc_hd__fa_1
XFILLER_5_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_105_2 pp_row105_12 pp_row105_13 c$1956 VGND VGND VPWR VPWR c$2682 s$2683
+ sky130_fd_sc_hd__fa_1
XFILLER_162_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_119_0 c$3868 c$3870 s$3873 VGND VGND VPWR VPWR c$4134 s$4135 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$950 final_adder.$signal$1112 final_adder.g_new$861 final_adder.$signal$46
+ VGND VGND VPWR VPWR final_adder.g_new$1078 sky130_fd_sc_hd__a21o_1
XFILLER_180_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$961 final_adder.$signal$1 net1890 VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__xor2_1
XU$$800 t$4813 net1417 VGND VGND VPWR VPWR booth_b10_m54 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$972 final_adder.$signal$1101 final_adder.g_new$1084 VGND VGND VPWR
+ VPWR net279 sky130_fd_sc_hd__xor2_2
XFILLER_28_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$811 net1582 net408 net1555 net674 VGND VGND VPWR VPWR t$4819 sky130_fd_sc_hd__a22o_1
XU$$822 net1417 VGND VGND VPWR VPWR notblock$4825\[0\] sky130_fd_sc_hd__inv_1
Xdadda_fa_3_39_3 s$1199 s$1201 s$1203 VGND VGND VPWR VPWR c$2156 s$2157 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$983 final_adder.$signal$1112 final_adder.g_new$861 VGND VGND VPWR
+ VPWR net299 sky130_fd_sc_hd__xor2_2
XU$$833 t$4831 net1312 VGND VGND VPWR VPWR booth_b12_m2 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$994 final_adder.$signal$1123 final_adder.g_new$1073 VGND VGND VPWR
+ VPWR net311 sky130_fd_sc_hd__xor2_2
XU$$844 net1515 net396 net1508 net662 VGND VGND VPWR VPWR t$4837 sky130_fd_sc_hd__a22o_1
XFILLER_73_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$855 t$4842 net1310 VGND VGND VPWR VPWR booth_b12_m13 sky130_fd_sc_hd__xor2_1
XFILLER_44_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$866 net1138 net393 net1130 net659 VGND VGND VPWR VPWR t$4848 sky130_fd_sc_hd__a22o_1
XU$$1005 net1133 net387 net1117 net653 VGND VGND VPWR VPWR t$4919 sky130_fd_sc_hd__a22o_1
XFILLER_17_979 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1016 t$4924 net1185 VGND VGND VPWR VPWR booth_b14_m25 sky130_fd_sc_hd__xor2_1
XU$$877 t$4853 net1314 VGND VGND VPWR VPWR booth_b12_m24 sky130_fd_sc_hd__xor2_1
XU$$888 net1039 net393 net1023 net659 VGND VGND VPWR VPWR t$4859 sky130_fd_sc_hd__a22o_1
XU$$1027 net1023 net388 net1015 net654 VGND VGND VPWR VPWR t$4930 sky130_fd_sc_hd__a22o_1
XU$$899 t$4864 net1311 VGND VGND VPWR VPWR booth_b12_m35 sky130_fd_sc_hd__xor2_1
XU$$1038 t$4935 net1186 VGND VGND VPWR VPWR booth_b14_m36 sky130_fd_sc_hd__xor2_1
XU$$1049 net1749 net392 net1741 net658 VGND VGND VPWR VPWR t$4941 sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_191_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_191_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_129_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0600_ clknet_leaf_188_clk booth_b40_m43 VGND VGND VPWR VPWR pp_row83_11 sky130_fd_sc_hd__dfxtp_1
X_1580_ clknet_leaf_243_clk booth_b8_m33 VGND VGND VPWR VPWR pp_row41_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_125_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0531_ clknet_leaf_162_clk notsign$5034 VGND VGND VPWR VPWR pp_row81_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_153_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0462_ clknet_leaf_157_clk booth_b50_m28 VGND VGND VPWR VPWR pp_row78_19 sky130_fd_sc_hd__dfxtp_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2201_ clknet_leaf_223_clk booth_b26_m35 VGND VGND VPWR VPWR pp_row61_13 sky130_fd_sc_hd__dfxtp_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0393_ clknet_leaf_191_clk booth_b34_m42 VGND VGND VPWR VPWR pp_row76_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1066 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1150 net1154 VGND VGND VPWR VPWR net1150 sky130_fd_sc_hd__buf_4
XFILLER_121_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_ha_2_28_3 pp_row28_9 pp_row28_10 VGND VGND VPWR VPWR c$1080 s$1081 sky130_fd_sc_hd__ha_1
XFILLER_6_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1161 net1163 VGND VGND VPWR VPWR net1161 sky130_fd_sc_hd__clkbuf_8
Xfanout1172 net71 VGND VGND VPWR VPWR net1172 sky130_fd_sc_hd__clkbuf_8
XFILLER_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2132_ clknet_leaf_32_clk booth_b30_m29 VGND VGND VPWR VPWR pp_row59_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1183 net1184 VGND VGND VPWR VPWR net1183 sky130_fd_sc_hd__buf_6
XFILLER_94_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_879 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1194 net1195 VGND VGND VPWR VPWR net1194 sky130_fd_sc_hd__buf_4
XFILLER_26_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_41_3 pp_row41_20 pp_row41_21 c$228 VGND VGND VPWR VPWR c$1224 s$1225 sky130_fd_sc_hd__fa_1
XFILLER_54_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2063_ clknet_leaf_43_clk booth_b28_m29 VGND VGND VPWR VPWR pp_row57_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_75_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_34_2 pp_row34_8 pp_row34_9 pp_row34_10 VGND VGND VPWR VPWR c$1138 s$1139
+ sky130_fd_sc_hd__fa_1
X_1014_ clknet_leaf_182_clk net131 VGND VGND VPWR VPWR pp_row101_15 sky130_fd_sc_hd__dfxtp_4
XFILLER_35_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2240 net1118 net571 net1108 net844 VGND VGND VPWR VPWR t$5550 sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_11_1 c$2756 s$2759 s$2761 VGND VGND VPWR VPWR c$3442 s$3443 sky130_fd_sc_hd__fa_1
XU$$2251 t$5555 net1433 VGND VGND VPWR VPWR booth_b32_m26 sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_27_1 pp_row27_3 pp_row27_4 pp_row27_5 VGND VGND VPWR VPWR c$1070 s$1071
+ sky130_fd_sc_hd__fa_1
XU$$2262 net1018 net570 net1001 net843 VGND VGND VPWR VPWR t$5561 sky130_fd_sc_hd__a22o_1
XFILLER_179_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2273 t$5566 net1437 VGND VGND VPWR VPWR booth_b32_m37 sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_182_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_182_clk
+ sky130_fd_sc_hd__clkbuf_16
XU$$2284 net1739 net573 net1731 net846 VGND VGND VPWR VPWR t$5572 sky130_fd_sc_hd__a22o_1
XU$$2295 t$5577 net1434 VGND VGND VPWR VPWR booth_b32_m48 sky130_fd_sc_hd__xor2_1
XU$$1550 t$5197 net1476 VGND VGND VPWR VPWR booth_b22_m18 sky130_fd_sc_hd__xor2_1
XU$$1561 net1089 net611 net1081 net884 VGND VGND VPWR VPWR t$5203 sky130_fd_sc_hd__a22o_1
XU$$1572 t$5208 net1480 VGND VGND VPWR VPWR booth_b22_m29 sky130_fd_sc_hd__xor2_1
XFILLER_50_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1583 net987 net613 net977 net886 VGND VGND VPWR VPWR t$5214 sky130_fd_sc_hd__a22o_1
XU$$1594 t$5219 net1477 VGND VGND VPWR VPWR booth_b22_m40 sky130_fd_sc_hd__xor2_1
XFILLER_188_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1916_ clknet_leaf_138_clk booth_b64_m43 VGND VGND VPWR VPWR pp_row107_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_175_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1847_ clknet_leaf_70_clk booth_b44_m6 VGND VGND VPWR VPWR pp_row50_22 sky130_fd_sc_hd__dfxtp_1
XFILLER_162_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1778_ clknet_leaf_220_clk booth_b26_m22 VGND VGND VPWR VPWR pp_row48_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0729_ clknet_leaf_135_clk booth_b40_m48 VGND VGND VPWR VPWR pp_row88_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_131_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_79_4 pp_row79_12 pp_row79_13 pp_row79_14 VGND VGND VPWR VPWR c$878 s$879
+ sky130_fd_sc_hd__fa_1
XFILLER_98_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$202 final_adder.$signal$107 final_adder.$signal$109 VGND VGND VPWR
+ VPWR final_adder.p_new$330 sky130_fd_sc_hd__and2_1
XTAP_4229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$213 final_adder.$signal$1133 final_adder.$signal$86 final_adder.$signal$88
+ VGND VGND VPWR VPWR final_adder.g_new$341 sky130_fd_sc_hd__a21o_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$224 final_adder.$signal$1120 final_adder.$signal$1121 VGND VGND VPWR
+ VPWR final_adder.p_new$352 sky130_fd_sc_hd__and2_1
Xdadda_fa_4_49_2 s$2233 s$2235 s$2237 VGND VGND VPWR VPWR c$2988 s$2989 sky130_fd_sc_hd__fa_1
XTAP_3506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$235 final_adder.$signal$1111 final_adder.$signal$42 final_adder.$signal$44
+ VGND VGND VPWR VPWR final_adder.g_new$363 sky130_fd_sc_hd__a21o_1
XTAP_3517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$246 final_adder.$signal$1098 final_adder.$signal$1099 VGND VGND VPWR
+ VPWR final_adder.p_new$374 sky130_fd_sc_hd__and2_1
XFILLER_100_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$268 final_adder.p_new$270 final_adder.p_new$268 VGND VGND VPWR VPWR
+ final_adder.p_new$396 sky130_fd_sc_hd__and2_1
XU$$107 t$4460 net1570 VGND VGND VPWR VPWR booth_b0_m50 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$279 final_adder.p_new$278 final_adder.g_new$281 final_adder.g_new$279
+ VGND VGND VPWR VPWR final_adder.g_new$407 sky130_fd_sc_hd__a21o_1
XFILLER_45_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$118 net1615 net449 net1607 net691 VGND VGND VPWR VPWR t$4466 sky130_fd_sc_hd__a22o_1
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$129 t$4471 net1570 VGND VGND VPWR VPWR booth_b0_m61 sky130_fd_sc_hd__xor2_1
Xdadda_fa_7_19_0 s$3475 c$3932 s$3935 VGND VGND VPWR VPWR c$4190 s$4191 sky130_fd_sc_hd__fa_1
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$682_1884 VGND VGND VPWR VPWR U$$682_1884/HI net1884 sky130_fd_sc_hd__conb_1
XFILLER_26_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_173_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_173_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_129_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_718 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_807 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_110_0 net1909 pp_row110_1 pp_row110_2 VGND VGND VPWR VPWR c$2718 s$2719
+ sky130_fd_sc_hd__fa_1
XFILLER_175_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_1014 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput220 c[67] VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__clkbuf_1
Xinput231 c[77] VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__clkbuf_1
Xinput242 c[87] VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_51_2 c$1336 s$1339 s$1341 VGND VGND VPWR VPWR c$2250 s$2251 sky130_fd_sc_hd__fa_2
XFILLER_103_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_0_67_2 pp_row67_6 pp_row67_7 pp_row67_8 VGND VGND VPWR VPWR c$124 s$125
+ sky130_fd_sc_hd__fa_1
Xinput253 c[97] VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_44_1 c$1246 c$1248 c$1250 VGND VGND VPWR VPWR c$2192 s$2193 sky130_fd_sc_hd__fa_1
XFILLER_124_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_21_0 c$3476 c$3478 s$3481 VGND VGND VPWR VPWR c$3938 s$3939 sky130_fd_sc_hd__fa_1
Xdadda_fa_3_37_0 s$215 c$1158 c$1160 VGND VGND VPWR VPWR c$2134 s$2135 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$780 final_adder.p_new$828 final_adder.p_new$796 VGND VGND VPWR VPWR
+ final_adder.p_new$908 sky130_fd_sc_hd__and2_1
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$630 net956 net409 net948 net675 VGND VGND VPWR VPWR t$4727 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$791 final_adder.p_new$806 final_adder.g_new$839 final_adder.g_new$807
+ VGND VGND VPWR VPWR final_adder.g_new$919 sky130_fd_sc_hd__a21o_1
XU$$641 t$4732 net1242 VGND VGND VPWR VPWR booth_b8_m43 sky130_fd_sc_hd__xor2_1
XFILLER_112_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$652 net1690 net416 net1682 net682 VGND VGND VPWR VPWR t$4738 sky130_fd_sc_hd__a22o_1
XU$$663 t$4743 net1237 VGND VGND VPWR VPWR booth_b8_m54 sky130_fd_sc_hd__xor2_1
XFILLER_16_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_1004 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$674 net1582 net416 net1555 net682 VGND VGND VPWR VPWR t$4749 sky130_fd_sc_hd__a22o_1
XFILLER_32_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$685 net1238 VGND VGND VPWR VPWR notblock$4755\[0\] sky130_fd_sc_hd__inv_1
XFILLER_56_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_164_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_164_clk
+ sky130_fd_sc_hd__clkbuf_16
XU$$696 t$4761 net1414 VGND VGND VPWR VPWR booth_b10_m2 sky130_fd_sc_hd__xor2_1
XFILLER_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_913 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1701_ clknet_leaf_22_clk booth_b38_m7 VGND VGND VPWR VPWR pp_row45_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1632_ clknet_leaf_242_clk booth_b8_m35 VGND VGND VPWR VPWR pp_row43_4 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_96_4 pp_row96_14 pp_row96_15 pp_row96_16 VGND VGND VPWR VPWR c$1886 s$1887
+ sky130_fd_sc_hd__fa_1
XFILLER_172_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1563_ clknet_leaf_7_clk booth_b22_m18 VGND VGND VPWR VPWR pp_row40_11 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_89_3 pp_row89_21 c$1000 c$1002 VGND VGND VPWR VPWR c$1800 s$1801 sky130_fd_sc_hd__fa_1
XFILLER_98_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0514_ clknet_leaf_191_clk booth_b36_m44 VGND VGND VPWR VPWR pp_row80_11 sky130_fd_sc_hd__dfxtp_1
Xfanout409 net412 VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__buf_4
XFILLER_141_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1494_ clknet_leaf_122_clk notsign$5874 VGND VGND VPWR VPWR pp_row105_0 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_59_1 s$3045 s$3047 s$3049 VGND VGND VPWR VPWR c$3634 s$3635 sky130_fd_sc_hd__fa_2
XFILLER_141_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0445_ clknet_leaf_207_clk booth_b18_m60 VGND VGND VPWR VPWR pp_row78_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_98_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0376_ clknet_leaf_203_clk booth_b62_m13 VGND VGND VPWR VPWR pp_row75_26 sky130_fd_sc_hd__dfxtp_1
XFILLER_95_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2115_ clknet_leaf_218_clk booth_b0_m59 VGND VGND VPWR VPWR pp_row59_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_27_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2046_ clknet_leaf_82_clk booth_b0_m57 VGND VGND VPWR VPWR pp_row57_0 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_105_1 pp_row105_3 pp_row105_4 pp_row105_5 VGND VGND VPWR VPWR c$1964 s$1965
+ sky130_fd_sc_hd__fa_1
XFILLER_63_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_155_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_155_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_74_1126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2070 t$5463 net1441 VGND VGND VPWR VPWR booth_b30_m4 sky130_fd_sc_hd__xor2_1
XU$$2081 net1494 net577 net1219 net850 VGND VGND VPWR VPWR t$5469 sky130_fd_sc_hd__a22o_1
XU$$2092 t$5474 net1440 VGND VGND VPWR VPWR booth_b30_m15 sky130_fd_sc_hd__xor2_1
XFILLER_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1380 net1126 net629 net1036 net902 VGND VGND VPWR VPWR t$5111 sky130_fd_sc_hd__a22o_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1391 t$5116 net1485 VGND VGND VPWR VPWR booth_b20_m7 sky130_fd_sc_hd__xor2_1
XFILLER_167_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_902 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_84_2 pp_row84_6 pp_row84_7 pp_row84_8 VGND VGND VPWR VPWR c$956 s$957
+ sky130_fd_sc_hd__fa_1
XFILLER_145_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_61_1 c$2322 c$2324 s$2327 VGND VGND VPWR VPWR c$3058 s$3059 sky130_fd_sc_hd__fa_1
Xfanout910 net911 VGND VGND VPWR VPWR net910 sky130_fd_sc_hd__buf_4
XFILLER_104_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout921 net923 VGND VGND VPWR VPWR net921 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_77_1 pp_row77_6 pp_row77_7 pp_row77_8 VGND VGND VPWR VPWR c$836 s$837
+ sky130_fd_sc_hd__fa_2
Xfanout932 net934 VGND VGND VPWR VPWR net932 sky130_fd_sc_hd__clkbuf_4
XFILLER_104_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout943 net947 VGND VGND VPWR VPWR net943 sky130_fd_sc_hd__buf_4
Xfanout954 net96 VGND VGND VPWR VPWR net954 sky130_fd_sc_hd__buf_4
Xdadda_fa_4_54_0 s$1385 c$2262 c$2264 VGND VGND VPWR VPWR c$3014 s$3015 sky130_fd_sc_hd__fa_1
XTAP_4004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout965 net968 VGND VGND VPWR VPWR net965 sky130_fd_sc_hd__buf_6
XTAP_4015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout976 net981 VGND VGND VPWR VPWR net976 sky130_fd_sc_hd__buf_4
XTAP_4026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout987 net989 VGND VGND VPWR VPWR net987 sky130_fd_sc_hd__buf_4
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout998 net999 VGND VGND VPWR VPWR net998 sky130_fd_sc_hd__buf_4
XTAP_4048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_303 net421 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_314 net564 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_325 net658 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_336 net740 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_347 net865 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_358 net967 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_146_clk clknet_5_25__leaf_clk VGND VGND VPWR VPWR clknet_leaf_146_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_369 net1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$4481_1861 VGND VGND VPWR VPWR U$$4481_1861/HI net1861 sky130_fd_sc_hd__conb_1
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_99_2 c$1910 c$1912 s$1915 VGND VGND VPWR VPWR c$2634 s$2635 sky130_fd_sc_hd__fa_1
XFILLER_155_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_69_0 c$3668 c$3670 s$3673 VGND VGND VPWR VPWR c$4034 s$4035 sky130_fd_sc_hd__fa_1
XFILLER_150_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_0_72_0 net1893 pp_row72_1 pp_row72_2 VGND VGND VPWR VPWR c$172 s$173 sky130_fd_sc_hd__fa_1
XFILLER_27_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0230_ clknet_leaf_153_clk booth_b34_m37 VGND VGND VPWR VPWR pp_row71_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_62_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_996 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$460 t$4640 net1244 VGND VGND VPWR VPWR booth_b6_m21 sky130_fd_sc_hd__xor2_1
XU$$471 net1066 net429 net1057 net711 VGND VGND VPWR VPWR t$4646 sky130_fd_sc_hd__a22o_1
XU$$482 t$4651 net1245 VGND VGND VPWR VPWR booth_b6_m32 sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_137_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_137_clk
+ sky130_fd_sc_hd__clkbuf_16
XU$$493 net956 net427 net948 net709 VGND VGND VPWR VPWR t$4657 sky130_fd_sc_hd__a22o_1
XFILLER_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0994_ clknet_leaf_121_clk booth_b62_m38 VGND VGND VPWR VPWR pp_row100_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_94_1 pp_row94_8 pp_row94_9 pp_row94_10 VGND VGND VPWR VPWR c$1856 s$1857
+ sky130_fd_sc_hd__fa_1
XFILLER_105_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1615_ clknet_leaf_241_clk booth_b28_m14 VGND VGND VPWR VPWR pp_row42_14 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_71_0 c$3110 c$3112 c$3114 VGND VGND VPWR VPWR c$3680 s$3681 sky130_fd_sc_hd__fa_1
XFILLER_99_521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_87_0 pp_row87_15 pp_row87_16 pp_row87_17 VGND VGND VPWR VPWR c$1770 s$1771
+ sky130_fd_sc_hd__fa_1
X_1546_ clknet_leaf_20_clk booth_b34_m5 VGND VGND VPWR VPWR pp_row39_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_114_876 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_70_8 s$157 s$159 s$161 VGND VGND VPWR VPWR c$724 s$725 sky130_fd_sc_hd__fa_1
XFILLER_115_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1477_ clknet_leaf_38_clk booth_b36_m0 VGND VGND VPWR VPWR pp_row36_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_63_7 c$70 s$73 s$75 VGND VGND VPWR VPWR c$596 s$597 sky130_fd_sc_hd__fa_1
XFILLER_189_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0428_ clknet_leaf_207_clk booth_b42_m35 VGND VGND VPWR VPWR pp_row77_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_41_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_56_6 pp_row56_26 pp_row56_27 pp_row56_28 VGND VGND VPWR VPWR c$468 s$469
+ sky130_fd_sc_hd__fa_1
XFILLER_39_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0359_ clknet_leaf_192_clk booth_b30_m45 VGND VGND VPWR VPWR pp_row75_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_27_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_49_5 pp_row49_15 pp_row49_16 pp_row49_17 VGND VGND VPWR VPWR c$342 s$343
+ sky130_fd_sc_hd__fa_1
XFILLER_54_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_8_0 s$3431 c$3910 s$3913 VGND VGND VPWR VPWR c$4168 s$4169 sky130_fd_sc_hd__fa_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2029_ clknet_leaf_76_clk booth_b30_m26 VGND VGND VPWR VPWR pp_row56_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_128_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_128_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_35_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_86_0 s$3743 c$4066 s$4069 VGND VGND VPWR VPWR c$4324 s$4325 sky130_fd_sc_hd__fa_2
XFILLER_136_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1705 net105 VGND VGND VPWR VPWR net1705 sky130_fd_sc_hd__buf_6
XFILLER_120_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1716 net104 VGND VGND VPWR VPWR net1716 sky130_fd_sc_hd__clkbuf_2
XFILLER_46_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1727 net1728 VGND VGND VPWR VPWR net1727 sky130_fd_sc_hd__buf_6
Xfanout1738 net101 VGND VGND VPWR VPWR net1738 sky130_fd_sc_hd__buf_6
Xfanout740 sel_1$6368 VGND VGND VPWR VPWR net740 sky130_fd_sc_hd__buf_6
Xfanout1749 net1752 VGND VGND VPWR VPWR net1749 sky130_fd_sc_hd__buf_6
Xfanout751 net752 VGND VGND VPWR VPWR net751 sky130_fd_sc_hd__buf_2
XFILLER_120_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout762 net764 VGND VGND VPWR VPWR net762 sky130_fd_sc_hd__buf_4
XU$$4208 net1717 net439 net1708 net721 VGND VGND VPWR VPWR t$6555 sky130_fd_sc_hd__a22o_1
Xfanout773 sel_1$6088 VGND VGND VPWR VPWR net773 sky130_fd_sc_hd__buf_6
XU$$4219 t$6560 net1270 VGND VGND VPWR VPWR booth_b60_m51 sky130_fd_sc_hd__xor2_1
Xfanout784 net791 VGND VGND VPWR VPWR net784 sky130_fd_sc_hd__buf_4
Xfanout795 sel_1$5878 VGND VGND VPWR VPWR net795 sky130_fd_sc_hd__buf_6
XU$$3507 net959 net486 net951 net759 VGND VGND VPWR VPWR t$6197 sky130_fd_sc_hd__a22o_1
XTAP_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3518 t$6202 net1335 VGND VGND VPWR VPWR booth_b50_m43 sky130_fd_sc_hd__xor2_1
XTAP_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3529 net1693 net490 net1684 net763 VGND VGND VPWR VPWR t$6208 sky130_fd_sc_hd__a22o_1
Xdadda_fa_6_101_0 c$3796 c$3798 s$3801 VGND VGND VPWR VPWR c$4098 s$4099 sky130_fd_sc_hd__fa_1
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2806 net1043 net538 net1027 net811 VGND VGND VPWR VPWR t$5839 sky130_fd_sc_hd__a22o_1
XTAP_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_100 net550 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2817 t$5844 net1378 VGND VGND VPWR VPWR booth_b40_m35 sky130_fd_sc_hd__xor2_1
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_111 net622 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2828 net927 net538 net1748 net811 VGND VGND VPWR VPWR t$5850 sky130_fd_sc_hd__a22o_1
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2839 t$5855 net1379 VGND VGND VPWR VPWR booth_b40_m46 sky130_fd_sc_hd__xor2_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_122 net674 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_133 net710 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_119_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_119_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_57_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_144 net769 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_155 net803 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_166 net891 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_177 net931 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_188 net972 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_199 net1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_14__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_5_14__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_114_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1400_ clknet_leaf_53_clk booth_b10_m23 VGND VGND VPWR VPWR pp_row33_5 sky130_fd_sc_hd__dfxtp_1
X_2380_ clknet_leaf_127_clk booth_b56_m55 VGND VGND VPWR VPWR pp_row111_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_69_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1331_ clknet_leaf_246_clk booth_b28_m1 VGND VGND VPWR VPWR pp_row29_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_2_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_66_5 s$647 s$649 s$651 VGND VGND VPWR VPWR c$1528 s$1529 sky130_fd_sc_hd__fa_1
XFILLER_110_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1262_ clknet_leaf_2_clk booth_b0_m26 VGND VGND VPWR VPWR pp_row26_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_84_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_59_4 s$515 s$517 s$519 VGND VGND VPWR VPWR c$1442 s$1443 sky130_fd_sc_hd__fa_1
Xinput6 a[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_2
X_0213_ clknet_leaf_152_clk booth_b64_m6 VGND VGND VPWR VPWR pp_row70_30 sky130_fd_sc_hd__dfxtp_1
XFILLER_37_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1193_ clknet_leaf_51_clk booth_b12_m9 VGND VGND VPWR VPWR pp_row21_6 sky130_fd_sc_hd__dfxtp_1
XTAP_4390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$290 net1675 net531 net1565 net804 VGND VGND VPWR VPWR t$4554 sky130_fd_sc_hd__a22o_1
XFILLER_189_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0977_ clknet_leaf_180_clk booth_b64_m57 VGND VGND VPWR VPWR pp_row121_4 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$4 c$4158 s$4161 VGND VGND VPWR VPWR final_adder.$signal$10 final_adder.$signal$1094
+ sky130_fd_sc_hd__ha_1
XFILLER_146_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput310 net310 VGND VGND VPWR VPWR o[32] sky130_fd_sc_hd__buf_2
XFILLER_173_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput321 net321 VGND VGND VPWR VPWR o[42] sky130_fd_sc_hd__buf_2
XFILLER_161_746 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput332 net332 VGND VGND VPWR VPWR o[52] sky130_fd_sc_hd__buf_2
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput343 net343 VGND VGND VPWR VPWR o[62] sky130_fd_sc_hd__buf_2
Xoutput354 net354 VGND VGND VPWR VPWR o[72] sky130_fd_sc_hd__buf_2
Xoutput365 net365 VGND VGND VPWR VPWR o[82] sky130_fd_sc_hd__buf_2
XFILLER_142_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput376 net376 VGND VGND VPWR VPWR o[92] sky130_fd_sc_hd__buf_2
XFILLER_102_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1529_ clknet_leaf_18_clk booth_b2_m37 VGND VGND VPWR VPWR pp_row39_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_101_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_61_4 pp_row61_26 pp_row61_27 pp_row61_28 VGND VGND VPWR VPWR c$554 s$555
+ sky130_fd_sc_hd__fa_1
XFILLER_142_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_54_3 pp_row54_14 pp_row54_15 pp_row54_16 VGND VGND VPWR VPWR c$426 s$427
+ sky130_fd_sc_hd__fa_1
XFILLER_67_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_31_2 s$2089 s$2091 s$2093 VGND VGND VPWR VPWR c$2880 s$2881 sky130_fd_sc_hd__fa_1
Xdadda_fa_1_47_2 pp_row47_6 pp_row47_7 pp_row47_8 VGND VGND VPWR VPWR c$306 s$307
+ sky130_fd_sc_hd__fa_1
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_24_1 c$2026 c$2028 s$2031 VGND VGND VPWR VPWR c$2836 s$2837 sky130_fd_sc_hd__fa_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_17_0 pp_row17_5 pp_row17_6 pp_row17_7 VGND VGND VPWR VPWR c$2792 s$2793
+ sky130_fd_sc_hd__fa_1
XFILLER_71_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$961_1890 VGND VGND VPWR VPWR final_adder.U$$961_1890/HI net1890 sky130_fd_sc_hd__conb_1
XFILLER_42_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_857 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1502 net128 VGND VGND VPWR VPWR net1502 sky130_fd_sc_hd__buf_6
Xfanout1513 net1514 VGND VGND VPWR VPWR net1513 sky130_fd_sc_hd__buf_4
Xdadda_fa_3_69_3 s$1559 s$1561 s$1563 VGND VGND VPWR VPWR c$2396 s$2397 sky130_fd_sc_hd__fa_1
Xfanout1524 net1526 VGND VGND VPWR VPWR net1524 sky130_fd_sc_hd__buf_4
Xfanout1535 net1538 VGND VGND VPWR VPWR net1535 sky130_fd_sc_hd__buf_4
Xfanout1546 net122 VGND VGND VPWR VPWR net1546 sky130_fd_sc_hd__buf_4
Xfanout1557 net1559 VGND VGND VPWR VPWR net1557 sky130_fd_sc_hd__clkbuf_8
XU$$4005 net1205 net452 net1197 net725 VGND VGND VPWR VPWR t$6452 sky130_fd_sc_hd__a22o_1
Xfanout570 sel_0$5527 VGND VGND VPWR VPWR net570 sky130_fd_sc_hd__buf_8
Xfanout1568 net1577 VGND VGND VPWR VPWR net1568 sky130_fd_sc_hd__buf_6
XU$$4016 t$6457 net1282 VGND VGND VPWR VPWR booth_b58_m18 sky130_fd_sc_hd__xor2_1
XU$$4027 net1095 net454 net1085 net727 VGND VGND VPWR VPWR t$6463 sky130_fd_sc_hd__a22o_1
Xfanout1579 net1581 VGND VGND VPWR VPWR net1579 sky130_fd_sc_hd__buf_4
Xfanout581 net582 VGND VGND VPWR VPWR net581 sky130_fd_sc_hd__buf_6
Xfanout592 sel_0$5387 VGND VGND VPWR VPWR net592 sky130_fd_sc_hd__buf_6
XFILLER_65_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4038 t$6468 net1286 VGND VGND VPWR VPWR booth_b58_m29 sky130_fd_sc_hd__xor2_1
XFILLER_120_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3304 net1677 net497 net1566 net770 VGND VGND VPWR VPWR t$6094 sky130_fd_sc_hd__a22o_1
XU$$4049 net988 net452 net979 net725 VGND VGND VPWR VPWR t$6474 sky130_fd_sc_hd__a22o_1
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3315 t$6099 net1339 VGND VGND VPWR VPWR booth_b48_m10 sky130_fd_sc_hd__xor2_1
XU$$3326 net1172 net497 net1163 net770 VGND VGND VPWR VPWR t$6105 sky130_fd_sc_hd__a22o_1
XU$$3337 t$6110 net1343 VGND VGND VPWR VPWR booth_b48_m21 sky130_fd_sc_hd__xor2_1
XFILLER_18_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2603 net1408 VGND VGND VPWR VPWR notblock$5735\[0\] sky130_fd_sc_hd__inv_1
XFILLER_34_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3348 net1068 net494 net1060 net767 VGND VGND VPWR VPWR t$6116 sky130_fd_sc_hd__a22o_1
XU$$2614 t$5741 net1395 VGND VGND VPWR VPWR booth_b38_m2 sky130_fd_sc_hd__xor2_1
XU$$3359 t$6121 net1340 VGND VGND VPWR VPWR booth_b48_m32 sky130_fd_sc_hd__xor2_1
XFILLER_62_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2625 net1512 net543 net1504 net816 VGND VGND VPWR VPWR t$5747 sky130_fd_sc_hd__a22o_1
XU$$2636 t$5752 net1399 VGND VGND VPWR VPWR booth_b38_m13 sky130_fd_sc_hd__xor2_1
XU$$1902 t$5376 net1464 VGND VGND VPWR VPWR booth_b26_m57 sky130_fd_sc_hd__xor2_1
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2647 net1143 net544 net1134 net817 VGND VGND VPWR VPWR t$5758 sky130_fd_sc_hd__a22o_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2658 t$5763 net1397 VGND VGND VPWR VPWR booth_b38_m24 sky130_fd_sc_hd__xor2_1
XU$$1913 net1540 net600 net1532 net873 VGND VGND VPWR VPWR t$5382 sky130_fd_sc_hd__a22o_1
XU$$1924 net1769 net584 net1227 net857 VGND VGND VPWR VPWR t$5389 sky130_fd_sc_hd__a22o_1
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2669 net1045 net547 net1029 net820 VGND VGND VPWR VPWR t$5769 sky130_fd_sc_hd__a22o_1
XFILLER_15_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1935 t$5394 net1451 VGND VGND VPWR VPWR booth_b28_m5 sky130_fd_sc_hd__xor2_1
XU$$1946 net1221 net585 net1211 net858 VGND VGND VPWR VPWR t$5400 sky130_fd_sc_hd__a22o_1
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1957 t$5405 net1449 VGND VGND VPWR VPWR booth_b28_m16 sky130_fd_sc_hd__xor2_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1968 net1107 net585 net1098 net858 VGND VGND VPWR VPWR t$5411 sky130_fd_sc_hd__a22o_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1979 t$5416 net1452 VGND VGND VPWR VPWR booth_b28_m27 sky130_fd_sc_hd__xor2_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0900_ clknet_leaf_101_clk booth_b64_m31 VGND VGND VPWR VPWR pp_row95_17 sky130_fd_sc_hd__dfxtp_1
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1880_ clknet_leaf_27_clk booth_b48_m3 VGND VGND VPWR VPWR pp_row51_24 sky130_fd_sc_hd__dfxtp_1
XFILLER_186_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0831_ clknet_leaf_107_clk booth_b58_m34 VGND VGND VPWR VPWR pp_row92_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_186_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0762_ clknet_leaf_161_clk booth_b56_m33 VGND VGND VPWR VPWR pp_row89_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_143_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2501_ clknet_leaf_147_clk booth_b42_m27 VGND VGND VPWR VPWR pp_row69_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_170_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0693_ clknet_leaf_184_clk net241 VGND VGND VPWR VPWR pp_row86_23 sky130_fd_sc_hd__dfxtp_1
XFILLER_115_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2432_ clknet_leaf_96_clk booth_b44_m23 VGND VGND VPWR VPWR pp_row67_22 sky130_fd_sc_hd__dfxtp_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_71_3 c$724 s$727 s$729 VGND VGND VPWR VPWR c$1584 s$1585 sky130_fd_sc_hd__fa_1
X_2363_ clknet_leaf_98_clk booth_b54_m11 VGND VGND VPWR VPWR pp_row65_27 sky130_fd_sc_hd__dfxtp_1
XFILLER_29_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_64_2 c$592 c$594 c$596 VGND VGND VPWR VPWR c$1498 s$1499 sky130_fd_sc_hd__fa_2
X_1314_ clknet_leaf_244_clk net177 VGND VGND VPWR VPWR pp_row28_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_97_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$609 final_adder.p_new$612 final_adder.g_new$621 final_adder.g_new$613
+ VGND VGND VPWR VPWR final_adder.g_new$737 sky130_fd_sc_hd__a21o_1
XFILLER_69_579 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2294_ clknet_leaf_130_clk booth_b62_m48 VGND VGND VPWR VPWR pp_row110_9 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_41_1 s$2937 s$2939 s$2941 VGND VGND VPWR VPWR c$3562 s$3563 sky130_fd_sc_hd__fa_2
Xdadda_fa_2_57_1 c$460 c$462 c$464 VGND VGND VPWR VPWR c$1412 s$1413 sky130_fd_sc_hd__fa_2
XFILLER_110_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1245_ clknet_leaf_244_clk net173 VGND VGND VPWR VPWR pp_row24_14 sky130_fd_sc_hd__dfxtp_2
XFILLER_84_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_34_0 c$2888 c$2890 c$2892 VGND VGND VPWR VPWR c$3532 s$3533 sky130_fd_sc_hd__fa_1
XU$$20 net1524 net446 net1516 net688 VGND VGND VPWR VPWR t$4417 sky130_fd_sc_hd__a22o_1
XFILLER_110_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$31 t$4422 net1573 VGND VGND VPWR VPWR booth_b0_m12 sky130_fd_sc_hd__xor2_1
XU$$42 net1147 net442 net1139 net684 VGND VGND VPWR VPWR t$4428 sky130_fd_sc_hd__a22o_1
XFILLER_38_988 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$53 t$4433 net1575 VGND VGND VPWR VPWR booth_b0_m23 sky130_fd_sc_hd__xor2_1
XFILLER_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1176_ clknet_leaf_50_clk booth_b6_m14 VGND VGND VPWR VPWR pp_row20_3 sky130_fd_sc_hd__dfxtp_1
XU$$64 net1047 net442 net1039 net684 VGND VGND VPWR VPWR t$4439 sky130_fd_sc_hd__a22o_1
XU$$3860 net1510 net464 net1501 net737 VGND VGND VPWR VPWR t$6378 sky130_fd_sc_hd__a22o_1
XFILLER_37_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$75 t$4444 net1574 VGND VGND VPWR VPWR booth_b0_m34 sky130_fd_sc_hd__xor2_1
XFILLER_24_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3871 t$6383 net1295 VGND VGND VPWR VPWR booth_b56_m14 sky130_fd_sc_hd__xor2_1
XU$$86 net940 net442 net924 net684 VGND VGND VPWR VPWR t$4450 sky130_fd_sc_hd__a22o_1
XU$$3882 net1135 net460 net1119 net733 VGND VGND VPWR VPWR t$6389 sky130_fd_sc_hd__a22o_1
XU$$97 t$4455 net1572 VGND VGND VPWR VPWR booth_b0_m45 sky130_fd_sc_hd__xor2_1
XU$$3893 t$6394 net1294 VGND VGND VPWR VPWR booth_b56_m25 sky130_fd_sc_hd__xor2_1
XFILLER_75_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_11 final_adder.p_new$734 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_33 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_44 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_55 net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_66 net417 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_77 net467 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_88 net518 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_99 net542 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_79_2 s$2473 s$2475 s$2477 VGND VGND VPWR VPWR c$3168 s$3169 sky130_fd_sc_hd__fa_1
XFILLER_99_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_49_0 s$3595 c$3992 s$3995 VGND VGND VPWR VPWR c$4250 s$4251 sky130_fd_sc_hd__fa_2
XFILLER_82_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_52_0 pp_row52_2 pp_row52_3 pp_row52_4 VGND VGND VPWR VPWR c$384 s$385
+ sky130_fd_sc_hd__fa_2
XFILLER_44_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1209 t$5022 net1014 VGND VGND VPWR VPWR booth_b16_m53 sky130_fd_sc_hd__xor2_1
XFILLER_180_1132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_50_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_50_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_168_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$1003 final_adder.$signal$1132 final_adder.g_new$953 VGND VGND VPWR
+ VPWR net321 sky130_fd_sc_hd__xor2_2
XFILLER_184_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1014 final_adder.$signal$109 final_adder.g_new$1063 VGND VGND VPWR
+ VPWR net333 sky130_fd_sc_hd__xor2_2
XFILLER_7_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1025 final_adder.$signal$1154 final_adder.g_new$931 VGND VGND VPWR
+ VPWR net345 sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$1036 final_adder.$signal$1165 final_adder.g_new$1052 VGND VGND VPWR
+ VPWR net357 sky130_fd_sc_hd__xor2_2
XFILLER_183_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1047 final_adder.$signal$1176 final_adder.g_new$1005 VGND VGND VPWR
+ VPWR net369 sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$1058 final_adder.$signal$1187 final_adder.g_new$1041 VGND VGND VPWR
+ VPWR net381 sky130_fd_sc_hd__xor2_2
XFILLER_165_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$1069 final_adder.$signal$1198 final_adder.g_new$983 VGND VGND VPWR
+ VPWR net266 sky130_fd_sc_hd__xor2_2
XFILLER_178_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_81_2 c$1696 s$1699 s$1701 VGND VGND VPWR VPWR c$2490 s$2491 sky130_fd_sc_hd__fa_1
XFILLER_152_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_74_1 c$1606 c$1608 c$1610 VGND VGND VPWR VPWR c$2432 s$2433 sky130_fd_sc_hd__fa_1
XFILLER_140_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_51_0 c$3596 c$3598 s$3601 VGND VGND VPWR VPWR c$3998 s$3999 sky130_fd_sc_hd__fa_2
XFILLER_78_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1310 net1311 VGND VGND VPWR VPWR net1310 sky130_fd_sc_hd__buf_6
Xdadda_fa_3_67_0 s$671 c$1518 c$1520 VGND VGND VPWR VPWR c$2374 s$2375 sky130_fd_sc_hd__fa_1
Xfanout1321 net1322 VGND VGND VPWR VPWR net1321 sky130_fd_sc_hd__clkbuf_8
XFILLER_79_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1332 net47 VGND VGND VPWR VPWR net1332 sky130_fd_sc_hd__buf_8
Xfanout1343 net1346 VGND VGND VPWR VPWR net1343 sky130_fd_sc_hd__clkbuf_8
XFILLER_78_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1354 net42 VGND VGND VPWR VPWR net1354 sky130_fd_sc_hd__buf_4
Xfanout1365 net1366 VGND VGND VPWR VPWR net1365 sky130_fd_sc_hd__buf_4
Xfanout1376 net1377 VGND VGND VPWR VPWR net1376 sky130_fd_sc_hd__buf_6
Xfanout1387 net1388 VGND VGND VPWR VPWR net1387 sky130_fd_sc_hd__buf_6
XU$$3101 t$5989 net1359 VGND VGND VPWR VPWR booth_b44_m40 sky130_fd_sc_hd__xor2_1
Xfanout1398 net33 VGND VGND VPWR VPWR net1398 sky130_fd_sc_hd__clkbuf_4
XFILLER_94_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3112 net1714 net513 net1705 net786 VGND VGND VPWR VPWR t$5995 sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_110_2 s$2721 s$2723 s$2725 VGND VGND VPWR VPWR c$3354 s$3355 sky130_fd_sc_hd__fa_1
XU$$3123 t$6000 net1363 VGND VGND VPWR VPWR booth_b44_m51 sky130_fd_sc_hd__xor2_1
X_1030_ clknet_leaf_61_clk booth_b0_m4 VGND VGND VPWR VPWR pp_row4_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3134 net1609 net516 net1602 net789 VGND VGND VPWR VPWR t$6006 sky130_fd_sc_hd__a22o_1
XU$$2400 t$5631 net1424 VGND VGND VPWR VPWR booth_b34_m32 sky130_fd_sc_hd__xor2_1
XFILLER_19_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3145 t$6011 net1365 VGND VGND VPWR VPWR booth_b44_m62 sky130_fd_sc_hd__xor2_1
XFILLER_185_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3156 net41 net1361 VGND VGND VPWR VPWR sel_1$6018 sky130_fd_sc_hd__xor2_1
XU$$2411 net958 net562 net949 net835 VGND VGND VPWR VPWR t$5637 sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_103_1 c$2658 c$2660 s$2663 VGND VGND VPWR VPWR c$3310 s$3311 sky130_fd_sc_hd__fa_1
XU$$2422 t$5642 net1425 VGND VGND VPWR VPWR booth_b34_m43 sky130_fd_sc_hd__xor2_1
XU$$3167 net1678 net505 net1567 net778 VGND VGND VPWR VPWR t$6024 sky130_fd_sc_hd__a22o_1
XFILLER_35_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2433 net1688 net565 net1680 net838 VGND VGND VPWR VPWR t$5648 sky130_fd_sc_hd__a22o_1
XU$$3178 t$6029 net1354 VGND VGND VPWR VPWR booth_b46_m10 sky130_fd_sc_hd__xor2_1
XFILLER_61_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3189 net1168 net502 net1160 net775 VGND VGND VPWR VPWR t$6035 sky130_fd_sc_hd__a22o_1
XU$$2444 t$5653 net1427 VGND VGND VPWR VPWR booth_b34_m54 sky130_fd_sc_hd__xor2_1
XFILLER_185_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2455 net1582 net567 net1555 net840 VGND VGND VPWR VPWR t$5659 sky130_fd_sc_hd__a22o_1
XU$$1710 net1041 net606 net1026 net879 VGND VGND VPWR VPWR t$5279 sky130_fd_sc_hd__a22o_1
XU$$2466 net1426 VGND VGND VPWR VPWR notblock$5665\[0\] sky130_fd_sc_hd__inv_1
XU$$1721 t$5284 net1468 VGND VGND VPWR VPWR booth_b24_m35 sky130_fd_sc_hd__xor2_1
XFILLER_179_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2477 t$5671 net1403 VGND VGND VPWR VPWR booth_b36_m2 sky130_fd_sc_hd__xor2_1
XFILLER_62_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1732 net928 net609 net1749 net882 VGND VGND VPWR VPWR t$5290 sky130_fd_sc_hd__a22o_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1743 t$5295 net1474 VGND VGND VPWR VPWR booth_b24_m46 sky130_fd_sc_hd__xor2_1
XFILLER_146_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2488 net1511 net551 net1503 net824 VGND VGND VPWR VPWR t$5677 sky130_fd_sc_hd__a22o_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1754 net1646 net607 net1638 net880 VGND VGND VPWR VPWR t$5301 sky130_fd_sc_hd__a22o_1
XU$$2499 t$5682 net1404 VGND VGND VPWR VPWR booth_b36_m13 sky130_fd_sc_hd__xor2_1
XFILLER_61_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1765 t$5306 net1472 VGND VGND VPWR VPWR booth_b24_m57 sky130_fd_sc_hd__xor2_1
XU$$1776 net1536 net608 net1528 net881 VGND VGND VPWR VPWR t$5312 sky130_fd_sc_hd__a22o_1
X_1932_ clknet_leaf_62_clk booth_b30_m23 VGND VGND VPWR VPWR pp_row53_15 sky130_fd_sc_hd__dfxtp_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1787 net1767 net594 net1228 net867 VGND VGND VPWR VPWR t$5319 sky130_fd_sc_hd__a22o_1
XU$$1798 t$5324 net1457 VGND VGND VPWR VPWR booth_b26_m5 sky130_fd_sc_hd__xor2_1
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_124_0 s$3895 c$4142 s$4145 VGND VGND VPWR VPWR c$4400 s$4401 sky130_fd_sc_hd__fa_1
Xclkbuf_leaf_41_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_187_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1863_ clknet_leaf_66_clk booth_b16_m35 VGND VGND VPWR VPWR pp_row51_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_147_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput20 a[27] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_6
X_0814_ clknet_leaf_194_clk net247 VGND VGND VPWR VPWR pp_row91_20 sky130_fd_sc_hd__dfxtp_2
Xinput31 a[37] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_4
Xinput42 a[47] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__buf_4
X_1794_ clknet_leaf_142_clk notsign$5944 VGND VGND VPWR VPWR pp_row107_0 sky130_fd_sc_hd__dfxtp_1
Xinput53 a[57] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput64 a[9] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_6
XFILLER_174_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_89_1 s$3225 s$3227 s$3229 VGND VGND VPWR VPWR c$3754 s$3755 sky130_fd_sc_hd__fa_1
Xinput75 b[19] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_4
XFILLER_143_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0745_ clknet_leaf_143_clk notsign$5314 VGND VGND VPWR VPWR pp_row89_0 sky130_fd_sc_hd__dfxtp_1
Xinput86 b[29] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_2
XFILLER_115_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput97 b[39] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0676_ clknet_leaf_176_clk booth_b36_m50 VGND VGND VPWR VPWR pp_row86_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_118_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2415_ clknet_leaf_92_clk booth_b12_m55 VGND VGND VPWR VPWR pp_row67_6 sky130_fd_sc_hd__dfxtp_1
X_2346_ clknet_leaf_88_clk booth_b24_m41 VGND VGND VPWR VPWR pp_row65_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_112_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$406 final_adder.p_new$412 final_adder.p_new$408 VGND VGND VPWR VPWR
+ final_adder.p_new$534 sky130_fd_sc_hd__and2_1
XFILLER_69_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$417 final_adder.p_new$418 final_adder.g_new$423 final_adder.g_new$419
+ VGND VGND VPWR VPWR final_adder.g_new$545 sky130_fd_sc_hd__a21o_1
XFILLER_29_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$428 final_adder.p_new$434 final_adder.p_new$430 VGND VGND VPWR VPWR
+ final_adder.p_new$556 sky130_fd_sc_hd__and2_1
X_2277_ clknet_leaf_212_clk booth_b32_m31 VGND VGND VPWR VPWR pp_row63_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_123_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$439 final_adder.p_new$440 final_adder.g_new$445 final_adder.g_new$441
+ VGND VGND VPWR VPWR final_adder.g_new$567 sky130_fd_sc_hd__a21o_1
XFILLER_42_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1228_ clknet_leaf_49_clk booth_b22_m1 VGND VGND VPWR VPWR pp_row23_11 sky130_fd_sc_hd__dfxtp_1
XU$$4380 t$6642 net1255 VGND VGND VPWR VPWR booth_b62_m63 sky130_fd_sc_hd__xor2_1
XU$$4391 t$6649 net1816 VGND VGND VPWR VPWR booth_b64_m0 sky130_fd_sc_hd__xor2_1
XFILLER_25_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1159_ clknet_leaf_46_clk booth_b0_m19 VGND VGND VPWR VPWR pp_row19_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_80_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3690 net1556 net483 net1549 net756 VGND VGND VPWR VPWR t$6290 sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_32_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_21_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_91_1 c$2562 c$2564 s$2567 VGND VGND VPWR VPWR c$3238 s$3239 sky130_fd_sc_hd__fa_1
XFILLER_107_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_84_0 s$1745 c$2502 c$2504 VGND VGND VPWR VPWR c$3194 s$3195 sky130_fd_sc_hd__fa_1
XFILLER_162_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_105_3 c$1958 c$1960 s$1963 VGND VGND VPWR VPWR c$2684 s$2685 sky130_fd_sc_hd__fa_1
Xclkbuf_leaf_99_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_99_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$940 final_adder.$signal$1132 final_adder.g_new$953 final_adder.$signal$86
+ VGND VGND VPWR VPWR final_adder.g_new$1068 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$951 final_adder.$signal$1110 final_adder.g_new$863 final_adder.$signal$42
+ VGND VGND VPWR VPWR final_adder.g_new$1079 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$962 final_adder.$signal$1091 final_adder.$signal VGND VGND VPWR VPWR
+ net296 sky130_fd_sc_hd__xor2_1
XFILLER_75_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$801 net1623 net407 net1615 net673 VGND VGND VPWR VPWR t$4814 sky130_fd_sc_hd__a22o_1
XU$$812 t$4819 net1419 VGND VGND VPWR VPWR booth_b10_m60 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$973 final_adder.$signal$1102 final_adder.g_new$751 VGND VGND VPWR
+ VPWR net288 sky130_fd_sc_hd__xor2_2
XFILLER_17_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$823 net4 VGND VGND VPWR VPWR notblock$4825\[1\] sky130_fd_sc_hd__inv_1
Xfinal_adder.U$$984 final_adder.$signal$1113 final_adder.g_new$1078 VGND VGND VPWR
+ VPWR net300 sky130_fd_sc_hd__xor2_2
XFILLER_28_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$834 net1032 net396 net933 net662 VGND VGND VPWR VPWR t$4832 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$995 final_adder.$signal$1124 final_adder.g_new$961 VGND VGND VPWR
+ VPWR net312 sky130_fd_sc_hd__xor2_2
XU$$845 t$4837 net1312 VGND VGND VPWR VPWR booth_b12_m8 sky130_fd_sc_hd__xor2_1
XU$$856 net1192 net393 net1173 net659 VGND VGND VPWR VPWR t$4843 sky130_fd_sc_hd__a22o_1
XU$$867 t$4848 net1310 VGND VGND VPWR VPWR booth_b12_m19 sky130_fd_sc_hd__xor2_1
XFILLER_73_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1006 t$4919 net1185 VGND VGND VPWR VPWR booth_b14_m20 sky130_fd_sc_hd__xor2_1
XFILLER_189_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4445_1843 VGND VGND VPWR VPWR U$$4445_1843/HI net1843 sky130_fd_sc_hd__conb_1
XU$$1017 net1071 net386 net1063 net652 VGND VGND VPWR VPWR t$4925 sky130_fd_sc_hd__a22o_1
XU$$878 net1083 net398 net1074 net664 VGND VGND VPWR VPWR t$4854 sky130_fd_sc_hd__a22o_1
XU$$889 t$4859 net1311 VGND VGND VPWR VPWR booth_b12_m30 sky130_fd_sc_hd__xor2_1
XU$$1028 t$4930 net1186 VGND VGND VPWR VPWR booth_b14_m31 sky130_fd_sc_hd__xor2_1
XU$$1039 net969 net389 net961 net655 VGND VGND VPWR VPWR t$4936 sky130_fd_sc_hd__a22o_1
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_23_clk clknet_5_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_169_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_99_0 c$3788 c$3790 s$3793 VGND VGND VPWR VPWR c$4094 s$4095 sky130_fd_sc_hd__fa_1
XFILLER_8_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0530_ clknet_leaf_194_clk net235 VGND VGND VPWR VPWR pp_row80_26 sky130_fd_sc_hd__dfxtp_1
XFILLER_140_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0461_ clknet_leaf_157_clk booth_b48_m30 VGND VGND VPWR VPWR pp_row78_18 sky130_fd_sc_hd__dfxtp_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2200_ clknet_leaf_228_clk booth_b24_m37 VGND VGND VPWR VPWR pp_row61_12 sky130_fd_sc_hd__dfxtp_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0392_ clknet_leaf_191_clk booth_b32_m44 VGND VGND VPWR VPWR pp_row76_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1140 net74 VGND VGND VPWR VPWR net1140 sky130_fd_sc_hd__clkbuf_4
Xfanout1151 net1153 VGND VGND VPWR VPWR net1151 sky130_fd_sc_hd__buf_4
Xfanout1162 net1163 VGND VGND VPWR VPWR net1162 sky130_fd_sc_hd__clkbuf_2
XFILLER_26_1078 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2131_ clknet_leaf_32_clk booth_b28_m31 VGND VGND VPWR VPWR pp_row59_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_152_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1173 net1174 VGND VGND VPWR VPWR net1173 sky130_fd_sc_hd__buf_4
Xfanout1184 net7 VGND VGND VPWR VPWR net1184 sky130_fd_sc_hd__buf_8
Xfanout1195 net1197 VGND VGND VPWR VPWR net1195 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_2_41_4 c$230 c$232 c$234 VGND VGND VPWR VPWR c$1226 s$1227 sky130_fd_sc_hd__fa_1
X_2062_ clknet_leaf_36_clk booth_b26_m31 VGND VGND VPWR VPWR pp_row57_13 sky130_fd_sc_hd__dfxtp_1
X_1013_ clknet_leaf_115_clk booth_b64_m37 VGND VGND VPWR VPWR pp_row101_14 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_34_3 pp_row34_11 pp_row34_12 pp_row34_13 VGND VGND VPWR VPWR c$1140 s$1141
+ sky130_fd_sc_hd__fa_1
XU$$2230 net1165 net569 net1156 net842 VGND VGND VPWR VPWR t$5545 sky130_fd_sc_hd__a22o_1
XFILLER_34_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2241 t$5550 net1433 VGND VGND VPWR VPWR booth_b32_m21 sky130_fd_sc_hd__xor2_1
XU$$2252 net1067 net572 net1058 net845 VGND VGND VPWR VPWR t$5556 sky130_fd_sc_hd__a22o_1
XU$$2263 t$5561 net1431 VGND VGND VPWR VPWR booth_b32_m32 sky130_fd_sc_hd__xor2_1
XU$$2274 net958 net573 net950 net846 VGND VGND VPWR VPWR t$5567 sky130_fd_sc_hd__a22o_1
XFILLER_179_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1540 t$5192 net1479 VGND VGND VPWR VPWR booth_b22_m13 sky130_fd_sc_hd__xor2_1
XU$$2285 t$5572 net1434 VGND VGND VPWR VPWR booth_b32_m43 sky130_fd_sc_hd__xor2_1
XFILLER_62_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1551 net1138 net610 net1130 net883 VGND VGND VPWR VPWR t$5198 sky130_fd_sc_hd__a22o_1
XU$$2296 net1688 net574 net1681 net847 VGND VGND VPWR VPWR t$5578 sky130_fd_sc_hd__a22o_1
XU$$1562 t$5203 net1476 VGND VGND VPWR VPWR booth_b22_m24 sky130_fd_sc_hd__xor2_1
XFILLER_37_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1573 net1041 net614 net1025 net887 VGND VGND VPWR VPWR t$5209 sky130_fd_sc_hd__a22o_1
XFILLER_50_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_14_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_16
XU$$1584 t$5214 net1478 VGND VGND VPWR VPWR booth_b22_m35 sky130_fd_sc_hd__xor2_1
XU$$1595 net925 net616 net1746 net889 VGND VGND VPWR VPWR t$5220 sky130_fd_sc_hd__a22o_1
XFILLER_188_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1915_ clknet_leaf_67_clk booth_b0_m53 VGND VGND VPWR VPWR pp_row53_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_187_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1846_ clknet_leaf_71_clk booth_b42_m8 VGND VGND VPWR VPWR pp_row50_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_147_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1777_ clknet_leaf_221_clk booth_b24_m24 VGND VGND VPWR VPWR pp_row48_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0728_ clknet_leaf_161_clk booth_b38_m50 VGND VGND VPWR VPWR pp_row88_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_143_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0659_ clknet_leaf_175_clk booth_b50_m35 VGND VGND VPWR VPWR pp_row85_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_103_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_79_5 pp_row79_15 pp_row79_16 pp_row79_17 VGND VGND VPWR VPWR c$880 s$881
+ sky130_fd_sc_hd__fa_1
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$203 final_adder.$signal$109 final_adder.$signal$106 final_adder.$signal$108
+ VGND VGND VPWR VPWR final_adder.g_new$331 sky130_fd_sc_hd__a21o_1
X_2329_ clknet_leaf_74_clk booth_b58_m6 VGND VGND VPWR VPWR pp_row64_29 sky130_fd_sc_hd__dfxtp_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$214 final_adder.$signal$1130 final_adder.$signal$1131 VGND VGND VPWR
+ VPWR final_adder.p_new$342 sky130_fd_sc_hd__and2_1
XFILLER_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$225 final_adder.$signal$1121 final_adder.$signal$62 final_adder.$signal$64
+ VGND VGND VPWR VPWR final_adder.g_new$353 sky130_fd_sc_hd__a21o_1
XTAP_3507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$236 final_adder.$signal$1108 final_adder.$signal$1109 VGND VGND VPWR
+ VPWR final_adder.p_new$364 sky130_fd_sc_hd__and2_1
XTAP_3518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$247 final_adder.$signal$1099 final_adder.$signal$18 final_adder.$signal$20
+ VGND VGND VPWR VPWR final_adder.g_new$375 sky130_fd_sc_hd__a21o_1
XFILLER_27_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$258 final_adder.p_new$260 final_adder.p_new$258 VGND VGND VPWR VPWR
+ final_adder.p_new$386 sky130_fd_sc_hd__and2_1
XU$$108 net1658 net449 net1649 net691 VGND VGND VPWR VPWR t$4461 sky130_fd_sc_hd__a22o_1
XFILLER_150_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$269 final_adder.p_new$268 final_adder.g_new$271 final_adder.g_new$269
+ VGND VGND VPWR VPWR final_adder.g_new$397 sky130_fd_sc_hd__a21o_1
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$119 t$4466 net1576 VGND VGND VPWR VPWR booth_b0_m56 sky130_fd_sc_hd__xor2_1
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_110_1 pp_row110_3 pp_row110_4 pp_row110_5 VGND VGND VPWR VPWR c$2720 s$2721
+ sky130_fd_sc_hd__fa_1
XFILLER_153_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4475_1858 VGND VGND VPWR VPWR U$$4475_1858/HI net1858 sky130_fd_sc_hd__conb_1
XFILLER_88_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_103_0 pp_row103_9 pp_row103_10 pp_row103_11 VGND VGND VPWR VPWR c$2662
+ s$2663 sky130_fd_sc_hd__fa_1
Xdadda_ha_0_68_5 pp_row68_15 pp_row68_16 VGND VGND VPWR VPWR c$142 s$143 sky130_fd_sc_hd__ha_1
XFILLER_150_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput210 c[58] VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkbuf_1
XFILLER_191_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput221 c[68] VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__clkbuf_1
Xinput232 c[78] VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_3_51_3 s$1343 s$1345 s$1347 VGND VGND VPWR VPWR c$2252 s$2253 sky130_fd_sc_hd__fa_2
Xinput243 c[88] VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput254 c[98] VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_0_67_3 pp_row67_9 pp_row67_10 pp_row67_11 VGND VGND VPWR VPWR c$126 s$127
+ sky130_fd_sc_hd__fa_2
Xdadda_fa_3_44_2 c$1252 s$1255 s$1257 VGND VGND VPWR VPWR c$2194 s$2195 sky130_fd_sc_hd__fa_1
XFILLER_91_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$770 final_adder.p_new$818 final_adder.p_new$786 VGND VGND VPWR VPWR
+ final_adder.p_new$898 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$781 final_adder.p_new$796 final_adder.g_new$829 final_adder.g_new$797
+ VGND VGND VPWR VPWR final_adder.g_new$909 sky130_fd_sc_hd__a21o_1
XU$$620 net998 net409 net990 net675 VGND VGND VPWR VPWR t$4722 sky130_fd_sc_hd__a22o_1
XFILLER_84_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_37_1 c$1162 c$1164 c$1166 VGND VGND VPWR VPWR c$2136 s$2137 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$792 final_adder.p_new$840 final_adder.p_new$808 VGND VGND VPWR VPWR
+ final_adder.p_new$920 sky130_fd_sc_hd__and2_1
XU$$631 t$4727 net1235 VGND VGND VPWR VPWR booth_b8_m38 sky130_fd_sc_hd__xor2_1
XU$$642 net1736 net414 net1725 net680 VGND VGND VPWR VPWR t$4733 sky130_fd_sc_hd__a22o_1
Xdadda_fa_6_14_0 c$3448 c$3450 s$3453 VGND VGND VPWR VPWR c$3924 s$3925 sky130_fd_sc_hd__fa_1
XFILLER_72_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$653 t$4738 net1242 VGND VGND VPWR VPWR booth_b8_m49 sky130_fd_sc_hd__xor2_1
XFILLER_182_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$664 net1620 net411 net1612 net677 VGND VGND VPWR VPWR t$4744 sky130_fd_sc_hd__a22o_1
XFILLER_56_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$675 t$4749 net1243 VGND VGND VPWR VPWR booth_b8_m60 sky130_fd_sc_hd__xor2_1
XU$$686 net2 VGND VGND VPWR VPWR notblock$4755\[1\] sky130_fd_sc_hd__inv_1
XU$$697 net1036 net404 net936 net670 VGND VGND VPWR VPWR t$4762 sky130_fd_sc_hd__a22o_1
XFILLER_71_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1700_ clknet_leaf_22_clk booth_b36_m9 VGND VGND VPWR VPWR pp_row45_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_12_493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1631_ clknet_leaf_246_clk booth_b6_m37 VGND VGND VPWR VPWR pp_row43_3 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_96_5 pp_row96_17 pp_row96_18 c$1046 VGND VGND VPWR VPWR c$1888 s$1889
+ sky130_fd_sc_hd__fa_1
XFILLER_193_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1562_ clknet_leaf_7_clk booth_b20_m20 VGND VGND VPWR VPWR pp_row40_10 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_89_4 c$1004 c$1006 c$1008 VGND VGND VPWR VPWR c$1802 s$1803 sky130_fd_sc_hd__fa_1
X_0513_ clknet_leaf_191_clk booth_b34_m46 VGND VGND VPWR VPWR pp_row80_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_4_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1493_ clknet_leaf_45_clk booth_b24_m13 VGND VGND VPWR VPWR pp_row37_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_140_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_3_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_16
X_0444_ clknet_leaf_131_clk booth_b52_m63 VGND VGND VPWR VPWR pp_row115_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_67_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0375_ clknet_leaf_203_clk booth_b60_m15 VGND VGND VPWR VPWR pp_row75_25 sky130_fd_sc_hd__dfxtp_1
X_2114_ clknet_leaf_231_clk net210 VGND VGND VPWR VPWR pp_row58_31 sky130_fd_sc_hd__dfxtp_2
XFILLER_39_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2045_ clknet_leaf_231_clk net208 VGND VGND VPWR VPWR pp_row56_30 sky130_fd_sc_hd__dfxtp_2
Xdadda_fa_2_32_0 pp_row32_0 pp_row32_1 pp_row32_2 VGND VGND VPWR VPWR c$1110 s$1111
+ sky130_fd_sc_hd__fa_1
XFILLER_35_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2060 net24 net1453 VGND VGND VPWR VPWR sel_1$5458 sky130_fd_sc_hd__xor2_1
XFILLER_120_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2071 net1675 net580 net1565 net853 VGND VGND VPWR VPWR t$5464 sky130_fd_sc_hd__a22o_1
XFILLER_90_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2082 t$5469 net1439 VGND VGND VPWR VPWR booth_b30_m10 sky130_fd_sc_hd__xor2_1
XFILLER_50_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2093 net1165 net577 net1156 net850 VGND VGND VPWR VPWR t$5475 sky130_fd_sc_hd__a22o_1
XFILLER_11_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1370 net1668 VGND VGND VPWR VPWR notblock$5105\[0\] sky130_fd_sc_hd__inv_1
XU$$1381 t$5111 net1487 VGND VGND VPWR VPWR booth_b20_m2 sky130_fd_sc_hd__xor2_1
XU$$1392 net1511 net627 net1503 net900 VGND VGND VPWR VPWR t$5117 sky130_fd_sc_hd__a22o_1
XFILLER_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_119_0 pp_row119_6 c$3398 c$3400 VGND VGND VPWR VPWR c$3872 s$3873 sky130_fd_sc_hd__fa_1
XFILLER_129_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1829_ clknet_leaf_34_clk booth_b12_m38 VGND VGND VPWR VPWR pp_row50_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_191_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_84_3 pp_row84_9 pp_row84_10 pp_row84_11 VGND VGND VPWR VPWR c$958 s$959
+ sky130_fd_sc_hd__fa_1
XFILLER_116_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout900 net901 VGND VGND VPWR VPWR net900 sky130_fd_sc_hd__buf_4
Xdadda_fa_4_61_2 s$2329 s$2331 s$2333 VGND VGND VPWR VPWR c$3060 s$3061 sky130_fd_sc_hd__fa_1
Xfanout911 net912 VGND VGND VPWR VPWR net911 sky130_fd_sc_hd__buf_6
Xfanout922 net923 VGND VGND VPWR VPWR net922 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_1_77_2 pp_row77_9 pp_row77_10 pp_row77_11 VGND VGND VPWR VPWR c$838 s$839
+ sky130_fd_sc_hd__fa_1
Xfanout933 net934 VGND VGND VPWR VPWR net933 sky130_fd_sc_hd__buf_4
Xfanout944 net947 VGND VGND VPWR VPWR net944 sky130_fd_sc_hd__buf_4
Xdadda_fa_4_54_1 c$2266 c$2268 s$2271 VGND VGND VPWR VPWR c$3016 s$3017 sky130_fd_sc_hd__fa_1
Xfanout955 net96 VGND VGND VPWR VPWR net955 sky130_fd_sc_hd__buf_4
XTAP_4005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout966 net968 VGND VGND VPWR VPWR net966 sky130_fd_sc_hd__buf_4
XTAP_4016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout977 net980 VGND VGND VPWR VPWR net977 sky130_fd_sc_hd__buf_6
XTAP_4027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_31_0 s$3523 c$3956 s$3959 VGND VGND VPWR VPWR c$4214 s$4215 sky130_fd_sc_hd__fa_2
XFILLER_86_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout988 net989 VGND VGND VPWR VPWR net988 sky130_fd_sc_hd__buf_6
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_47_0 s$1301 c$2206 c$2208 VGND VGND VPWR VPWR c$2972 s$2973 sky130_fd_sc_hd__fa_1
Xfanout999 net1005 VGND VGND VPWR VPWR net999 sky130_fd_sc_hd__buf_6
XTAP_4049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_304 net421 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_315 net583 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_326 net674 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_337 net765 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_348 net865 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_359 net967 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_1047 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_99_3 s$1917 s$1919 s$1921 VGND VGND VPWR VPWR c$2636 s$2637 sky130_fd_sc_hd__fa_1
XFILLER_108_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_0_72_1 pp_row72_3 pp_row72_4 pp_row72_5 VGND VGND VPWR VPWR c$174 s$175
+ sky130_fd_sc_hd__fa_1
XFILLER_0_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_65_0 pp_row0_1 pp_row65_1 pp_row65_2 VGND VGND VPWR VPWR c$96 s$97 sky130_fd_sc_hd__fa_1
XFILLER_76_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$450 t$4635 net1249 VGND VGND VPWR VPWR booth_b6_m16 sky130_fd_sc_hd__xor2_1
XTAP_3893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$461 net1105 net426 net1097 net708 VGND VGND VPWR VPWR t$4641 sky130_fd_sc_hd__a22o_1
XFILLER_51_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$472 t$4646 net1249 VGND VGND VPWR VPWR booth_b6_m27 sky130_fd_sc_hd__xor2_1
XU$$483 net1000 net431 net992 net713 VGND VGND VPWR VPWR t$4652 sky130_fd_sc_hd__a22o_1
XU$$494 t$4657 net1253 VGND VGND VPWR VPWR booth_b6_m38 sky130_fd_sc_hd__xor2_1
X_0993_ clknet_leaf_116_clk booth_b60_m40 VGND VGND VPWR VPWR pp_row100_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_158_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1614_ clknet_leaf_239_clk booth_b26_m16 VGND VGND VPWR VPWR pp_row42_13 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_94_2 pp_row94_11 pp_row94_12 pp_row94_13 VGND VGND VPWR VPWR c$1858 s$1859
+ sky130_fd_sc_hd__fa_1
XFILLER_126_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_71_1 s$3117 s$3119 s$3121 VGND VGND VPWR VPWR c$3682 s$3683 sky130_fd_sc_hd__fa_1
Xdadda_fa_2_87_1 pp_row87_18 pp_row87_19 pp_row87_20 VGND VGND VPWR VPWR c$1772 s$1773
+ sky130_fd_sc_hd__fa_1
XFILLER_99_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1545_ clknet_leaf_17_clk booth_b32_m7 VGND VGND VPWR VPWR pp_row39_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_99_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_64_0 c$3068 c$3070 c$3072 VGND VGND VPWR VPWR c$3652 s$3653 sky130_fd_sc_hd__fa_1
XFILLER_114_888 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1476_ clknet_leaf_38_clk booth_b34_m2 VGND VGND VPWR VPWR pp_row36_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_141_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0427_ clknet_leaf_207_clk booth_b40_m37 VGND VGND VPWR VPWR pp_row77_14 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_63_8 s$77 s$79 s$81 VGND VGND VPWR VPWR c$598 s$599 sky130_fd_sc_hd__fa_2
XFILLER_95_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_56_7 pp_row56_29 pp_row56_30 c$8 VGND VGND VPWR VPWR c$470 s$471 sky130_fd_sc_hd__fa_1
X_0358_ clknet_leaf_192_clk booth_b28_m47 VGND VGND VPWR VPWR pp_row75_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_39_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_49_6 pp_row49_18 pp_row49_19 pp_row49_20 VGND VGND VPWR VPWR c$344 s$345
+ sky130_fd_sc_hd__fa_1
XFILLER_27_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0289_ clknet_leaf_128_clk booth_b60_m53 VGND VGND VPWR VPWR pp_row113_6 sky130_fd_sc_hd__dfxtp_1
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2028_ clknet_leaf_76_clk booth_b28_m28 VGND VGND VPWR VPWR pp_row56_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_23_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_1_90_3 pp_row90_9 pp_row90_10 VGND VGND VPWR VPWR c$1024 s$1025 sky130_fd_sc_hd__ha_1
XFILLER_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_79_0 s$3715 c$4052 s$4055 VGND VGND VPWR VPWR c$4310 s$4311 sky130_fd_sc_hd__fa_2
XFILLER_3_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_82_0 net1897 pp_row82_1 pp_row82_2 VGND VGND VPWR VPWR c$922 s$923 sky130_fd_sc_hd__fa_1
Xfanout1706 net105 VGND VGND VPWR VPWR net1706 sky130_fd_sc_hd__buf_8
Xfanout1717 net1719 VGND VGND VPWR VPWR net1717 sky130_fd_sc_hd__buf_4
XFILLER_120_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1728 net103 VGND VGND VPWR VPWR net1728 sky130_fd_sc_hd__buf_4
Xfanout730 net731 VGND VGND VPWR VPWR net730 sky130_fd_sc_hd__clkbuf_4
XFILLER_49_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout741 net744 VGND VGND VPWR VPWR net741 sky130_fd_sc_hd__buf_6
Xfanout1739 net101 VGND VGND VPWR VPWR net1739 sky130_fd_sc_hd__buf_6
Xfanout752 sel_1$6228 VGND VGND VPWR VPWR net752 sky130_fd_sc_hd__buf_4
Xfanout763 net764 VGND VGND VPWR VPWR net763 sky130_fd_sc_hd__buf_4
XU$$4209 t$6555 net1270 VGND VGND VPWR VPWR booth_b60_m46 sky130_fd_sc_hd__xor2_1
Xfanout774 net775 VGND VGND VPWR VPWR net774 sky130_fd_sc_hd__buf_4
Xfanout785 net791 VGND VGND VPWR VPWR net785 sky130_fd_sc_hd__buf_4
Xfanout796 net799 VGND VGND VPWR VPWR net796 sky130_fd_sc_hd__buf_4
XFILLER_19_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3508 t$6197 net1330 VGND VGND VPWR VPWR booth_b50_m38 sky130_fd_sc_hd__xor2_1
XTAP_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3519 net1735 net489 net1727 net762 VGND VGND VPWR VPWR t$6203 sky130_fd_sc_hd__a22o_1
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2807 t$5839 net1380 VGND VGND VPWR VPWR booth_b40_m30 sky130_fd_sc_hd__xor2_1
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_101 net550 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2818 net975 net537 net966 net810 VGND VGND VPWR VPWR t$5845 sky130_fd_sc_hd__a22o_1
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_112 net622 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2829 t$5850 net1380 VGND VGND VPWR VPWR booth_b40_m41 sky130_fd_sc_hd__xor2_1
XTAP_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_123 net674 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_134 net723 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_145 net773 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_156 net803 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_167 net895 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_178 net947 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_189 net981 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_6_81_0 c$3716 c$3718 s$3721 VGND VGND VPWR VPWR c$4058 s$4059 sky130_fd_sc_hd__fa_1
Xdadda_fa_3_97_0 c$1048 c$1878 c$1880 VGND VGND VPWR VPWR c$2614 s$2615 sky130_fd_sc_hd__fa_1
XFILLER_143_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1330_ clknet_leaf_4_clk booth_b26_m3 VGND VGND VPWR VPWR pp_row29_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_110_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1261_ clknet_leaf_248_clk net174 VGND VGND VPWR VPWR pp_row25_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_110_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_59_5 s$521 s$523 s$525 VGND VGND VPWR VPWR c$1444 s$1445 sky130_fd_sc_hd__fa_1
XFILLER_77_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0212_ clknet_leaf_145_clk booth_b62_m8 VGND VGND VPWR VPWR pp_row70_29 sky130_fd_sc_hd__dfxtp_1
XFILLER_83_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput7 a[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_8
X_1192_ clknet_leaf_52_clk booth_b10_m11 VGND VGND VPWR VPWR pp_row21_5 sky130_fd_sc_hd__dfxtp_1
XTAP_4380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$280 net1783 net531 net1231 net804 VGND VGND VPWR VPWR t$4549 sky130_fd_sc_hd__a22o_1
XFILLER_17_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$291 t$4554 net1277 VGND VGND VPWR VPWR booth_b4_m5 sky130_fd_sc_hd__xor2_1
XFILLER_32_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0976_ clknet_leaf_116_clk booth_b62_m37 VGND VGND VPWR VPWR pp_row99_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_9_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$5 c$4160 s$4163 VGND VGND VPWR VPWR final_adder.$signal$12 final_adder.$signal$1095
+ sky130_fd_sc_hd__ha_1
XFILLER_133_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput300 net300 VGND VGND VPWR VPWR o[23] sky130_fd_sc_hd__buf_2
Xoutput311 net311 VGND VGND VPWR VPWR o[33] sky130_fd_sc_hd__buf_2
Xoutput322 net322 VGND VGND VPWR VPWR o[43] sky130_fd_sc_hd__buf_2
Xoutput333 net333 VGND VGND VPWR VPWR o[53] sky130_fd_sc_hd__buf_2
XFILLER_161_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput344 net344 VGND VGND VPWR VPWR o[63] sky130_fd_sc_hd__buf_2
Xoutput355 net355 VGND VGND VPWR VPWR o[73] sky130_fd_sc_hd__buf_2
XFILLER_114_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput366 net366 VGND VGND VPWR VPWR o[83] sky130_fd_sc_hd__buf_2
Xoutput377 net377 VGND VGND VPWR VPWR o[93] sky130_fd_sc_hd__buf_2
XFILLER_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1528_ clknet_leaf_121_clk booth_b46_m59 VGND VGND VPWR VPWR pp_row105_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_19_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1459_ clknet_leaf_40_clk booth_b4_m32 VGND VGND VPWR VPWR pp_row36_2 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_61_5 pp_row61_29 pp_row61_30 pp_row61_31 VGND VGND VPWR VPWR c$556 s$557
+ sky130_fd_sc_hd__fa_1
XFILLER_132_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_54_4 pp_row54_17 pp_row54_18 pp_row54_19 VGND VGND VPWR VPWR c$428 s$429
+ sky130_fd_sc_hd__fa_1
XFILLER_67_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_47_3 pp_row47_9 pp_row47_10 pp_row47_11 VGND VGND VPWR VPWR c$308 s$309
+ sky130_fd_sc_hd__fa_1
XFILLER_56_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_24_2 s$2033 s$2035 s$2037 VGND VGND VPWR VPWR c$2838 s$2839 sky130_fd_sc_hd__fa_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_17_1 pp_row17_8 pp_row17_9 c$1978 VGND VGND VPWR VPWR c$2794 s$2795 sky130_fd_sc_hd__fa_1
Xclkbuf_5_20__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_5_20__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_169_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1503 net1506 VGND VGND VPWR VPWR net1503 sky130_fd_sc_hd__buf_4
Xfanout1514 net1518 VGND VGND VPWR VPWR net1514 sky130_fd_sc_hd__buf_6
Xfanout1525 net1526 VGND VGND VPWR VPWR net1525 sky130_fd_sc_hd__buf_4
Xfanout1536 net1538 VGND VGND VPWR VPWR net1536 sky130_fd_sc_hd__buf_4
XFILLER_78_558 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1547 net122 VGND VGND VPWR VPWR net1547 sky130_fd_sc_hd__buf_4
Xfanout560 net562 VGND VGND VPWR VPWR net560 sky130_fd_sc_hd__buf_4
Xfanout1558 net1559 VGND VGND VPWR VPWR net1558 sky130_fd_sc_hd__buf_2
XU$$4006 t$6452 net1283 VGND VGND VPWR VPWR booth_b58_m13 sky130_fd_sc_hd__xor2_1
Xdadda_ha_3_20_3 pp_row20_9 pp_row20_10 VGND VGND VPWR VPWR c$2004 s$2005 sky130_fd_sc_hd__ha_1
Xfanout1569 net1577 VGND VGND VPWR VPWR net1569 sky130_fd_sc_hd__clkbuf_4
XU$$4017 net1142 net452 net1135 net725 VGND VGND VPWR VPWR t$6458 sky130_fd_sc_hd__a22o_1
Xfanout571 net572 VGND VGND VPWR VPWR net571 sky130_fd_sc_hd__buf_4
XU$$4028 t$6463 net1286 VGND VGND VPWR VPWR booth_b58_m24 sky130_fd_sc_hd__xor2_1
Xfanout582 net583 VGND VGND VPWR VPWR net582 sky130_fd_sc_hd__buf_6
Xfanout593 net595 VGND VGND VPWR VPWR net593 sky130_fd_sc_hd__buf_4
XFILLER_59_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4039 net1045 net453 net1028 net726 VGND VGND VPWR VPWR t$6469 sky130_fd_sc_hd__a22o_1
XU$$3305 t$6094 net1343 VGND VGND VPWR VPWR booth_b48_m5 sky130_fd_sc_hd__xor2_1
XU$$3316 net1222 net493 net1214 net766 VGND VGND VPWR VPWR t$6100 sky130_fd_sc_hd__a22o_1
XU$$3327 t$6105 net1343 VGND VGND VPWR VPWR booth_b48_m16 sky130_fd_sc_hd__xor2_1
XU$$3338 net1111 net495 net1102 net768 VGND VGND VPWR VPWR t$6111 sky130_fd_sc_hd__a22o_1
XU$$3349 t$6116 net1341 VGND VGND VPWR VPWR booth_b48_m27 sky130_fd_sc_hd__xor2_1
XU$$2604 net32 VGND VGND VPWR VPWR notblock$5735\[1\] sky130_fd_sc_hd__inv_1
XU$$2615 net1031 net543 net932 net816 VGND VGND VPWR VPWR t$5742 sky130_fd_sc_hd__a22o_1
XU$$2626 t$5747 net1395 VGND VGND VPWR VPWR booth_b38_m8 sky130_fd_sc_hd__xor2_1
XFILLER_94_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4409_1825 VGND VGND VPWR VPWR U$$4409_1825/HI net1825 sky130_fd_sc_hd__conb_1
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2637 net1199 net549 net1180 net822 VGND VGND VPWR VPWR t$5753 sky130_fd_sc_hd__a22o_1
XFILLER_18_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1903 net1597 net599 net1588 net872 VGND VGND VPWR VPWR t$5377 sky130_fd_sc_hd__a22o_1
XU$$2648 t$5758 net1402 VGND VGND VPWR VPWR booth_b38_m19 sky130_fd_sc_hd__xor2_1
XU$$2659 net1086 net544 net1076 net817 VGND VGND VPWR VPWR t$5764 sky130_fd_sc_hd__a22o_1
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1914 t$5382 net1465 VGND VGND VPWR VPWR booth_b26_m63 sky130_fd_sc_hd__xor2_1
XU$$1925 t$5389 net1448 VGND VGND VPWR VPWR booth_b28_m0 sky130_fd_sc_hd__xor2_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1936 net1565 net587 net1524 net860 VGND VGND VPWR VPWR t$5395 sky130_fd_sc_hd__a22o_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1947 t$5400 net1449 VGND VGND VPWR VPWR booth_b28_m11 sky130_fd_sc_hd__xor2_1
XFILLER_92_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1958 net1158 net585 net1147 net858 VGND VGND VPWR VPWR t$5406 sky130_fd_sc_hd__a22o_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1969 t$5411 net1449 VGND VGND VPWR VPWR booth_b28_m22 sky130_fd_sc_hd__xor2_1
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0830_ clknet_leaf_108_clk booth_b56_m36 VGND VGND VPWR VPWR pp_row92_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0761_ clknet_leaf_161_clk booth_b54_m35 VGND VGND VPWR VPWR pp_row89_15 sky130_fd_sc_hd__dfxtp_1
X_2500_ clknet_leaf_147_clk booth_b40_m29 VGND VGND VPWR VPWR pp_row69_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_115_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0692_ clknet_leaf_167_clk booth_b64_m22 VGND VGND VPWR VPWR pp_row86_22 sky130_fd_sc_hd__dfxtp_1
XFILLER_170_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2431_ clknet_leaf_96_clk booth_b42_m25 VGND VGND VPWR VPWR pp_row67_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_115_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2362_ clknet_leaf_74_clk booth_b52_m13 VGND VGND VPWR VPWR pp_row65_26 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_71_4 s$731 s$733 s$735 VGND VGND VPWR VPWR c$1586 s$1587 sky130_fd_sc_hd__fa_1
X_1313_ clknet_leaf_246_clk net1448 VGND VGND VPWR VPWR pp_row28_15 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_64_3 c$598 s$601 s$603 VGND VGND VPWR VPWR c$1500 s$1501 sky130_fd_sc_hd__fa_1
X_2293_ clknet_leaf_212_clk booth_b60_m3 VGND VGND VPWR VPWR pp_row63_30 sky130_fd_sc_hd__dfxtp_1
XFILLER_84_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1244_ clknet_leaf_14_clk net1467 VGND VGND VPWR VPWR pp_row24_13 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_57_2 c$466 c$468 c$470 VGND VGND VPWR VPWR c$1414 s$1415 sky130_fd_sc_hd__fa_1
XU$$10 net1127 net447 net1035 net689 VGND VGND VPWR VPWR t$4412 sky130_fd_sc_hd__a22o_1
XFILLER_77_591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_34_1 s$2895 s$2897 s$2899 VGND VGND VPWR VPWR c$3534 s$3535 sky130_fd_sc_hd__fa_1
XU$$21 t$4417 net1573 VGND VGND VPWR VPWR booth_b0_m7 sky130_fd_sc_hd__xor2_1
XU$$32 net1207 net447 net1199 net689 VGND VGND VPWR VPWR t$4423 sky130_fd_sc_hd__a22o_1
XFILLER_37_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$43 t$4428 net1569 VGND VGND VPWR VPWR booth_b0_m18 sky130_fd_sc_hd__xor2_1
X_1175_ clknet_leaf_45_clk booth_b4_m16 VGND VGND VPWR VPWR pp_row20_2 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_200_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_200_clk
+ sky130_fd_sc_hd__clkbuf_16
XU$$3850 net935 net460 net1674 net733 VGND VGND VPWR VPWR t$6373 sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_27_0 c$2846 c$2848 c$2850 VGND VGND VPWR VPWR c$3504 s$3505 sky130_fd_sc_hd__fa_1
XU$$54 net1089 net443 net1081 net685 VGND VGND VPWR VPWR t$4434 sky130_fd_sc_hd__a22o_1
XU$$65 t$4439 net1568 VGND VGND VPWR VPWR booth_b0_m29 sky130_fd_sc_hd__xor2_1
XU$$3861 t$6378 net1296 VGND VGND VPWR VPWR booth_b56_m9 sky130_fd_sc_hd__xor2_1
XU$$76 net987 net448 net977 net690 VGND VGND VPWR VPWR t$4445 sky130_fd_sc_hd__a22o_1
XU$$87 t$4450 net1568 VGND VGND VPWR VPWR booth_b0_m40 sky130_fd_sc_hd__xor2_1
XFILLER_37_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3872 net1178 net461 net1169 net734 VGND VGND VPWR VPWR t$6384 sky130_fd_sc_hd__a22o_1
XU$$3883 t$6389 net1291 VGND VGND VPWR VPWR booth_b56_m20 sky130_fd_sc_hd__xor2_1
XU$$98 net1711 net444 net1703 net686 VGND VGND VPWR VPWR t$4456 sky130_fd_sc_hd__a22o_1
XU$$3894 net1076 net460 net1068 net733 VGND VGND VPWR VPWR t$6395 sky130_fd_sc_hd__a22o_1
XFILLER_21_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_12 pp_row54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_23 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_34 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_45 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_56 net240 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_67 net425 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_78 net472 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_89 net526 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0959_ clknet_leaf_114_clk booth_b64_m34 VGND VGND VPWR VPWR pp_row98_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_137_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_101_0 c$3290 c$3292 c$3294 VGND VGND VPWR VPWR c$3800 s$3801 sky130_fd_sc_hd__fa_1
XFILLER_146_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_934 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_52_1 pp_row52_5 pp_row52_6 pp_row52_7 VGND VGND VPWR VPWR c$386 s$387
+ sky130_fd_sc_hd__fa_1
XFILLER_90_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_45_0 pp_row45_0 pp_row45_1 pp_row45_2 VGND VGND VPWR VPWR c$276 s$277
+ sky130_fd_sc_hd__fa_1
XFILLER_44_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_5_126_0_1920 VGND VGND VPWR VPWR net1920 dadda_ha_5_126_0_1920/LO sky130_fd_sc_hd__conb_1
XFILLER_102_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1004 final_adder.$signal$1133 final_adder.g_new$1068 VGND VGND VPWR
+ VPWR net322 sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$1015 final_adder.$signal$111 final_adder.g_new$941 VGND VGND VPWR
+ VPWR net334 sky130_fd_sc_hd__xor2_2
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1026 final_adder.$signal$1155 final_adder.g_new$1057 VGND VGND VPWR
+ VPWR net346 sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$1037 final_adder.$signal$1166 final_adder.g_new$1015 VGND VGND VPWR
+ VPWR net358 sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$1048 final_adder.$signal$1177 final_adder.g_new$1046 VGND VGND VPWR
+ VPWR net370 sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$1059 final_adder.$signal$1188 final_adder.g_new$993 VGND VGND VPWR
+ VPWR net382 sky130_fd_sc_hd__xor2_1
XFILLER_137_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_81_3 s$1703 s$1705 s$1707 VGND VGND VPWR VPWR c$2492 s$2493 sky130_fd_sc_hd__fa_1
XFILLER_11_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_74_2 c$1612 s$1615 s$1617 VGND VGND VPWR VPWR c$2434 s$2435 sky130_fd_sc_hd__fa_1
XFILLER_112_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1300 net1309 VGND VGND VPWR VPWR net1300 sky130_fd_sc_hd__buf_8
XFILLER_105_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1311 net5 VGND VGND VPWR VPWR net1311 sky130_fd_sc_hd__buf_6
Xdadda_fa_3_67_1 c$1522 c$1524 c$1526 VGND VGND VPWR VPWR c$2376 s$2377 sky130_fd_sc_hd__fa_1
Xfanout1322 net1323 VGND VGND VPWR VPWR net1322 sky130_fd_sc_hd__buf_4
Xfanout1333 net1337 VGND VGND VPWR VPWR net1333 sky130_fd_sc_hd__buf_6
Xfanout1344 net1345 VGND VGND VPWR VPWR net1344 sky130_fd_sc_hd__buf_6
Xdadda_fa_6_44_0 c$3568 c$3570 s$3573 VGND VGND VPWR VPWR c$3984 s$3985 sky130_fd_sc_hd__fa_1
Xfanout1355 net1356 VGND VGND VPWR VPWR net1355 sky130_fd_sc_hd__buf_6
XFILLER_78_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1366 net40 VGND VGND VPWR VPWR net1366 sky130_fd_sc_hd__buf_6
XFILLER_94_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1377 net1384 VGND VGND VPWR VPWR net1377 sky130_fd_sc_hd__buf_6
Xfanout390 net391 VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__clkbuf_8
Xfanout1388 net1393 VGND VGND VPWR VPWR net1388 sky130_fd_sc_hd__buf_6
Xfanout1399 net1402 VGND VGND VPWR VPWR net1399 sky130_fd_sc_hd__buf_6
XU$$3102 net926 net512 net1747 net785 VGND VGND VPWR VPWR t$5990 sky130_fd_sc_hd__a22o_1
XU$$3113 t$5995 net1360 VGND VGND VPWR VPWR booth_b44_m46 sky130_fd_sc_hd__xor2_1
XFILLER_115_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3124 net1650 net515 net1642 net788 VGND VGND VPWR VPWR t$6001 sky130_fd_sc_hd__a22o_1
XFILLER_19_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3135 t$6006 net1365 VGND VGND VPWR VPWR booth_b44_m57 sky130_fd_sc_hd__xor2_1
XU$$2401 net1001 net564 net993 net837 VGND VGND VPWR VPWR t$5632 sky130_fd_sc_hd__a22o_1
XFILLER_74_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3146 net1539 net516 net1531 net789 VGND VGND VPWR VPWR t$6012 sky130_fd_sc_hd__a22o_1
XU$$3157 net1789 net502 net1229 net775 VGND VGND VPWR VPWR t$6019 sky130_fd_sc_hd__a22o_1
XU$$2412 t$5637 net1422 VGND VGND VPWR VPWR booth_b34_m38 sky130_fd_sc_hd__xor2_1
XFILLER_185_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3168 t$6024 net1353 VGND VGND VPWR VPWR booth_b46_m5 sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_103_2 s$2665 s$2667 s$2669 VGND VGND VPWR VPWR c$3312 s$3313 sky130_fd_sc_hd__fa_1
XU$$2423 net1731 net566 net1722 net839 VGND VGND VPWR VPWR t$5643 sky130_fd_sc_hd__a22o_1
XU$$2434 t$5648 net1425 VGND VGND VPWR VPWR booth_b34_m49 sky130_fd_sc_hd__xor2_1
XU$$3179 net1226 net506 net1217 net779 VGND VGND VPWR VPWR t$6030 sky130_fd_sc_hd__a22o_1
XU$$2445 net1628 net565 net1614 net838 VGND VGND VPWR VPWR t$5654 sky130_fd_sc_hd__a22o_1
XU$$1700 net1082 net602 net1073 net875 VGND VGND VPWR VPWR t$5274 sky130_fd_sc_hd__a22o_1
XU$$1711 t$5279 net1470 VGND VGND VPWR VPWR booth_b24_m30 sky130_fd_sc_hd__xor2_1
XU$$2456 t$5659 net1428 VGND VGND VPWR VPWR booth_b34_m60 sky130_fd_sc_hd__xor2_1
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2467 net30 VGND VGND VPWR VPWR notblock$5665\[1\] sky130_fd_sc_hd__inv_1
XU$$1722 net974 net606 net965 net879 VGND VGND VPWR VPWR t$5285 sky130_fd_sc_hd__a22o_1
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2478 net1032 net551 net933 net824 VGND VGND VPWR VPWR t$5672 sky130_fd_sc_hd__a22o_1
XU$$1733 t$5290 net1474 VGND VGND VPWR VPWR booth_b24_m41 sky130_fd_sc_hd__xor2_1
XU$$2489 t$5677 net1403 VGND VGND VPWR VPWR booth_b36_m8 sky130_fd_sc_hd__xor2_1
XU$$1744 net1705 net607 net1695 net880 VGND VGND VPWR VPWR t$5296 sky130_fd_sc_hd__a22o_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1755 t$5301 net1473 VGND VGND VPWR VPWR booth_b24_m52 sky130_fd_sc_hd__xor2_1
XFILLER_15_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1766 net1597 net607 net1588 net880 VGND VGND VPWR VPWR t$5307 sky130_fd_sc_hd__a22o_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1931_ clknet_leaf_62_clk booth_b28_m25 VGND VGND VPWR VPWR pp_row53_14 sky130_fd_sc_hd__dfxtp_1
XU$$1777 t$5312 net1471 VGND VGND VPWR VPWR booth_b24_m63 sky130_fd_sc_hd__xor2_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1788 t$5319 net1457 VGND VGND VPWR VPWR booth_b26_m0 sky130_fd_sc_hd__xor2_1
XFILLER_30_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1799 net1564 net596 net1524 net869 VGND VGND VPWR VPWR t$5325 sky130_fd_sc_hd__a22o_1
XFILLER_30_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1862_ clknet_leaf_66_clk booth_b14_m37 VGND VGND VPWR VPWR pp_row51_7 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_7_117_0 s$3867 c$4128 s$4131 VGND VGND VPWR VPWR c$4386 s$4387 sky130_fd_sc_hd__fa_1
Xinput10 a[18] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_2
X_0813_ clknet_leaf_94_clk booth_b64_m27 VGND VGND VPWR VPWR pp_row91_19 sky130_fd_sc_hd__dfxtp_1
Xinput21 a[28] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput32 a[38] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dlymetal6s2s_1
X_1793_ clknet_leaf_35_clk booth_b0_m49 VGND VGND VPWR VPWR pp_row49_0 sky130_fd_sc_hd__dfxtp_1
Xinput43 a[48] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_249_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_249_clk
+ sky130_fd_sc_hd__clkbuf_16
Xinput54 a[58] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput65 b[0] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_2
Xinput76 b[1] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_6
X_0744_ clknet_leaf_131_clk booth_b60_m58 VGND VGND VPWR VPWR pp_row118_4 sky130_fd_sc_hd__dfxtp_1
Xinput87 b[2] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_4
XFILLER_155_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput98 b[3] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__buf_4
X_0675_ clknet_leaf_170_clk booth_b34_m52 VGND VGND VPWR VPWR pp_row86_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_192_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2414_ clknet_leaf_127_clk booth_b62_m49 VGND VGND VPWR VPWR pp_row111_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_143_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2345_ clknet_leaf_87_clk booth_b22_m43 VGND VGND VPWR VPWR pp_row65_11 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_62_0 s$71 c$546 c$548 VGND VGND VPWR VPWR c$1470 s$1471 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$407 final_adder.p_new$408 final_adder.g_new$413 final_adder.g_new$409
+ VGND VGND VPWR VPWR final_adder.g_new$535 sky130_fd_sc_hd__a21o_1
XFILLER_96_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_997 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$418 final_adder.p_new$424 final_adder.p_new$420 VGND VGND VPWR VPWR
+ final_adder.p_new$546 sky130_fd_sc_hd__and2_1
XFILLER_38_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2276_ clknet_leaf_213_clk booth_b30_m33 VGND VGND VPWR VPWR pp_row63_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_84_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_848 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$429 final_adder.p_new$430 final_adder.g_new$435 final_adder.g_new$431
+ VGND VGND VPWR VPWR final_adder.g_new$557 sky130_fd_sc_hd__a21o_1
X_1227_ clknet_leaf_143_clk booth_b48_m55 VGND VGND VPWR VPWR pp_row103_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_37_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4370 t$6637 net1257 VGND VGND VPWR VPWR booth_b62_m58 sky130_fd_sc_hd__xor2_1
XU$$4381 net1528 net419 net1809 net701 VGND VGND VPWR VPWR t$6643 sky130_fd_sc_hd__a22o_1
XU$$4392 net1234 sel_0$6647 net1129 net698 VGND VGND VPWR VPWR t$6650 sky130_fd_sc_hd__a22o_1
XFILLER_38_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1158_ clknet_leaf_245_clk net166 VGND VGND VPWR VPWR pp_row18_11 sky130_fd_sc_hd__dfxtp_2
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3680 net1616 net483 net1608 net756 VGND VGND VPWR VPWR t$6285 sky130_fd_sc_hd__a22o_1
XFILLER_16_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3691 t$6290 net1327 VGND VGND VPWR VPWR booth_b52_m61 sky130_fd_sc_hd__xor2_1
XFILLER_41_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1089_ clknet_leaf_59_clk booth_b10_m2 VGND VGND VPWR VPWR pp_row12_5 sky130_fd_sc_hd__dfxtp_1
XU$$2990 t$5932 net1375 VGND VGND VPWR VPWR booth_b42_m53 sky130_fd_sc_hd__xor2_1
XFILLER_40_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_91_2 s$2569 s$2571 s$2573 VGND VGND VPWR VPWR c$3240 s$3241 sky130_fd_sc_hd__fa_1
XFILLER_10_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_102_0_1905 VGND VGND VPWR VPWR net1905 dadda_fa_2_102_0_1905/LO sky130_fd_sc_hd__conb_1
Xdadda_fa_4_84_1 c$2506 c$2508 s$2511 VGND VGND VPWR VPWR c$3196 s$3197 sky130_fd_sc_hd__fa_1
XFILLER_134_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_61_0 s$3643 c$4016 s$4019 VGND VGND VPWR VPWR c$4274 s$4275 sky130_fd_sc_hd__fa_1
Xdadda_fa_4_77_0 s$1661 c$2446 c$2448 VGND VGND VPWR VPWR c$3152 s$3153 sky130_fd_sc_hd__fa_1
XFILLER_122_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$930 final_adder.$signal$1152 final_adder.g_new$933 final_adder.$signal$126
+ VGND VGND VPWR VPWR final_adder.g_new$1058 sky130_fd_sc_hd__a21o_1
XFILLER_189_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$941 final_adder.$signal$1130 final_adder.g_new$955 final_adder.$signal$82
+ VGND VGND VPWR VPWR final_adder.g_new$1069 sky130_fd_sc_hd__a21o_1
XFILLER_63_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$952 final_adder.$signal$1108 final_adder.g_new$865 final_adder.$signal$38
+ VGND VGND VPWR VPWR final_adder.g_new$1080 sky130_fd_sc_hd__a21o_1
XFILLER_169_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$963 final_adder.$signal$1092 final_adder.g_new$383 VGND VGND VPWR
+ VPWR net307 sky130_fd_sc_hd__xor2_1
XU$$802 t$4814 net1419 VGND VGND VPWR VPWR booth_b10_m55 sky130_fd_sc_hd__xor2_1
XFILLER_29_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$813 net1551 net403 net1543 net669 VGND VGND VPWR VPWR t$4820 sky130_fd_sc_hd__a22o_1
XFILLER_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$974 final_adder.$signal$1103 final_adder.g_new$1083 VGND VGND VPWR
+ VPWR net289 sky130_fd_sc_hd__xor2_2
XU$$824 net1316 VGND VGND VPWR VPWR notblock$4825\[2\] sky130_fd_sc_hd__inv_1
XFILLER_56_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$985 final_adder.$signal$1114 final_adder.g_new$859 VGND VGND VPWR
+ VPWR net301 sky130_fd_sc_hd__xor2_2
XFILLER_73_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$835 t$4832 net1312 VGND VGND VPWR VPWR booth_b12_m3 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$996 final_adder.$signal$1125 final_adder.g_new$1072 VGND VGND VPWR
+ VPWR net313 sky130_fd_sc_hd__xor2_2
XFILLER_113_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$846 net1508 net397 net1499 net663 VGND VGND VPWR VPWR t$4838 sky130_fd_sc_hd__a22o_1
XU$$857 t$4843 net1310 VGND VGND VPWR VPWR booth_b12_m14 sky130_fd_sc_hd__xor2_1
XU$$868 net1134 net396 net1118 net662 VGND VGND VPWR VPWR t$4849 sky130_fd_sc_hd__a22o_1
XU$$1007 net1117 net389 net1108 net655 VGND VGND VPWR VPWR t$4920 sky130_fd_sc_hd__a22o_1
XU$$1018 t$4925 net1183 VGND VGND VPWR VPWR booth_b14_m26 sky130_fd_sc_hd__xor2_1
XFILLER_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$879 t$4854 net1314 VGND VGND VPWR VPWR booth_b12_m25 sky130_fd_sc_hd__xor2_1
XU$$1029 net1015 net386 net998 net652 VGND VGND VPWR VPWR t$4931 sky130_fd_sc_hd__a22o_1
XFILLER_189_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0460_ clknet_leaf_157_clk booth_b46_m32 VGND VGND VPWR VPWR pp_row78_17 sky130_fd_sc_hd__dfxtp_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0391_ clknet_leaf_196_clk booth_b30_m46 VGND VGND VPWR VPWR pp_row76_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_94_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1130 net1132 VGND VGND VPWR VPWR net1130 sky130_fd_sc_hd__buf_4
Xfanout1141 net74 VGND VGND VPWR VPWR net1141 sky130_fd_sc_hd__buf_4
XFILLER_6_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2130_ clknet_leaf_29_clk booth_b26_m33 VGND VGND VPWR VPWR pp_row59_13 sky130_fd_sc_hd__dfxtp_1
Xfanout1152 net1153 VGND VGND VPWR VPWR net1152 sky130_fd_sc_hd__buf_4
XFILLER_78_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1163 net72 VGND VGND VPWR VPWR net1163 sky130_fd_sc_hd__buf_4
Xfanout1174 net1176 VGND VGND VPWR VPWR net1174 sky130_fd_sc_hd__clkbuf_4
Xfanout1185 net1187 VGND VGND VPWR VPWR net1185 sky130_fd_sc_hd__buf_6
X_2061_ clknet_leaf_164_clk booth_b62_m62 VGND VGND VPWR VPWR pp_row124_2 sky130_fd_sc_hd__dfxtp_1
Xfanout1196 net1197 VGND VGND VPWR VPWR net1196 sky130_fd_sc_hd__clkbuf_8
Xdadda_fa_2_41_5 s$237 s$239 s$241 VGND VGND VPWR VPWR c$1228 s$1229 sky130_fd_sc_hd__fa_2
XFILLER_47_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_829 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1012_ clknet_leaf_115_clk booth_b62_m39 VGND VGND VPWR VPWR pp_row101_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_19_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_34_4 pp_row34_14 pp_row34_15 pp_row34_16 VGND VGND VPWR VPWR c$1142 s$1143
+ sky130_fd_sc_hd__fa_1
XU$$2220 net1220 net569 net1210 net842 VGND VGND VPWR VPWR t$5540 sky130_fd_sc_hd__a22o_1
XU$$2231 t$5545 net1430 VGND VGND VPWR VPWR booth_b32_m16 sky130_fd_sc_hd__xor2_1
XFILLER_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2242 net1108 net571 net1101 net844 VGND VGND VPWR VPWR t$5551 sky130_fd_sc_hd__a22o_1
XFILLER_34_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2253 t$5556 net1433 VGND VGND VPWR VPWR booth_b32_m27 sky130_fd_sc_hd__xor2_1
XU$$2264 net1001 net572 net993 net845 VGND VGND VPWR VPWR t$5562 sky130_fd_sc_hd__a22o_1
XU$$1530 t$5187 net1475 VGND VGND VPWR VPWR booth_b22_m8 sky130_fd_sc_hd__xor2_1
XFILLER_50_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2275 t$5567 net1434 VGND VGND VPWR VPWR booth_b32_m38 sky130_fd_sc_hd__xor2_1
XFILLER_179_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2286 net1731 net573 net1722 net846 VGND VGND VPWR VPWR t$5573 sky130_fd_sc_hd__a22o_1
XFILLER_16_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1541 net1198 net613 net1179 net886 VGND VGND VPWR VPWR t$5193 sky130_fd_sc_hd__a22o_1
XU$$1552 t$5198 net1475 VGND VGND VPWR VPWR booth_b22_m19 sky130_fd_sc_hd__xor2_1
XU$$2297 t$5578 net1435 VGND VGND VPWR VPWR booth_b32_m49 sky130_fd_sc_hd__xor2_1
XU$$1563 net1082 net612 net1073 net885 VGND VGND VPWR VPWR t$5204 sky130_fd_sc_hd__a22o_1
XU$$1574 t$5209 net1479 VGND VGND VPWR VPWR booth_b22_m30 sky130_fd_sc_hd__xor2_1
XU$$1585 net977 net618 net965 net891 VGND VGND VPWR VPWR t$5215 sky130_fd_sc_hd__a22o_1
XFILLER_37_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1596 t$5220 net1483 VGND VGND VPWR VPWR booth_b22_m41 sky130_fd_sc_hd__xor2_1
XFILLER_147_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1914_ clknet_leaf_232_clk net204 VGND VGND VPWR VPWR pp_row52_28 sky130_fd_sc_hd__dfxtp_2
XFILLER_147_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1845_ clknet_leaf_71_clk booth_b40_m10 VGND VGND VPWR VPWR pp_row50_20 sky130_fd_sc_hd__dfxtp_1
XFILLER_175_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_94_0 c$3248 c$3250 c$3252 VGND VGND VPWR VPWR c$3772 s$3773 sky130_fd_sc_hd__fa_1
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1776_ clknet_leaf_238_clk booth_b22_m26 VGND VGND VPWR VPWR pp_row48_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0727_ clknet_leaf_161_clk booth_b36_m52 VGND VGND VPWR VPWR pp_row88_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_143_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0658_ clknet_leaf_177_clk booth_b48_m37 VGND VGND VPWR VPWR pp_row85_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_170_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_79_6 pp_row79_18 pp_row79_19 pp_row79_20 VGND VGND VPWR VPWR c$882 s$883
+ sky130_fd_sc_hd__fa_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0589_ clknet_leaf_186_clk booth_b20_m63 VGND VGND VPWR VPWR pp_row83_1 sky130_fd_sc_hd__dfxtp_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$204 final_adder.$signal$103 final_adder.$signal$105 VGND VGND VPWR
+ VPWR final_adder.p_new$332 sky130_fd_sc_hd__and2_1
X_2328_ clknet_leaf_74_clk booth_b56_m8 VGND VGND VPWR VPWR pp_row64_28 sky130_fd_sc_hd__dfxtp_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$215 final_adder.$signal$1131 final_adder.$signal$82 final_adder.$signal$84
+ VGND VGND VPWR VPWR final_adder.g_new$343 sky130_fd_sc_hd__a21o_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$226 final_adder.$signal$1118 final_adder.$signal$1119 VGND VGND VPWR
+ VPWR final_adder.p_new$354 sky130_fd_sc_hd__and2_1
XTAP_3508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$237 final_adder.$signal$1109 final_adder.$signal$38 final_adder.$signal$40
+ VGND VGND VPWR VPWR final_adder.g_new$365 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$248 final_adder.$signal$1096 final_adder.$signal$1097 VGND VGND VPWR
+ VPWR final_adder.p_new$376 sky130_fd_sc_hd__and2_1
XTAP_3519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$259 final_adder.p_new$258 final_adder.g_new$261 final_adder.g_new$259
+ VGND VGND VPWR VPWR final_adder.g_new$387 sky130_fd_sc_hd__a21o_1
XU$$109 t$4461 net1576 VGND VGND VPWR VPWR booth_b0_m51 sky130_fd_sc_hd__xor2_1
X_2259_ clknet_leaf_230_clk booth_b0_m63 VGND VGND VPWR VPWR pp_row63_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_26_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_110_2 pp_row110_6 pp_row110_7 pp_row110_8 VGND VGND VPWR VPWR c$2722 s$2723
+ sky130_fd_sc_hd__fa_1
XFILLER_107_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_103_1 pp_row103_12 pp_row103_13 pp_row103_14 VGND VGND VPWR VPWR c$2664
+ s$2665 sky130_fd_sc_hd__fa_1
XFILLER_104_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput200 c[49] VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__clkbuf_1
Xinput211 c[59] VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput222 c[69] VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_124_0 c$3888 c$3890 s$3893 VGND VGND VPWR VPWR c$4144 s$4145 sky130_fd_sc_hd__fa_1
Xinput233 c[79] VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput244 c[89] VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__clkbuf_1
Xinput255 c[99] VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_0_67_4 pp_row67_12 pp_row67_13 pp_row67_14 VGND VGND VPWR VPWR c$128 s$129
+ sky130_fd_sc_hd__fa_1
Xdadda_fa_3_44_3 s$1259 s$1261 s$1263 VGND VGND VPWR VPWR c$2196 s$2197 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$760 final_adder.p_new$808 final_adder.p_new$776 VGND VGND VPWR VPWR
+ final_adder.p_new$888 sky130_fd_sc_hd__and2_1
XFILLER_29_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$610 net1057 net413 net1049 net679 VGND VGND VPWR VPWR t$4717 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$771 final_adder.p_new$786 final_adder.g_new$819 final_adder.g_new$787
+ VGND VGND VPWR VPWR final_adder.g_new$899 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$782 final_adder.p_new$830 final_adder.p_new$798 VGND VGND VPWR VPWR
+ final_adder.p_new$910 sky130_fd_sc_hd__and2_1
XU$$621 t$4722 net1235 VGND VGND VPWR VPWR booth_b8_m33 sky130_fd_sc_hd__xor2_1
XFILLER_84_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_37_2 c$1168 s$1171 s$1173 VGND VGND VPWR VPWR c$2138 s$2139 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$793 final_adder.p_new$808 final_adder.g_new$841 final_adder.g_new$809
+ VGND VGND VPWR VPWR final_adder.g_new$921 sky130_fd_sc_hd__a21o_1
XU$$632 net948 net411 net940 net677 VGND VGND VPWR VPWR t$4728 sky130_fd_sc_hd__a22o_1
XFILLER_17_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$643 t$4733 net1241 VGND VGND VPWR VPWR booth_b8_m44 sky130_fd_sc_hd__xor2_1
XFILLER_189_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$654 net1682 net416 net1657 net682 VGND VGND VPWR VPWR t$4739 sky130_fd_sc_hd__a22o_1
XFILLER_186_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$665 t$4744 net1237 VGND VGND VPWR VPWR booth_b8_m55 sky130_fd_sc_hd__xor2_1
XFILLER_44_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$676 net1555 net416 net1547 net682 VGND VGND VPWR VPWR t$4750 sky130_fd_sc_hd__a22o_1
XU$$687 net1417 VGND VGND VPWR VPWR notblock$4755\[2\] sky130_fd_sc_hd__inv_1
XU$$698 t$4762 net1414 VGND VGND VPWR VPWR booth_b10_m3 sky130_fd_sc_hd__xor2_1
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2189_1772 VGND VGND VPWR VPWR U$$2189_1772/HI net1772 sky130_fd_sc_hd__conb_1
XFILLER_9_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1630_ clknet_leaf_239_clk booth_b4_m39 VGND VGND VPWR VPWR pp_row43_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1561_ clknet_leaf_108_clk booth_b52_m53 VGND VGND VPWR VPWR pp_row105_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_153_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_89_5 s$1011 s$1013 s$1015 VGND VGND VPWR VPWR c$1804 s$1805 sky130_fd_sc_hd__fa_2
X_0512_ clknet_leaf_190_clk booth_b32_m48 VGND VGND VPWR VPWR pp_row80_9 sky130_fd_sc_hd__dfxtp_1
X_1492_ clknet_leaf_45_clk booth_b22_m15 VGND VGND VPWR VPWR pp_row37_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_4_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0443_ clknet_leaf_155_clk booth_b16_m62 VGND VGND VPWR VPWR pp_row78_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_39_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_932 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0374_ clknet_leaf_204_clk booth_b58_m17 VGND VGND VPWR VPWR pp_row75_24 sky130_fd_sc_hd__dfxtp_1
XFILLER_67_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_ha_2_26_2 pp_row26_6 pp_row26_7 VGND VGND VPWR VPWR c$1066 s$1067 sky130_fd_sc_hd__ha_1
X_2113_ clknet_leaf_85_clk net1287 VGND VGND VPWR VPWR pp_row58_30 sky130_fd_sc_hd__dfxtp_1
XFILLER_94_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2044_ clknet_leaf_83_clk net1296 VGND VGND VPWR VPWR pp_row56_29 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_32_1 pp_row32_3 pp_row32_4 pp_row32_5 VGND VGND VPWR VPWR c$1112 s$1113
+ sky130_fd_sc_hd__fa_1
XFILLER_50_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_25_0 pp_row25_0 pp_row25_1 pp_row25_2 VGND VGND VPWR VPWR c$1058 s$1059
+ sky130_fd_sc_hd__fa_1
XU$$2050 net1539 net591 net1531 net864 VGND VGND VPWR VPWR t$5452 sky130_fd_sc_hd__a22o_1
Xclkbuf_5_1__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_5_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XU$$2061 net1771 net576 net1227 net849 VGND VGND VPWR VPWR t$5459 sky130_fd_sc_hd__a22o_1
XU$$2072 t$5464 net1441 VGND VGND VPWR VPWR booth_b30_m5 sky130_fd_sc_hd__xor2_1
XU$$2083 net1220 net576 net1210 net849 VGND VGND VPWR VPWR t$5470 sky130_fd_sc_hd__a22o_1
XU$$2094 t$5475 net1440 VGND VGND VPWR VPWR booth_b30_m16 sky130_fd_sc_hd__xor2_1
XU$$1360 t$5099 net1668 VGND VGND VPWR VPWR booth_b18_m60 sky130_fd_sc_hd__xor2_1
XU$$1371 net13 VGND VGND VPWR VPWR notblock$5105\[1\] sky130_fd_sc_hd__inv_1
XU$$1382 net1036 net629 net933 net902 VGND VGND VPWR VPWR t$5112 sky130_fd_sc_hd__a22o_1
XU$$1393 t$5117 net1485 VGND VGND VPWR VPWR booth_b20_m8 sky130_fd_sc_hd__xor2_1
XFILLER_50_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_119_1 c$3402 s$3405 s$3407 VGND VGND VPWR VPWR c$3874 s$3875 sky130_fd_sc_hd__fa_1
XFILLER_148_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1828_ clknet_leaf_234_clk booth_b10_m40 VGND VGND VPWR VPWR pp_row50_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1759_ clknet_leaf_23_clk booth_b42_m5 VGND VGND VPWR VPWR pp_row47_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_84_4 pp_row84_12 pp_row84_13 pp_row84_14 VGND VGND VPWR VPWR c$960 s$961
+ sky130_fd_sc_hd__fa_1
Xfanout901 net904 VGND VGND VPWR VPWR net901 sky130_fd_sc_hd__buf_6
Xfanout912 sel_1$5038 VGND VGND VPWR VPWR net912 sky130_fd_sc_hd__buf_6
Xfanout923 sel_1$4968 VGND VGND VPWR VPWR net923 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_77_3 pp_row77_12 pp_row77_13 pp_row77_14 VGND VGND VPWR VPWR c$840 s$841
+ sky130_fd_sc_hd__fa_1
XFILLER_89_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout934 net935 VGND VGND VPWR VPWR net934 sky130_fd_sc_hd__clkbuf_4
Xfanout945 net946 VGND VGND VPWR VPWR net945 sky130_fd_sc_hd__buf_4
Xdadda_fa_4_54_2 s$2273 s$2275 s$2277 VGND VGND VPWR VPWR c$3018 s$3019 sky130_fd_sc_hd__fa_1
Xfanout956 net957 VGND VGND VPWR VPWR net956 sky130_fd_sc_hd__buf_4
XTAP_4006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout967 net968 VGND VGND VPWR VPWR net967 sky130_fd_sc_hd__buf_4
XTAP_4017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout978 net980 VGND VGND VPWR VPWR net978 sky130_fd_sc_hd__buf_2
XFILLER_161_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout989 net92 VGND VGND VPWR VPWR net989 sky130_fd_sc_hd__clkbuf_8
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_47_1 c$2210 c$2212 s$2215 VGND VGND VPWR VPWR c$2974 s$2975 sky130_fd_sc_hd__fa_1
XFILLER_57_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_24_0 s$3495 c$3942 s$3945 VGND VGND VPWR VPWR c$4200 s$4201 sky130_fd_sc_hd__fa_1
XTAP_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_305 net421 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_316 net588 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_327 net680 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_338 net773 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_349 net874 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1093_1754 VGND VGND VPWR VPWR U$$1093_1754/HI net1754 sky130_fd_sc_hd__conb_1
XFILLER_122_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_0_72_2 pp_row72_6 pp_row72_7 pp_row72_8 VGND VGND VPWR VPWR c$176 s$177
+ sky130_fd_sc_hd__fa_1
XFILLER_114_1111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_0_65_1 pp_row65_3 pp_row65_4 pp_row65_5 VGND VGND VPWR VPWR c$98 s$99 sky130_fd_sc_hd__fa_1
XFILLER_114_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_42_0 s$253 c$1218 c$1220 VGND VGND VPWR VPWR c$2174 s$2175 sky130_fd_sc_hd__fa_1
XFILLER_49_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_58_0 pp_row58_0 pp_row58_1 pp_row58_2 VGND VGND VPWR VPWR c$24 s$25 sky130_fd_sc_hd__fa_1
XFILLER_48_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$590 final_adder.p_new$602 final_adder.p_new$594 VGND VGND VPWR VPWR
+ final_adder.p_new$718 sky130_fd_sc_hd__and2_1
XTAP_3872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$440 t$4630 net1245 VGND VGND VPWR VPWR booth_b6_m11 sky130_fd_sc_hd__xor2_1
XTAP_3883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$451 net1161 net431 net1149 net713 VGND VGND VPWR VPWR t$4636 sky130_fd_sc_hd__a22o_1
XTAP_3894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$462 t$4641 net1244 VGND VGND VPWR VPWR booth_b6_m22 sky130_fd_sc_hd__xor2_1
XFILLER_45_884 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$473 net1058 net429 net1050 net711 VGND VGND VPWR VPWR t$4647 sky130_fd_sc_hd__a22o_1
XU$$484 t$4652 net1250 VGND VGND VPWR VPWR booth_b6_m33 sky130_fd_sc_hd__xor2_1
XU$$495 net949 net427 net941 net709 VGND VGND VPWR VPWR t$4658 sky130_fd_sc_hd__a22o_1
X_0992_ clknet_leaf_116_clk booth_b58_m42 VGND VGND VPWR VPWR pp_row100_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_13_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_786 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1613_ clknet_leaf_239_clk booth_b24_m18 VGND VGND VPWR VPWR pp_row42_12 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_94_3 pp_row94_14 pp_row94_15 pp_row94_16 VGND VGND VPWR VPWR c$1860 s$1861
+ sky130_fd_sc_hd__fa_1
XFILLER_172_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_87_2 pp_row87_21 pp_row87_22 c$978 VGND VGND VPWR VPWR c$1774 s$1775 sky130_fd_sc_hd__fa_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1544_ clknet_leaf_16_clk booth_b30_m9 VGND VGND VPWR VPWR pp_row39_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_141_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_64_1 s$3075 s$3077 s$3079 VGND VGND VPWR VPWR c$3654 s$3655 sky130_fd_sc_hd__fa_1
XFILLER_5_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1475_ clknet_leaf_39_clk booth_b32_m4 VGND VGND VPWR VPWR pp_row36_16 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_57_0 c$3026 c$3028 c$3030 VGND VGND VPWR VPWR c$3624 s$3625 sky130_fd_sc_hd__fa_1
X_0426_ clknet_leaf_207_clk booth_b38_m39 VGND VGND VPWR VPWR pp_row77_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_189_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_56_8 c$10 s$13 s$15 VGND VGND VPWR VPWR c$472 s$473 sky130_fd_sc_hd__fa_1
X_0357_ clknet_leaf_196_clk booth_b26_m49 VGND VGND VPWR VPWR pp_row75_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_67_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$271_1780 VGND VGND VPWR VPWR U$$271_1780/HI net1780 sky130_fd_sc_hd__conb_1
XFILLER_36_840 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0288_ clknet_leaf_202_clk booth_b18_m55 VGND VGND VPWR VPWR pp_row73_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_42_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2027_ clknet_leaf_135_clk booth_b60_m48 VGND VGND VPWR VPWR pp_row108_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_36_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_103_0 pp_row103_0 pp_row103_1 pp_row103_2 VGND VGND VPWR VPWR c$1950 s$1951
+ sky130_fd_sc_hd__fa_1
XFILLER_51_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1190 net1730 net648 net1721 net921 VGND VGND VPWR VPWR t$5013 sky130_fd_sc_hd__a22o_1
XFILLER_148_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_82_1 pp_row82_3 pp_row82_4 pp_row82_5 VGND VGND VPWR VPWR c$924 s$925
+ sky130_fd_sc_hd__fa_1
XFILLER_137_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1707 net105 VGND VGND VPWR VPWR net1707 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout720 net723 VGND VGND VPWR VPWR net720 sky130_fd_sc_hd__clkbuf_4
Xfanout1718 net1719 VGND VGND VPWR VPWR net1718 sky130_fd_sc_hd__clkbuf_2
Xdadda_fa_1_75_0 pp_row75_6 pp_row75_7 pp_row75_8 VGND VGND VPWR VPWR c$798 s$799
+ sky130_fd_sc_hd__fa_1
XFILLER_172_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1729 net1732 VGND VGND VPWR VPWR net1729 sky130_fd_sc_hd__buf_4
Xfanout731 net732 VGND VGND VPWR VPWR net731 sky130_fd_sc_hd__buf_4
XFILLER_120_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout742 net744 VGND VGND VPWR VPWR net742 sky130_fd_sc_hd__buf_4
Xfanout753 net754 VGND VGND VPWR VPWR net753 sky130_fd_sc_hd__buf_4
Xfanout764 net765 VGND VGND VPWR VPWR net764 sky130_fd_sc_hd__buf_2
Xfanout775 net782 VGND VGND VPWR VPWR net775 sky130_fd_sc_hd__clkbuf_4
Xfanout786 net791 VGND VGND VPWR VPWR net786 sky130_fd_sc_hd__buf_4
Xfanout797 net798 VGND VGND VPWR VPWR net797 sky130_fd_sc_hd__buf_6
XFILLER_92_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3509 net951 net486 net943 net759 VGND VGND VPWR VPWR t$6198 sky130_fd_sc_hd__a22o_1
XTAP_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2808 net1027 net538 net1019 net811 VGND VGND VPWR VPWR t$5840 sky130_fd_sc_hd__a22o_1
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2819 t$5845 net1378 VGND VGND VPWR VPWR booth_b40_m36 sky130_fd_sc_hd__xor2_1
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_102 net568 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_113 net628 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_124 net674 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_135 net723 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_146 net773 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_157 net815 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_168 net895 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_179 net947 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1047 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_97_1 c$1882 c$1884 c$1886 VGND VGND VPWR VPWR c$2616 s$2617 sky130_fd_sc_hd__fa_1
XFILLER_155_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_74_0 c$3688 c$3690 s$3693 VGND VGND VPWR VPWR c$4044 s$4045 sky130_fd_sc_hd__fa_1
XFILLER_64_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1260_ clknet_leaf_109_clk booth_b54_m49 VGND VGND VPWR VPWR pp_row103_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_1_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0211_ clknet_leaf_184_clk net143 VGND VGND VPWR VPWR pp_row112_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1191_ clknet_leaf_59_clk booth_b8_m13 VGND VGND VPWR VPWR pp_row21_4 sky130_fd_sc_hd__dfxtp_1
Xinput8 a[16] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_4
XFILLER_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_119_0 pp_row119_0 pp_row119_1 pp_row119_2 VGND VGND VPWR VPWR c$3404 s$3405
+ sky130_fd_sc_hd__fa_1
XTAP_4370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$270 t$4542 net1392 VGND VGND VPWR VPWR booth_b2_m63 sky130_fd_sc_hd__xor2_1
XU$$281 t$4549 net1277 VGND VGND VPWR VPWR booth_b4_m0 sky130_fd_sc_hd__xor2_1
XFILLER_45_692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$292 net1564 net531 net1523 net804 VGND VGND VPWR VPWR t$4555 sky130_fd_sc_hd__a22o_1
XTAP_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0975_ clknet_leaf_116_clk booth_b60_m39 VGND VGND VPWR VPWR pp_row99_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_186_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1081 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$6 c$4162 s$4165 VGND VGND VPWR VPWR final_adder.$signal$14 final_adder.$signal$1096
+ sky130_fd_sc_hd__ha_1
XFILLER_134_907 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput301 net301 VGND VGND VPWR VPWR o[24] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_92_0 pp_row92_8 pp_row92_9 pp_row92_10 VGND VGND VPWR VPWR c$1830 s$1831
+ sky130_fd_sc_hd__fa_1
Xoutput312 net312 VGND VGND VPWR VPWR o[34] sky130_fd_sc_hd__buf_2
XU$$4391_1816 VGND VGND VPWR VPWR U$$4391_1816/HI net1816 sky130_fd_sc_hd__conb_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput323 net323 VGND VGND VPWR VPWR o[44] sky130_fd_sc_hd__buf_2
Xoutput334 net334 VGND VGND VPWR VPWR o[54] sky130_fd_sc_hd__buf_2
Xoutput345 net345 VGND VGND VPWR VPWR o[64] sky130_fd_sc_hd__buf_2
Xoutput356 net356 VGND VGND VPWR VPWR o[74] sky130_fd_sc_hd__buf_2
Xoutput367 net367 VGND VGND VPWR VPWR o[84] sky130_fd_sc_hd__buf_2
Xoutput378 net378 VGND VGND VPWR VPWR o[94] sky130_fd_sc_hd__buf_2
Xdadda_ha_4_118_2 pp_row118_6 pp_row118_7 VGND VGND VPWR VPWR c$3402 s$3403 sky130_fd_sc_hd__ha_1
XFILLER_114_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1527_ clknet_leaf_18_clk booth_b0_m39 VGND VGND VPWR VPWR pp_row39_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_113_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1458_ clknet_leaf_42_clk booth_b2_m34 VGND VGND VPWR VPWR pp_row36_1 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_61_6 c$40 c$42 c$44 VGND VGND VPWR VPWR c$558 s$559 sky130_fd_sc_hd__fa_1
XFILLER_171_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0409_ clknet_leaf_208_clk booth_b64_m12 VGND VGND VPWR VPWR pp_row76_27 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_54_5 pp_row54_20 pp_row54_21 pp_row54_22 VGND VGND VPWR VPWR c$430 s$431
+ sky130_fd_sc_hd__fa_1
X_1389_ clknet_leaf_45_clk booth_b32_m0 VGND VGND VPWR VPWR pp_row32_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_95_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_47_4 pp_row47_12 pp_row47_13 pp_row47_14 VGND VGND VPWR VPWR c$310 s$311
+ sky130_fd_sc_hd__fa_1
XFILLER_55_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_1148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_17_2 c$1980 s$1983 s$1985 VGND VGND VPWR VPWR c$2796 s$2797 sky130_fd_sc_hd__fa_1
XFILLER_35_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_91_0 s$3763 c$4076 s$4079 VGND VGND VPWR VPWR c$4334 s$4335 sky130_fd_sc_hd__fa_1
XFILLER_167_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1504 net1506 VGND VGND VPWR VPWR net1504 sky130_fd_sc_hd__buf_2
Xfanout1515 net1516 VGND VGND VPWR VPWR net1515 sky130_fd_sc_hd__buf_4
XFILLER_120_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1526 net125 VGND VGND VPWR VPWR net1526 sky130_fd_sc_hd__buf_4
Xfanout1537 net1538 VGND VGND VPWR VPWR net1537 sky130_fd_sc_hd__buf_2
XFILLER_120_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout550 sel_0$5737 VGND VGND VPWR VPWR net550 sky130_fd_sc_hd__buf_6
Xfanout1548 net1550 VGND VGND VPWR VPWR net1548 sky130_fd_sc_hd__buf_4
Xfanout1559 net121 VGND VGND VPWR VPWR net1559 sky130_fd_sc_hd__buf_8
XU$$4007 net1196 net451 net1177 net724 VGND VGND VPWR VPWR t$6453 sky130_fd_sc_hd__a22o_1
Xfanout561 net562 VGND VGND VPWR VPWR net561 sky130_fd_sc_hd__clkbuf_2
XU$$4018 t$6458 net1283 VGND VGND VPWR VPWR booth_b58_m19 sky130_fd_sc_hd__xor2_1
Xfanout572 sel_0$5527 VGND VGND VPWR VPWR net572 sky130_fd_sc_hd__buf_6
XFILLER_47_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout583 sel_0$5457 VGND VGND VPWR VPWR net583 sky130_fd_sc_hd__buf_6
XU$$4029 net1085 net454 net1077 net727 VGND VGND VPWR VPWR t$6464 sky130_fd_sc_hd__a22o_1
Xfanout594 net595 VGND VGND VPWR VPWR net594 sky130_fd_sc_hd__clkbuf_2
XFILLER_58_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3306 net1566 net497 net1525 net770 VGND VGND VPWR VPWR t$6095 sky130_fd_sc_hd__a22o_1
XU$$3317 t$6100 net1338 VGND VGND VPWR VPWR booth_b48_m11 sky130_fd_sc_hd__xor2_1
XU$$3328 net1163 net497 net1153 net770 VGND VGND VPWR VPWR t$6106 sky130_fd_sc_hd__a22o_1
XFILLER_73_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3339 t$6111 net1340 VGND VGND VPWR VPWR booth_b48_m22 sky130_fd_sc_hd__xor2_1
XU$$2605 net1397 VGND VGND VPWR VPWR notblock$5735\[2\] sky130_fd_sc_hd__inv_1
XU$$2616 t$5742 net1394 VGND VGND VPWR VPWR booth_b38_m3 sky130_fd_sc_hd__xor2_1
XU$$2627 net1504 net543 net1495 net816 VGND VGND VPWR VPWR t$5748 sky130_fd_sc_hd__a22o_1
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2638 t$5753 net1399 VGND VGND VPWR VPWR booth_b38_m14 sky130_fd_sc_hd__xor2_1
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1904 t$5377 net1463 VGND VGND VPWR VPWR booth_b26_m58 sky130_fd_sc_hd__xor2_1
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2649 net1134 net544 net1118 net817 VGND VGND VPWR VPWR t$5759 sky130_fd_sc_hd__a22o_1
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1915 net1532 net600 net1768 net873 VGND VGND VPWR VPWR t$5383 sky130_fd_sc_hd__a22o_1
XFILLER_61_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1926 net1227 net584 net1122 net857 VGND VGND VPWR VPWR t$5390 sky130_fd_sc_hd__a22o_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1937 t$5395 net1451 VGND VGND VPWR VPWR booth_b28_m6 sky130_fd_sc_hd__xor2_1
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1948 net1211 net585 net1201 net858 VGND VGND VPWR VPWR t$5401 sky130_fd_sc_hd__a22o_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1959 t$5406 net1449 VGND VGND VPWR VPWR booth_b28_m17 sky130_fd_sc_hd__xor2_1
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0760_ clknet_leaf_153_clk booth_b52_m37 VGND VGND VPWR VPWR pp_row89_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_127_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0691_ clknet_leaf_168_clk booth_b62_m24 VGND VGND VPWR VPWR pp_row86_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_143_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2430_ clknet_leaf_96_clk booth_b40_m27 VGND VGND VPWR VPWR pp_row67_20 sky130_fd_sc_hd__dfxtp_1
XFILLER_143_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2361_ clknet_leaf_75_clk booth_b50_m15 VGND VGND VPWR VPWR pp_row65_25 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_71_5 s$737 s$739 s$741 VGND VGND VPWR VPWR c$1588 s$1589 sky130_fd_sc_hd__fa_1
XFILLER_155_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1312_ clknet_leaf_246_clk booth_b28_m0 VGND VGND VPWR VPWR pp_row28_14 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_64_4 s$605 s$607 s$609 VGND VGND VPWR VPWR c$1502 s$1503 sky130_fd_sc_hd__fa_2
X_2292_ clknet_leaf_212_clk booth_b58_m5 VGND VGND VPWR VPWR pp_row63_29 sky130_fd_sc_hd__dfxtp_1
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1243_ clknet_leaf_15_clk booth_b24_m0 VGND VGND VPWR VPWR pp_row24_12 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_57_3 c$472 s$475 s$477 VGND VGND VPWR VPWR c$1416 s$1417 sky130_fd_sc_hd__fa_1
XFILLER_2_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$11 t$4412 net1573 VGND VGND VPWR VPWR booth_b0_m2 sky130_fd_sc_hd__xor2_1
XU$$22 net1515 net446 net1508 net688 VGND VGND VPWR VPWR t$4418 sky130_fd_sc_hd__a22o_1
XU$$33 t$4423 net1574 VGND VGND VPWR VPWR booth_b0_m13 sky130_fd_sc_hd__xor2_1
X_1174_ clknet_leaf_46_clk booth_b2_m18 VGND VGND VPWR VPWR pp_row20_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_38_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$44 net1143 net448 net1133 net690 VGND VGND VPWR VPWR t$4429 sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_27_1 s$2853 s$2855 s$2857 VGND VGND VPWR VPWR c$3506 s$3507 sky130_fd_sc_hd__fa_2
XU$$55 t$4434 net1569 VGND VGND VPWR VPWR booth_b0_m24 sky130_fd_sc_hd__xor2_1
XU$$3840 notblock$6365\[2\] net52 net1302 t$6366 notblock$6365\[0\] VGND VGND VPWR
+ VPWR sel_0$6367 sky130_fd_sc_hd__a32o_4
XU$$66 net1039 net442 net1023 net684 VGND VGND VPWR VPWR t$4440 sky130_fd_sc_hd__a22o_1
XFILLER_37_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3851 t$6373 net1291 VGND VGND VPWR VPWR booth_b56_m4 sky130_fd_sc_hd__xor2_1
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3862 net1501 net467 net1226 net740 VGND VGND VPWR VPWR t$6379 sky130_fd_sc_hd__a22o_1
XU$$3873 t$6384 net1295 VGND VGND VPWR VPWR booth_b56_m15 sky130_fd_sc_hd__xor2_1
XU$$77 t$4445 net1575 VGND VGND VPWR VPWR booth_b0_m35 sky130_fd_sc_hd__xor2_1
XU$$88 net924 net444 net1745 net686 VGND VGND VPWR VPWR t$4451 sky130_fd_sc_hd__a22o_1
XU$$99 t$4456 net1570 VGND VGND VPWR VPWR booth_b0_m46 sky130_fd_sc_hd__xor2_1
XU$$3884 net1119 net460 net1111 net733 VGND VGND VPWR VPWR t$6390 sky130_fd_sc_hd__a22o_1
XU$$3895 t$6395 net1294 VGND VGND VPWR VPWR booth_b56_m26 sky130_fd_sc_hd__xor2_1
XFILLER_80_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_13 pp_row55_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_24 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_35 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_46 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_57 net243 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_68 net425 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_79 net487 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0958_ clknet_leaf_114_clk booth_b62_m36 VGND VGND VPWR VPWR pp_row98_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_174_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_101_1 s$3297 s$3299 s$3301 VGND VGND VPWR VPWR c$3802 s$3803 sky130_fd_sc_hd__fa_1
XFILLER_161_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_929 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0889_ clknet_leaf_100_clk booth_b44_m51 VGND VGND VPWR VPWR pp_row95_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_133_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_ha_1_39_2 pp_row39_6 pp_row39_7 VGND VGND VPWR VPWR c$226 s$227 sky130_fd_sc_hd__ha_1
Xdadda_fa_1_52_2 pp_row52_8 pp_row52_9 pp_row52_10 VGND VGND VPWR VPWR c$388 s$389
+ sky130_fd_sc_hd__fa_1
XFILLER_29_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_45_1 pp_row45_3 pp_row45_4 pp_row45_5 VGND VGND VPWR VPWR c$278 s$279
+ sky130_fd_sc_hd__fa_1
XFILLER_55_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_22_0 s$1051 c$2006 c$2008 VGND VGND VPWR VPWR c$2822 s$2823 sky130_fd_sc_hd__fa_1
Xdadda_fa_1_38_0 pp_row38_0 pp_row38_1 pp_row38_2 VGND VGND VPWR VPWR c$216 s$217
+ sky130_fd_sc_hd__fa_1
XFILLER_12_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1005 final_adder.$signal$1134 final_adder.g_new$951 VGND VGND VPWR
+ VPWR net323 sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$1016 final_adder.$signal$113 final_adder.g_new$1062 VGND VGND VPWR
+ VPWR net335 sky130_fd_sc_hd__xor2_2
XFILLER_11_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$1027 final_adder.$signal$1156 final_adder.g_new$1025 VGND VGND VPWR
+ VPWR net347 sky130_fd_sc_hd__xor2_2
XFILLER_109_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1038 final_adder.$signal$1167 final_adder.g_new$1051 VGND VGND VPWR
+ VPWR net359 sky130_fd_sc_hd__xor2_2
XFILLER_137_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1049 final_adder.$signal$1178 final_adder.g_new$1003 VGND VGND VPWR
+ VPWR net371 sky130_fd_sc_hd__xor2_2
XFILLER_152_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_74_3 s$1619 s$1621 s$1623 VGND VGND VPWR VPWR c$2436 s$2437 sky130_fd_sc_hd__fa_1
XFILLER_105_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1301 net1303 VGND VGND VPWR VPWR net1301 sky130_fd_sc_hd__buf_6
Xfanout1312 net1315 VGND VGND VPWR VPWR net1312 sky130_fd_sc_hd__buf_6
Xdadda_fa_3_67_2 c$1528 s$1531 s$1533 VGND VGND VPWR VPWR c$2378 s$2379 sky130_fd_sc_hd__fa_1
XFILLER_61_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1323 net1328 VGND VGND VPWR VPWR net1323 sky130_fd_sc_hd__buf_4
XFILLER_78_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1334 net1336 VGND VGND VPWR VPWR net1334 sky130_fd_sc_hd__buf_6
Xfanout1345 net1346 VGND VGND VPWR VPWR net1345 sky130_fd_sc_hd__buf_6
Xfanout1356 net42 VGND VGND VPWR VPWR net1356 sky130_fd_sc_hd__buf_6
XFILLER_47_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1367 net1368 VGND VGND VPWR VPWR net1367 sky130_fd_sc_hd__buf_6
XFILLER_66_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1378 net1380 VGND VGND VPWR VPWR net1378 sky130_fd_sc_hd__buf_6
XFILLER_94_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout391 net392 VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__buf_6
Xfanout1389 net1391 VGND VGND VPWR VPWR net1389 sky130_fd_sc_hd__buf_6
Xdadda_fa_6_37_0 c$3540 c$3542 s$3545 VGND VGND VPWR VPWR c$3970 s$3971 sky130_fd_sc_hd__fa_1
XU$$3103 t$5990 net1359 VGND VGND VPWR VPWR booth_b44_m41 sky130_fd_sc_hd__xor2_1
XU$$3114 net1708 net515 net1700 net788 VGND VGND VPWR VPWR t$5996 sky130_fd_sc_hd__a22o_1
XU$$3125 t$6001 net1364 VGND VGND VPWR VPWR booth_b44_m52 sky130_fd_sc_hd__xor2_1
XU$$3136 net1602 net516 net1593 net789 VGND VGND VPWR VPWR t$6007 sky130_fd_sc_hd__a22o_1
XFILLER_59_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2402 t$5632 net1424 VGND VGND VPWR VPWR booth_b34_m33 sky130_fd_sc_hd__xor2_1
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3147 t$6012 net1365 VGND VGND VPWR VPWR booth_b44_m63 sky130_fd_sc_hd__xor2_1
XU$$2413 net949 net562 net941 net835 VGND VGND VPWR VPWR t$5638 sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_194_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_194_clk
+ sky130_fd_sc_hd__clkbuf_16
XU$$3158 t$6019 net1349 VGND VGND VPWR VPWR booth_b46_m0 sky130_fd_sc_hd__xor2_1
XU$$3169 net1566 net505 net1526 net778 VGND VGND VPWR VPWR t$6025 sky130_fd_sc_hd__a22o_1
XU$$2424 t$5643 net1426 VGND VGND VPWR VPWR booth_b34_m44 sky130_fd_sc_hd__xor2_1
XFILLER_59_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2435 net1680 net566 net1655 net839 VGND VGND VPWR VPWR t$5649 sky130_fd_sc_hd__a22o_1
XFILLER_34_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1701 t$5274 net1468 VGND VGND VPWR VPWR booth_b24_m25 sky130_fd_sc_hd__xor2_1
XU$$2446 t$5654 net1425 VGND VGND VPWR VPWR booth_b34_m55 sky130_fd_sc_hd__xor2_1
XU$$2457 net1557 net568 net1550 net841 VGND VGND VPWR VPWR t$5660 sky130_fd_sc_hd__a22o_1
XU$$1712 net1026 net606 net1018 net879 VGND VGND VPWR VPWR t$5280 sky130_fd_sc_hd__a22o_1
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2468 net1408 VGND VGND VPWR VPWR notblock$5665\[2\] sky130_fd_sc_hd__inv_1
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1723 t$5285 net1470 VGND VGND VPWR VPWR booth_b24_m36 sky130_fd_sc_hd__xor2_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1734 net1749 net606 net1741 net879 VGND VGND VPWR VPWR t$5291 sky130_fd_sc_hd__a22o_1
XFILLER_185_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2479 t$5672 net1404 VGND VGND VPWR VPWR booth_b36_m3 sky130_fd_sc_hd__xor2_1
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1745 t$5296 net1473 VGND VGND VPWR VPWR booth_b24_m47 sky130_fd_sc_hd__xor2_1
XFILLER_15_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1756 net1639 net609 net1631 net882 VGND VGND VPWR VPWR t$5302 sky130_fd_sc_hd__a22o_1
X_1930_ clknet_leaf_62_clk booth_b26_m27 VGND VGND VPWR VPWR pp_row53_13 sky130_fd_sc_hd__dfxtp_1
XU$$1767 t$5307 net1471 VGND VGND VPWR VPWR booth_b24_m58 sky130_fd_sc_hd__xor2_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1778 net1529 net609 net1766 net882 VGND VGND VPWR VPWR t$5313 sky130_fd_sc_hd__a22o_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1789 net1227 net593 net1122 net866 VGND VGND VPWR VPWR t$5320 sky130_fd_sc_hd__a22o_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1861_ clknet_leaf_133_clk booth_b54_m53 VGND VGND VPWR VPWR pp_row107_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_187_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0812_ clknet_leaf_93_clk booth_b62_m29 VGND VGND VPWR VPWR pp_row91_18 sky130_fd_sc_hd__dfxtp_1
Xinput11 a[19] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_4
XFILLER_35_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput22 a[29] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
X_1792_ clknet_leaf_232_clk net199 VGND VGND VPWR VPWR pp_row48_26 sky130_fd_sc_hd__dfxtp_1
Xinput33 a[39] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_6
XFILLER_128_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput44 a[49] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_1
Xinput55 a[59] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_4
X_0743_ clknet_leaf_184_clk net243 VGND VGND VPWR VPWR pp_row88_22 sky130_fd_sc_hd__dfxtp_1
Xinput66 b[10] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__buf_6
XFILLER_143_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput77 b[20] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_6
Xinput88 b[30] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_2
XFILLER_192_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput99 b[40] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__dlymetal6s2s_1
X_0674_ clknet_leaf_170_clk booth_b32_m54 VGND VGND VPWR VPWR pp_row86_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_192_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2413_ clknet_leaf_84_clk booth_b10_m57 VGND VGND VPWR VPWR pp_row67_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2344_ clknet_leaf_87_clk booth_b20_m45 VGND VGND VPWR VPWR pp_row65_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_69_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_62_1 c$550 c$552 c$554 VGND VGND VPWR VPWR c$1472 s$1473 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$408 final_adder.p_new$414 final_adder.p_new$410 VGND VGND VPWR VPWR
+ final_adder.p_new$536 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$419 final_adder.p_new$420 final_adder.g_new$425 final_adder.g_new$421
+ VGND VGND VPWR VPWR final_adder.g_new$547 sky130_fd_sc_hd__a21o_1
X_2275_ clknet_leaf_217_clk booth_b28_m35 VGND VGND VPWR VPWR pp_row63_14 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_55_0 s$11 c$420 c$422 VGND VGND VPWR VPWR c$1386 s$1387 sky130_fd_sc_hd__fa_1
XFILLER_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1226_ clknet_leaf_48_clk booth_b20_m3 VGND VGND VPWR VPWR pp_row23_10 sky130_fd_sc_hd__dfxtp_1
XU$$4360 t$6632 net1260 VGND VGND VPWR VPWR booth_b62_m53 sky130_fd_sc_hd__xor2_1
XU$$4371 net1588 net419 net1579 net701 VGND VGND VPWR VPWR t$6638 sky130_fd_sc_hd__a22o_1
XU$$4382 t$6643 net1255 VGND VGND VPWR VPWR booth_b62_m64 sky130_fd_sc_hd__xor2_1
XU$$4393 t$6650 net1817 VGND VGND VPWR VPWR booth_b64_m1 sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_185_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_185_clk
+ sky130_fd_sc_hd__clkbuf_16
X_1157_ clknet_leaf_15_clk net1664 VGND VGND VPWR VPWR pp_row18_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_77_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3670 net1660 net482 net1652 net755 VGND VGND VPWR VPWR t$6280 sky130_fd_sc_hd__a22o_1
XFILLER_25_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3681 t$6285 net1327 VGND VGND VPWR VPWR booth_b52_m56 sky130_fd_sc_hd__xor2_1
XU$$3692 net1549 net483 net1541 net756 VGND VGND VPWR VPWR t$6291 sky130_fd_sc_hd__a22o_1
X_1088_ clknet_leaf_58_clk booth_b8_m4 VGND VGND VPWR VPWR pp_row12_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_80_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_9_0 pp_row9_2 pp_row9_3 pp_row9_4 VGND VGND VPWR VPWR c$3432 s$3433 sky130_fd_sc_hd__fa_1
XU$$2980 t$5927 net1371 VGND VGND VPWR VPWR booth_b42_m48 sky130_fd_sc_hd__xor2_1
XU$$2991 net1637 net524 net1627 net797 VGND VGND VPWR VPWR t$5933 sky130_fd_sc_hd__a22o_1
XFILLER_179_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_84_2 s$2513 s$2515 s$2517 VGND VGND VPWR VPWR c$3198 s$3199 sky130_fd_sc_hd__fa_1
XFILLER_164_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_77_1 c$2450 c$2452 s$2455 VGND VGND VPWR VPWR c$3154 s$3155 sky130_fd_sc_hd__fa_1
XFILLER_106_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_54_0 s$3615 c$4002 s$4005 VGND VGND VPWR VPWR c$4260 s$4261 sky130_fd_sc_hd__fa_1
XFILLER_115_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$920 final_adder.$signal$1172 final_adder.g_new$1009 final_adder.$signal$166
+ VGND VGND VPWR VPWR final_adder.g_new$1048 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$931 final_adder.$signal$1150 final_adder.g_new$935 final_adder.$signal$122
+ VGND VGND VPWR VPWR final_adder.g_new$1059 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$942 final_adder.$signal$1128 final_adder.g_new$957 final_adder.$signal$78
+ VGND VGND VPWR VPWR final_adder.g_new$1070 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$953 final_adder.$signal$1106 final_adder.g_new$747 final_adder.$signal$34
+ VGND VGND VPWR VPWR final_adder.g_new$1081 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$964 final_adder.$signal$1093 final_adder.g_new$1088 VGND VGND VPWR
+ VPWR net318 sky130_fd_sc_hd__xor2_1
XU$$803 net1615 net407 net1607 net673 VGND VGND VPWR VPWR t$4815 sky130_fd_sc_hd__a22o_1
XU$$814 t$4820 net1417 VGND VGND VPWR VPWR booth_b10_m61 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$975 final_adder.$signal$1104 final_adder.g_new$749 VGND VGND VPWR
+ VPWR net290 sky130_fd_sc_hd__xor2_2
XU$$825 net1316 notblock$4825\[1\] VGND VGND VPWR VPWR t$4826 sky130_fd_sc_hd__and2_1
XFILLER_16_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$986 final_adder.$signal$1115 final_adder.g_new$1077 VGND VGND VPWR
+ VPWR net302 sky130_fd_sc_hd__xor2_2
Xclkbuf_leaf_176_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_176_clk
+ sky130_fd_sc_hd__clkbuf_16
XU$$836 net933 net394 net1672 net660 VGND VGND VPWR VPWR t$4833 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$997 final_adder.$signal$1126 final_adder.g_new$959 VGND VGND VPWR
+ VPWR net314 sky130_fd_sc_hd__xor2_2
XU$$847 t$4838 net1313 VGND VGND VPWR VPWR booth_b12_m9 sky130_fd_sc_hd__xor2_1
XU$$858 net1173 net393 net1164 net659 VGND VGND VPWR VPWR t$4844 sky130_fd_sc_hd__a22o_1
XU$$1008 t$4920 net1187 VGND VGND VPWR VPWR booth_b14_m21 sky130_fd_sc_hd__xor2_1
XFILLER_44_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$869 t$4849 net1314 VGND VGND VPWR VPWR booth_b12_m20 sky130_fd_sc_hd__xor2_1
XFILLER_189_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1019 net1063 net386 net1055 net652 VGND VGND VPWR VPWR t$4926 sky130_fd_sc_hd__a22o_1
XFILLER_71_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1057 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_100_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_100_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_98_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_72_0 s$761 c$1578 c$1580 VGND VGND VPWR VPWR c$2414 s$2415 sky130_fd_sc_hd__fa_1
XFILLER_98_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1000 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0390_ clknet_leaf_196_clk booth_b28_m48 VGND VGND VPWR VPWR pp_row76_9 sky130_fd_sc_hd__dfxtp_1
Xfanout1120 net1121 VGND VGND VPWR VPWR net1120 sky130_fd_sc_hd__buf_6
Xfanout1131 net1132 VGND VGND VPWR VPWR net1131 sky130_fd_sc_hd__buf_2
Xfanout1142 net74 VGND VGND VPWR VPWR net1142 sky130_fd_sc_hd__clkbuf_4
Xfanout1153 net1154 VGND VGND VPWR VPWR net1153 sky130_fd_sc_hd__clkbuf_8
XFILLER_93_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1164 net1167 VGND VGND VPWR VPWR net1164 sky130_fd_sc_hd__buf_4
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1175 net1176 VGND VGND VPWR VPWR net1175 sky130_fd_sc_hd__buf_4
Xfanout1186 net1187 VGND VGND VPWR VPWR net1186 sky130_fd_sc_hd__clkbuf_8
X_2060_ clknet_leaf_184_clk net138 VGND VGND VPWR VPWR pp_row108_12 sky130_fd_sc_hd__dfxtp_2
Xfanout1197 net69 VGND VGND VPWR VPWR net1197 sky130_fd_sc_hd__clkbuf_4
XFILLER_19_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1011_ clknet_leaf_115_clk booth_b60_m41 VGND VGND VPWR VPWR pp_row101_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_47_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_167_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_167_clk
+ sky130_fd_sc_hd__clkbuf_16
XU$$2210 net1560 net569 net1519 net842 VGND VGND VPWR VPWR t$5535 sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_101_0 s$1941 c$2638 c$2640 VGND VGND VPWR VPWR c$3296 s$3297 sky130_fd_sc_hd__fa_1
XU$$2221 t$5540 net1430 VGND VGND VPWR VPWR booth_b32_m11 sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_34_5 pp_row34_17 pp_row34_18 pp_row34_19 VGND VGND VPWR VPWR c$1144 s$1145
+ sky130_fd_sc_hd__fa_1
XU$$2232 net1158 net569 net1148 net842 VGND VGND VPWR VPWR t$5546 sky130_fd_sc_hd__a22o_1
XU$$2243 t$5551 net1433 VGND VGND VPWR VPWR booth_b32_m22 sky130_fd_sc_hd__xor2_1
XFILLER_179_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2254 net1056 net570 net1048 net843 VGND VGND VPWR VPWR t$5557 sky130_fd_sc_hd__a22o_1
XU$$2265 t$5562 net1433 VGND VGND VPWR VPWR booth_b32_m33 sky130_fd_sc_hd__xor2_1
XU$$1520 t$5182 net1475 VGND VGND VPWR VPWR booth_b22_m3 sky130_fd_sc_hd__xor2_1
XU$$1531 net1503 net611 net1494 net884 VGND VGND VPWR VPWR t$5188 sky130_fd_sc_hd__a22o_1
XU$$2276 net951 net573 net942 net846 VGND VGND VPWR VPWR t$5568 sky130_fd_sc_hd__a22o_1
XU$$2287 t$5573 net1434 VGND VGND VPWR VPWR booth_b32_m44 sky130_fd_sc_hd__xor2_1
XFILLER_37_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1542 t$5193 net1478 VGND VGND VPWR VPWR booth_b22_m14 sky130_fd_sc_hd__xor2_1
XU$$1553 net1132 net610 net1116 net883 VGND VGND VPWR VPWR t$5199 sky130_fd_sc_hd__a22o_1
XU$$2298 net1680 net573 net1655 net846 VGND VGND VPWR VPWR t$5579 sky130_fd_sc_hd__a22o_1
XFILLER_16_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1564 t$5204 net1477 VGND VGND VPWR VPWR booth_b22_m25 sky130_fd_sc_hd__xor2_1
XFILLER_97_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1575 net1025 net614 net1017 net887 VGND VGND VPWR VPWR t$5210 sky130_fd_sc_hd__a22o_1
XFILLER_72_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1586 t$5215 net1484 VGND VGND VPWR VPWR booth_b22_m36 sky130_fd_sc_hd__xor2_1
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1913_ clknet_leaf_31_clk net1320 VGND VGND VPWR VPWR pp_row52_27 sky130_fd_sc_hd__dfxtp_1
XU$$1597 net1749 net618 net1741 net891 VGND VGND VPWR VPWR t$5221 sky130_fd_sc_hd__a22o_1
XFILLER_187_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1844_ clknet_leaf_71_clk booth_b38_m12 VGND VGND VPWR VPWR pp_row50_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_175_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_94_1 s$3255 s$3257 s$3259 VGND VGND VPWR VPWR c$3774 s$3775 sky130_fd_sc_hd__fa_1
XFILLER_147_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1775_ clknet_leaf_239_clk booth_b20_m28 VGND VGND VPWR VPWR pp_row48_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_129_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_87_0 c$3206 c$3208 c$3210 VGND VGND VPWR VPWR c$3744 s$3745 sky130_fd_sc_hd__fa_1
X_0726_ clknet_leaf_161_clk booth_b34_m54 VGND VGND VPWR VPWR pp_row88_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_171_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0657_ clknet_leaf_178_clk booth_b46_m39 VGND VGND VPWR VPWR pp_row85_13 sky130_fd_sc_hd__dfxtp_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_79_7 pp_row79_21 pp_row79_22 pp_row79_23 VGND VGND VPWR VPWR c$884 s$885
+ sky130_fd_sc_hd__fa_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0588_ clknet_leaf_120_clk booth_b62_m54 VGND VGND VPWR VPWR pp_row116_6 sky130_fd_sc_hd__dfxtp_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2327_ clknet_leaf_127_clk notsign$6084 VGND VGND VPWR VPWR pp_row111_0 sky130_fd_sc_hd__dfxtp_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$205 final_adder.$signal$105 final_adder.$signal$102 final_adder.$signal$104
+ VGND VGND VPWR VPWR final_adder.g_new$333 sky130_fd_sc_hd__a21o_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$216 final_adder.$signal$1128 final_adder.$signal$1129 VGND VGND VPWR
+ VPWR final_adder.p_new$344 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$227 final_adder.$signal$1119 final_adder.$signal$58 final_adder.$signal$60
+ VGND VGND VPWR VPWR final_adder.g_new$355 sky130_fd_sc_hd__a21o_1
XTAP_3509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$238 final_adder.$signal$1106 final_adder.$signal$1107 VGND VGND VPWR
+ VPWR final_adder.p_new$366 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$249 final_adder.$signal$1097 final_adder.$signal$14 final_adder.$signal$16
+ VGND VGND VPWR VPWR final_adder.g_new$377 sky130_fd_sc_hd__a21o_1
X_2258_ clknet_leaf_231_clk net215 VGND VGND VPWR VPWR pp_row62_33 sky130_fd_sc_hd__dfxtp_1
XFILLER_38_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1209_ clknet_leaf_49_clk booth_b16_m6 VGND VGND VPWR VPWR pp_row22_8 sky130_fd_sc_hd__dfxtp_1
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_158_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_158_clk
+ sky130_fd_sc_hd__clkbuf_16
XU$$4190 net971 net438 net962 net720 VGND VGND VPWR VPWR t$6546 sky130_fd_sc_hd__a22o_1
X_2189_ clknet_leaf_227_clk booth_b4_m57 VGND VGND VPWR VPWR pp_row61_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_168_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4509_1875 VGND VGND VPWR VPWR U$$4509_1875/HI net1875 sky130_fd_sc_hd__conb_1
XFILLER_26_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_790 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_103_2 c$1942 c$1944 c$1946 VGND VGND VPWR VPWR c$2666 s$2667 sky130_fd_sc_hd__fa_1
XFILLER_134_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_1088 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput201 c[4] VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkbuf_1
XFILLER_68_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput212 c[5] VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput223 c[6] VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__clkbuf_1
Xinput234 c[7] VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput245 c[8] VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_0_67_5 pp_row67_15 pp_row67_16 pp_row67_17 VGND VGND VPWR VPWR c$130 s$131
+ sky130_fd_sc_hd__fa_2
Xinput256 c[9] VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_117_0 c$3860 c$3862 s$3865 VGND VGND VPWR VPWR c$4130 s$4131 sky130_fd_sc_hd__fa_1
XFILLER_25_1080 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$750 final_adder.p_new$798 final_adder.p_new$766 VGND VGND VPWR VPWR
+ final_adder.p_new$878 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$761 final_adder.p_new$776 final_adder.g_new$809 final_adder.g_new$777
+ VGND VGND VPWR VPWR final_adder.g_new$889 sky130_fd_sc_hd__a21o_1
XU$$600 net1097 net410 net1088 net676 VGND VGND VPWR VPWR t$4712 sky130_fd_sc_hd__a22o_1
XFILLER_57_871 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$611 t$4717 net1239 VGND VGND VPWR VPWR booth_b8_m28 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$772 final_adder.p_new$820 final_adder.p_new$788 VGND VGND VPWR VPWR
+ final_adder.p_new$900 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$783 final_adder.p_new$798 final_adder.g_new$831 final_adder.g_new$799
+ VGND VGND VPWR VPWR final_adder.g_new$911 sky130_fd_sc_hd__a21o_1
XU$$622 net990 net409 net982 net675 VGND VGND VPWR VPWR t$4723 sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_149_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_149_clk
+ sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_3_37_3 s$1175 s$1177 s$1179 VGND VGND VPWR VPWR c$2140 s$2141 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$794 final_adder.p_new$842 final_adder.p_new$810 VGND VGND VPWR VPWR
+ final_adder.p_new$922 sky130_fd_sc_hd__and2_1
XU$$633 t$4728 net1235 VGND VGND VPWR VPWR booth_b8_m39 sky130_fd_sc_hd__xor2_1
XU$$644 net1725 net417 net1716 net683 VGND VGND VPWR VPWR t$4734 sky130_fd_sc_hd__a22o_1
XU$$655 t$4739 net1242 VGND VGND VPWR VPWR booth_b8_m50 sky130_fd_sc_hd__xor2_1
XU$$666 net1612 net411 net1604 net677 VGND VGND VPWR VPWR t$4745 sky130_fd_sc_hd__a22o_1
XU$$677 t$4750 net1242 VGND VGND VPWR VPWR booth_b8_m61 sky130_fd_sc_hd__xor2_1
XFILLER_140_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$688 net1417 notblock$4755\[1\] VGND VGND VPWR VPWR t$4756 sky130_fd_sc_hd__and2_1
XFILLER_72_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$699 net933 net406 net1672 net672 VGND VGND VPWR VPWR t$4763 sky130_fd_sc_hd__a22o_1
XFILLER_108_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_98_0_1908 VGND VGND VPWR VPWR net1908 dadda_fa_2_98_0_1908/LO sky130_fd_sc_hd__conb_1
X_1560_ clknet_leaf_7_clk booth_b18_m22 VGND VGND VPWR VPWR pp_row40_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0511_ clknet_leaf_126_clk booth_b64_m51 VGND VGND VPWR VPWR pp_row115_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_154_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1491_ clknet_leaf_18_clk booth_b20_m17 VGND VGND VPWR VPWR pp_row37_10 sky130_fd_sc_hd__dfxtp_1
X_0442_ clknet_leaf_151_clk booth_b14_m64 VGND VGND VPWR VPWR pp_row78_1 sky130_fd_sc_hd__dfxtp_1
X_0373_ clknet_leaf_204_clk booth_b56_m19 VGND VGND VPWR VPWR pp_row75_23 sky130_fd_sc_hd__dfxtp_1
XFILLER_95_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2112_ clknet_leaf_86_clk booth_b58_m0 VGND VGND VPWR VPWR pp_row58_29 sky130_fd_sc_hd__dfxtp_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2043_ clknet_leaf_85_clk booth_b56_m0 VGND VGND VPWR VPWR pp_row56_28 sky130_fd_sc_hd__dfxtp_1
XFILLER_35_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_32_2 pp_row32_6 pp_row32_7 pp_row32_8 VGND VGND VPWR VPWR c$1114 s$1115
+ sky130_fd_sc_hd__fa_1
XU$$2040 net1597 net590 net1588 net863 VGND VGND VPWR VPWR t$5447 sky130_fd_sc_hd__a22o_1
XU$$2051 t$5452 net1455 VGND VGND VPWR VPWR booth_b28_m63 sky130_fd_sc_hd__xor2_1
XU$$2062 t$5459 net1439 VGND VGND VPWR VPWR booth_b30_m0 sky130_fd_sc_hd__xor2_1
XU$$2073 net1565 net581 net1524 net854 VGND VGND VPWR VPWR t$5465 sky130_fd_sc_hd__a22o_1
XU$$2084 t$5470 net1439 VGND VGND VPWR VPWR booth_b30_m11 sky130_fd_sc_hd__xor2_1
XU$$2095 net1156 net576 net1148 net849 VGND VGND VPWR VPWR t$5476 sky130_fd_sc_hd__a22o_1
XU$$1350 t$5094 net1669 VGND VGND VPWR VPWR booth_b18_m55 sky130_fd_sc_hd__xor2_1
XU$$1361 net1552 net641 net1546 net914 VGND VGND VPWR VPWR t$5100 sky130_fd_sc_hd__a22o_1
XU$$1372 net1491 VGND VGND VPWR VPWR notblock$5105\[2\] sky130_fd_sc_hd__inv_1
XU$$1383 t$5112 net1487 VGND VGND VPWR VPWR booth_b20_m3 sky130_fd_sc_hd__xor2_1
XFILLER_188_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1394 net1503 net627 net1494 net900 VGND VGND VPWR VPWR t$5118 sky130_fd_sc_hd__a22o_1
XFILLER_149_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1827_ clknet_leaf_135_clk booth_b48_m59 VGND VGND VPWR VPWR pp_row107_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_117_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1758_ clknet_leaf_219_clk booth_b40_m7 VGND VGND VPWR VPWR pp_row47_20 sky130_fd_sc_hd__dfxtp_1
XFILLER_144_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0709_ clknet_leaf_168_clk booth_b50_m37 VGND VGND VPWR VPWR pp_row87_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_143_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_84_5 pp_row84_15 pp_row84_16 pp_row84_17 VGND VGND VPWR VPWR c$962 s$963
+ sky130_fd_sc_hd__fa_1
X_1689_ clknet_leaf_18_clk booth_b16_m29 VGND VGND VPWR VPWR pp_row45_8 sky130_fd_sc_hd__dfxtp_1
Xfanout902 net903 VGND VGND VPWR VPWR net902 sky130_fd_sc_hd__clkbuf_8
Xfanout913 net915 VGND VGND VPWR VPWR net913 sky130_fd_sc_hd__buf_4
Xfanout924 net925 VGND VGND VPWR VPWR net924 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_77_4 pp_row77_15 pp_row77_16 pp_row77_17 VGND VGND VPWR VPWR c$842 s$843
+ sky130_fd_sc_hd__fa_1
Xfanout935 net98 VGND VGND VPWR VPWR net935 sky130_fd_sc_hd__buf_6
Xfanout946 net947 VGND VGND VPWR VPWR net946 sky130_fd_sc_hd__buf_4
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout957 net960 VGND VGND VPWR VPWR net957 sky130_fd_sc_hd__buf_6
XTAP_4007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout968 net94 VGND VGND VPWR VPWR net968 sky130_fd_sc_hd__buf_6
XFILLER_135_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout979 net980 VGND VGND VPWR VPWR net979 sky130_fd_sc_hd__buf_6
XTAP_4029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_47_2 s$2217 s$2219 s$2221 VGND VGND VPWR VPWR c$2976 s$2977 sky130_fd_sc_hd__fa_1
XFILLER_86_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_306 net445 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_17_0 s$3467 c$3928 s$3931 VGND VGND VPWR VPWR c$4186 s$4187 sky130_fd_sc_hd__fa_2
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_317 net588 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_328 net680 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_339 net775 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$90 c$4330 s$4333 VGND VGND VPWR VPWR final_adder.$signal$182 final_adder.$signal$1180
+ sky130_fd_sc_hd__ha_2
XFILLER_13_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_857 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_0_59_3 pp_row59_9 pp_row59_10 VGND VGND VPWR VPWR c$38 s$39 sky130_fd_sc_hd__ha_1
XFILLER_110_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1044 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_0_65_2 pp_row65_6 pp_row65_7 pp_row65_8 VGND VGND VPWR VPWR c$100 s$101
+ sky130_fd_sc_hd__fa_1
XFILLER_92_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_42_1 c$1222 c$1224 c$1226 VGND VGND VPWR VPWR c$2176 s$2177 sky130_fd_sc_hd__fa_1
Xdadda_fa_0_58_1 pp_row58_3 pp_row58_4 pp_row58_5 VGND VGND VPWR VPWR c$26 s$27 sky130_fd_sc_hd__fa_1
XTAP_3840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_35_0 s$207 c$1134 c$1136 VGND VGND VPWR VPWR c$2118 s$2119 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$580 final_adder.p_new$592 final_adder.p_new$584 VGND VGND VPWR VPWR
+ final_adder.p_new$708 sky130_fd_sc_hd__and2_1
XTAP_3862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$591 final_adder.p_new$594 final_adder.g_new$603 final_adder.g_new$595
+ VGND VGND VPWR VPWR final_adder.g_new$719 sky130_fd_sc_hd__a21o_1
XU$$430 t$4625 net1248 VGND VGND VPWR VPWR booth_b6_m6 sky130_fd_sc_hd__xor2_1
XTAP_3873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$441 net1211 net431 net1203 net713 VGND VGND VPWR VPWR t$4631 sky130_fd_sc_hd__a22o_1
XFILLER_151_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$452 t$4636 net1250 VGND VGND VPWR VPWR booth_b6_m17 sky130_fd_sc_hd__xor2_1
XTAP_3895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$463 net1097 net426 net1088 net708 VGND VGND VPWR VPWR t$4642 sky130_fd_sc_hd__a22o_1
XFILLER_44_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$474 t$4647 net1248 VGND VGND VPWR VPWR booth_b6_m28 sky130_fd_sc_hd__xor2_1
XU$$485 net990 net428 net986 net710 VGND VGND VPWR VPWR t$4653 sky130_fd_sc_hd__a22o_1
XFILLER_17_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$496 t$4658 net1253 VGND VGND VPWR VPWR booth_b6_m39 sky130_fd_sc_hd__xor2_1
XFILLER_60_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2052_1770 VGND VGND VPWR VPWR U$$2052_1770/HI net1770 sky130_fd_sc_hd__conb_1
X_0991_ clknet_leaf_118_clk booth_b56_m44 VGND VGND VPWR VPWR pp_row100_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_160_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1612_ clknet_leaf_239_clk booth_b22_m20 VGND VGND VPWR VPWR pp_row42_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_145_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_94_4 pp_row94_17 pp_row94_18 pp_row94_19 VGND VGND VPWR VPWR c$1862 s$1863
+ sky130_fd_sc_hd__fa_1
XFILLER_114_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1543_ clknet_leaf_16_clk booth_b28_m11 VGND VGND VPWR VPWR pp_row39_14 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_87_3 c$980 c$982 c$984 VGND VGND VPWR VPWR c$1776 s$1777 sky130_fd_sc_hd__fa_1
XFILLER_113_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1474_ clknet_leaf_39_clk booth_b30_m6 VGND VGND VPWR VPWR pp_row36_15 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_57_1 s$3033 s$3035 s$3037 VGND VGND VPWR VPWR c$3626 s$3627 sky130_fd_sc_hd__fa_1
XFILLER_101_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0425_ clknet_leaf_207_clk booth_b36_m41 VGND VGND VPWR VPWR pp_row77_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_80_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0356_ clknet_leaf_196_clk booth_b24_m51 VGND VGND VPWR VPWR pp_row75_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_27_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0287_ clknet_leaf_202_clk booth_b16_m57 VGND VGND VPWR VPWR pp_row73_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_36_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2026_ clknet_leaf_35_clk booth_b26_m30 VGND VGND VPWR VPWR pp_row56_13 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_103_1 pp_row103_3 pp_row103_4 pp_row103_5 VGND VGND VPWR VPWR c$1952 s$1953
+ sky130_fd_sc_hd__fa_2
Xdadda_fa_1_92_0_1902 VGND VGND VPWR VPWR net1902 dadda_fa_1_92_0_1902/LO sky130_fd_sc_hd__conb_1
XFILLER_23_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1180 net955 net645 net944 net918 VGND VGND VPWR VPWR t$5008 sky130_fd_sc_hd__a22o_1
XU$$1191 t$5013 net1008 VGND VGND VPWR VPWR booth_b16_m44 sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_124_0 net1914 pp_row124_1 pp_row124_2 VGND VGND VPWR VPWR c$3892 s$3893
+ sky130_fd_sc_hd__fa_1
XFILLER_148_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_82_2 pp_row82_6 pp_row82_7 pp_row82_8 VGND VGND VPWR VPWR c$926 s$927
+ sky130_fd_sc_hd__fa_1
XFILLER_132_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_719 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1708 net1710 VGND VGND VPWR VPWR net1708 sky130_fd_sc_hd__buf_4
XFILLER_172_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout710 net715 VGND VGND VPWR VPWR net710 sky130_fd_sc_hd__buf_6
XFILLER_137_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1719 net104 VGND VGND VPWR VPWR net1719 sky130_fd_sc_hd__buf_6
Xfanout721 net722 VGND VGND VPWR VPWR net721 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_75_1 pp_row75_9 pp_row75_10 pp_row75_11 VGND VGND VPWR VPWR c$800 s$801
+ sky130_fd_sc_hd__fa_1
Xfanout732 sel_1$6438 VGND VGND VPWR VPWR net732 sky130_fd_sc_hd__clkbuf_4
Xfanout743 net744 VGND VGND VPWR VPWR net743 sky130_fd_sc_hd__clkbuf_4
Xfanout754 sel_1$6228 VGND VGND VPWR VPWR net754 sky130_fd_sc_hd__buf_4
Xdadda_fa_4_52_0 s$1361 c$2246 c$2248 VGND VGND VPWR VPWR c$3002 s$3003 sky130_fd_sc_hd__fa_1
Xdadda_fa_1_68_0 pp_row68_17 pp_row68_18 pp_row68_19 VGND VGND VPWR VPWR c$672 s$673
+ sky130_fd_sc_hd__fa_1
Xfanout765 sel_1$6158 VGND VGND VPWR VPWR net765 sky130_fd_sc_hd__clkbuf_8
Xdadda_ha_2_102_3 pp_row102_9 pp_row102_10 VGND VGND VPWR VPWR c$1948 s$1949 sky130_fd_sc_hd__ha_1
Xfanout776 net782 VGND VGND VPWR VPWR net776 sky130_fd_sc_hd__buf_4
Xfanout787 net790 VGND VGND VPWR VPWR net787 sky130_fd_sc_hd__buf_4
XFILLER_74_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout798 net799 VGND VGND VPWR VPWR net798 sky130_fd_sc_hd__buf_4
XFILLER_74_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2809 t$5840 net1380 VGND VGND VPWR VPWR booth_b40_m31 sky130_fd_sc_hd__xor2_1
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_103 net568 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_114 net631 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_125 net683 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_136 net728 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_147 net790 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_158 net815 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_169 net895 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_80_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_80_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_97_2 c$1888 s$1891 s$1893 VGND VGND VPWR VPWR c$2618 s$2619 sky130_fd_sc_hd__fa_1
XFILLER_170_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_67_0 c$3660 c$3662 s$3665 VGND VGND VPWR VPWR c$4030 s$4031 sky130_fd_sc_hd__fa_1
XFILLER_123_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_70_0 net1892 pp_row70_1 pp_row70_2 VGND VGND VPWR VPWR c$154 s$155 sky130_fd_sc_hd__fa_1
XFILLER_1_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0210_ clknet_leaf_154_clk booth_b60_m10 VGND VGND VPWR VPWR pp_row70_28 sky130_fd_sc_hd__dfxtp_1
X_1190_ clknet_leaf_59_clk booth_b6_m15 VGND VGND VPWR VPWR pp_row21_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput9 a[17] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_4
XTAP_4360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_119_1 pp_row119_3 pp_row119_4 pp_row119_5 VGND VGND VPWR VPWR c$3406 s$3407
+ sky130_fd_sc_hd__fa_1
XTAP_4371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_5_6_1 pp_row6_3 pp_row6_4 VGND VGND VPWR VPWR c$3422 s$3423 sky130_fd_sc_hd__ha_1
XTAP_3670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$260 t$4537 net1388 VGND VGND VPWR VPWR booth_b2_m58 sky130_fd_sc_hd__xor2_1
XU$$271 net1531 net626 net1780 net899 VGND VGND VPWR VPWR t$4543 sky130_fd_sc_hd__a22o_1
XU$$282 net1232 net531 net1127 net804 VGND VGND VPWR VPWR t$4550 sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_71_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_71_clk sky130_fd_sc_hd__clkbuf_16
XU$$293 t$4555 net1277 VGND VGND VPWR VPWR booth_b4_m6 sky130_fd_sc_hd__xor2_1
XTAP_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0974_ clknet_leaf_116_clk booth_b58_m41 VGND VGND VPWR VPWR pp_row99_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_192_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$7 c$4164 s$4167 VGND VGND VPWR VPWR final_adder.$signal$16 final_adder.$signal$1097
+ sky130_fd_sc_hd__ha_1
XFILLER_134_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput302 net302 VGND VGND VPWR VPWR o[25] sky130_fd_sc_hd__buf_2
XFILLER_161_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_92_1 pp_row92_11 pp_row92_12 pp_row92_13 VGND VGND VPWR VPWR c$1832 s$1833
+ sky130_fd_sc_hd__fa_1
Xoutput313 net313 VGND VGND VPWR VPWR o[35] sky130_fd_sc_hd__buf_2
XFILLER_133_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput324 net324 VGND VGND VPWR VPWR o[45] sky130_fd_sc_hd__buf_2
XFILLER_99_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput335 net335 VGND VGND VPWR VPWR o[55] sky130_fd_sc_hd__buf_2
Xoutput346 net346 VGND VGND VPWR VPWR o[65] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_85_0 pp_row85_18 pp_row85_19 pp_row85_20 VGND VGND VPWR VPWR c$1746 s$1747
+ sky130_fd_sc_hd__fa_1
Xoutput357 net357 VGND VGND VPWR VPWR o[75] sky130_fd_sc_hd__buf_2
Xoutput368 net368 VGND VGND VPWR VPWR o[85] sky130_fd_sc_hd__buf_2
X_1526_ clknet_leaf_236_clk net188 VGND VGND VPWR VPWR pp_row38_21 sky130_fd_sc_hd__dfxtp_1
Xoutput379 net379 VGND VGND VPWR VPWR o[95] sky130_fd_sc_hd__buf_2
XFILLER_113_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_1_48_7 pp_row48_21 pp_row48_22 VGND VGND VPWR VPWR c$330 s$331 sky130_fd_sc_hd__ha_1
XFILLER_99_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1457_ clknet_leaf_41_clk booth_b0_m36 VGND VGND VPWR VPWR pp_row36_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_61_7 c$46 c$48 s$51 VGND VGND VPWR VPWR c$560 s$561 sky130_fd_sc_hd__fa_1
XFILLER_45_1083 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0408_ clknet_leaf_206_clk booth_b62_m14 VGND VGND VPWR VPWR pp_row76_26 sky130_fd_sc_hd__dfxtp_1
XFILLER_142_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1388_ clknet_leaf_45_clk booth_b30_m2 VGND VGND VPWR VPWR pp_row32_15 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_54_6 pp_row54_23 pp_row54_24 pp_row54_25 VGND VGND VPWR VPWR c$432 s$433
+ sky130_fd_sc_hd__fa_1
XFILLER_83_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0339_ clknet_leaf_226_clk booth_b52_m22 VGND VGND VPWR VPWR pp_row74_22 sky130_fd_sc_hd__dfxtp_1
XFILLER_55_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_47_5 pp_row47_15 pp_row47_16 pp_row47_17 VGND VGND VPWR VPWR c$312 s$313
+ sky130_fd_sc_hd__fa_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_6_0 s$3423 c$3906 s$3909 VGND VGND VPWR VPWR c$4164 s$4165 sky130_fd_sc_hd__fa_1
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2009_ clknet_leaf_76_clk booth_b52_m3 VGND VGND VPWR VPWR pp_row55_26 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_62_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_62_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_23_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_84_0 s$3735 c$4062 s$4065 VGND VGND VPWR VPWR c$4320 s$4321 sky130_fd_sc_hd__fa_2
XFILLER_100_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1505 net1506 VGND VGND VPWR VPWR net1505 sky130_fd_sc_hd__buf_4
Xfanout1516 net1518 VGND VGND VPWR VPWR net1516 sky130_fd_sc_hd__buf_4
Xfanout1527 net1530 VGND VGND VPWR VPWR net1527 sky130_fd_sc_hd__buf_4
Xfanout540 net541 VGND VGND VPWR VPWR net540 sky130_fd_sc_hd__buf_4
Xfanout1538 net123 VGND VGND VPWR VPWR net1538 sky130_fd_sc_hd__buf_6
Xfanout551 net553 VGND VGND VPWR VPWR net551 sky130_fd_sc_hd__buf_4
XFILLER_116_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1549 net1550 VGND VGND VPWR VPWR net1549 sky130_fd_sc_hd__clkbuf_4
Xfanout562 net568 VGND VGND VPWR VPWR net562 sky130_fd_sc_hd__clkbuf_8
XU$$4008 t$6453 net1282 VGND VGND VPWR VPWR booth_b58_m14 sky130_fd_sc_hd__xor2_1
Xfanout573 net574 VGND VGND VPWR VPWR net573 sky130_fd_sc_hd__buf_4
XU$$4019 net1135 net451 net1119 net724 VGND VGND VPWR VPWR t$6459 sky130_fd_sc_hd__a22o_1
Xfanout584 net586 VGND VGND VPWR VPWR net584 sky130_fd_sc_hd__buf_4
Xfanout595 net601 VGND VGND VPWR VPWR net595 sky130_fd_sc_hd__buf_2
XFILLER_111_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3307 t$6095 net1343 VGND VGND VPWR VPWR booth_b48_m6 sky130_fd_sc_hd__xor2_1
XFILLER_101_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3318 net1214 net493 net1202 net766 VGND VGND VPWR VPWR t$6101 sky130_fd_sc_hd__a22o_1
XU$$3329 t$6106 net1343 VGND VGND VPWR VPWR booth_b48_m17 sky130_fd_sc_hd__xor2_1
XFILLER_100_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2606 net1397 notblock$5735\[1\] VGND VGND VPWR VPWR t$5736 sky130_fd_sc_hd__and2_1
XU$$2617 net932 net543 net1671 net816 VGND VGND VPWR VPWR t$5743 sky130_fd_sc_hd__a22o_1
XFILLER_74_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2628 t$5748 net1394 VGND VGND VPWR VPWR booth_b38_m9 sky130_fd_sc_hd__xor2_1
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2639 net1180 net549 net1171 net822 VGND VGND VPWR VPWR t$5754 sky130_fd_sc_hd__a22o_1
XU$$1905 net1588 net599 net1579 net872 VGND VGND VPWR VPWR t$5378 sky130_fd_sc_hd__a22o_1
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1916 t$5383 net1465 VGND VGND VPWR VPWR booth_b26_m64 sky130_fd_sc_hd__xor2_1
XU$$1927 t$5390 net1448 VGND VGND VPWR VPWR booth_b28_m1 sky130_fd_sc_hd__xor2_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1938 net1524 net587 net1516 net860 VGND VGND VPWR VPWR t$5396 sky130_fd_sc_hd__a22o_1
XFILLER_26_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_53_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_53_clk sky130_fd_sc_hd__clkbuf_16
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1949 t$5401 net1449 VGND VGND VPWR VPWR booth_b28_m12 sky130_fd_sc_hd__xor2_1
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0690_ clknet_leaf_168_clk booth_b60_m26 VGND VGND VPWR VPWR pp_row86_20 sky130_fd_sc_hd__dfxtp_1
XFILLER_127_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2360_ clknet_leaf_74_clk booth_b48_m17 VGND VGND VPWR VPWR pp_row65_24 sky130_fd_sc_hd__dfxtp_1
XFILLER_69_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1311_ clknet_leaf_3_clk booth_b26_m2 VGND VGND VPWR VPWR pp_row28_13 sky130_fd_sc_hd__dfxtp_1
X_2291_ clknet_leaf_214_clk booth_b56_m7 VGND VGND VPWR VPWR pp_row63_28 sky130_fd_sc_hd__dfxtp_1
XFILLER_116_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_64_5 s$611 s$613 s$615 VGND VGND VPWR VPWR c$1504 s$1505 sky130_fd_sc_hd__fa_2
X_1242_ clknet_leaf_15_clk booth_b22_m2 VGND VGND VPWR VPWR pp_row24_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_38_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_57_4 s$479 s$481 s$483 VGND VGND VPWR VPWR c$1418 s$1419 sky130_fd_sc_hd__fa_2
XFILLER_37_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$12 net1035 net446 net937 net688 VGND VGND VPWR VPWR t$4413 sky130_fd_sc_hd__a22o_1
XFILLER_38_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1173_ clknet_leaf_46_clk booth_b0_m20 VGND VGND VPWR VPWR pp_row20_0 sky130_fd_sc_hd__dfxtp_1
XU$$23 t$4418 net1573 VGND VGND VPWR VPWR booth_b0_m8 sky130_fd_sc_hd__xor2_1
XU$$34 net1194 net448 net1175 net690 VGND VGND VPWR VPWR t$4424 sky130_fd_sc_hd__a22o_1
XU$$3830 t$6361 net1306 VGND VGND VPWR VPWR booth_b54_m62 sky130_fd_sc_hd__xor2_1
XU$$3841 net52 net1302 VGND VGND VPWR VPWR sel_1$6368 sky130_fd_sc_hd__xor2_4
XU$$45 t$4429 net1575 VGND VGND VPWR VPWR booth_b0_m19 sky130_fd_sc_hd__xor2_1
XTAP_4190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$56 net1080 net443 net1071 net685 VGND VGND VPWR VPWR t$4435 sky130_fd_sc_hd__a22o_1
XU$$67 t$4440 net1568 VGND VGND VPWR VPWR booth_b0_m30 sky130_fd_sc_hd__xor2_1
XU$$3852 net1674 net461 net1563 net734 VGND VGND VPWR VPWR t$6374 sky130_fd_sc_hd__a22o_1
XU$$3863 t$6379 net1296 VGND VGND VPWR VPWR booth_b56_m10 sky130_fd_sc_hd__xor2_1
XU$$78 net977 net448 net969 net690 VGND VGND VPWR VPWR t$4446 sky130_fd_sc_hd__a22o_1
XU$$3874 net1168 net460 net1159 net733 VGND VGND VPWR VPWR t$6385 sky130_fd_sc_hd__a22o_1
XU$$89 t$4451 net1570 VGND VGND VPWR VPWR booth_b0_m41 sky130_fd_sc_hd__xor2_1
XFILLER_52_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3885 t$6390 net1294 VGND VGND VPWR VPWR booth_b56_m21 sky130_fd_sc_hd__xor2_1
XFILLER_18_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3896 net1069 net463 net1061 net736 VGND VGND VPWR VPWR t$6396 sky130_fd_sc_hd__a22o_1
XFILLER_80_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_44_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_44_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_75_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_14 s$4323 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_25 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_36 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_47 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_58 net283 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_69 net433 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0957_ clknet_leaf_114_clk booth_b60_m38 VGND VGND VPWR VPWR pp_row98_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_119_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0888_ clknet_leaf_130_clk booth_b60_m60 VGND VGND VPWR VPWR pp_row120_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_134_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1509_ clknet_leaf_17_clk booth_b10_m28 VGND VGND VPWR VPWR pp_row38_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_130_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2489_ clknet_leaf_90_clk booth_b20_m49 VGND VGND VPWR VPWR pp_row69_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_102_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_52_3 pp_row52_11 pp_row52_12 pp_row52_13 VGND VGND VPWR VPWR c$390 s$391
+ sky130_fd_sc_hd__fa_1
XFILLER_46_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_45_2 pp_row45_6 pp_row45_7 pp_row45_8 VGND VGND VPWR VPWR c$280 s$281
+ sky130_fd_sc_hd__fa_1
Xdadda_fa_4_22_1 c$2010 c$2012 s$2015 VGND VGND VPWR VPWR c$2824 s$2825 sky130_fd_sc_hd__fa_1
XFILLER_70_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_38_1 pp_row38_3 pp_row38_4 pp_row38_5 VGND VGND VPWR VPWR c$218 s$219
+ sky130_fd_sc_hd__fa_1
XFILLER_71_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_15_0 pp_row15_2 pp_row15_3 pp_row15_4 VGND VGND VPWR VPWR c$2780 s$2781
+ sky130_fd_sc_hd__fa_1
XFILLER_102_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_35_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_23_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1006 final_adder.$signal$1135 final_adder.g_new$1067 VGND VGND VPWR
+ VPWR net324 sky130_fd_sc_hd__xor2_2
XFILLER_183_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1017 final_adder.$signal$1146 final_adder.g_new$939 VGND VGND VPWR
+ VPWR net336 sky130_fd_sc_hd__xor2_1
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$1028 final_adder.$signal$1157 final_adder.g_new$1056 VGND VGND VPWR
+ VPWR net348 sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$1039 final_adder.$signal$1168 final_adder.g_new$1013 VGND VGND VPWR
+ VPWR net360 sky130_fd_sc_hd__xor2_2
XFILLER_178_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_760 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1302 net1303 VGND VGND VPWR VPWR net1302 sky130_fd_sc_hd__clkbuf_4
Xfanout1313 net1315 VGND VGND VPWR VPWR net1313 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_3_67_3 s$1535 s$1537 s$1539 VGND VGND VPWR VPWR c$2380 s$2381 sky130_fd_sc_hd__fa_1
Xfanout1324 net1325 VGND VGND VPWR VPWR net1324 sky130_fd_sc_hd__buf_6
Xfanout1335 net1336 VGND VGND VPWR VPWR net1335 sky130_fd_sc_hd__buf_6
XFILLER_78_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3285_1790 VGND VGND VPWR VPWR U$$3285_1790/HI net1790 sky130_fd_sc_hd__conb_1
Xfanout1346 net1347 VGND VGND VPWR VPWR net1346 sky130_fd_sc_hd__buf_6
Xfanout1357 net1366 VGND VGND VPWR VPWR net1357 sky130_fd_sc_hd__buf_6
XFILLER_8_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1368 net38 VGND VGND VPWR VPWR net1368 sky130_fd_sc_hd__buf_6
XFILLER_47_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1379 net1380 VGND VGND VPWR VPWR net1379 sky130_fd_sc_hd__buf_4
Xfanout392 sel_0$4897 VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__buf_8
XFILLER_87_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3104 net1747 net512 net1739 net785 VGND VGND VPWR VPWR t$5991 sky130_fd_sc_hd__a22o_1
XU$$3115 t$5996 net1364 VGND VGND VPWR VPWR booth_b44_m47 sky130_fd_sc_hd__xor2_1
XFILLER_86_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3126 net1644 net515 net1635 net788 VGND VGND VPWR VPWR t$6002 sky130_fd_sc_hd__a22o_1
XU$$3137 t$6007 net1365 VGND VGND VPWR VPWR booth_b44_m58 sky130_fd_sc_hd__xor2_1
XU$$2403 net996 net567 net988 net840 VGND VGND VPWR VPWR t$5633 sky130_fd_sc_hd__a22o_1
XU$$3148 net1532 net513 net1788 net786 VGND VGND VPWR VPWR t$6013 sky130_fd_sc_hd__a22o_1
XU$$2414 t$5638 net1422 VGND VGND VPWR VPWR booth_b34_m39 sky130_fd_sc_hd__xor2_1
XU$$3159 net1229 net501 net1125 net774 VGND VGND VPWR VPWR t$6020 sky130_fd_sc_hd__a22o_1
XU$$2425 net1722 net565 net1713 net838 VGND VGND VPWR VPWR t$5644 sky130_fd_sc_hd__a22o_1
XU$$2436 t$5649 net1426 VGND VGND VPWR VPWR booth_b34_m50 sky130_fd_sc_hd__xor2_1
XFILLER_61_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1702 net1073 net604 net1064 net877 VGND VGND VPWR VPWR t$5275 sky130_fd_sc_hd__a22o_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2447 net1615 net567 net1607 net840 VGND VGND VPWR VPWR t$5655 sky130_fd_sc_hd__a22o_1
XU$$2458 t$5660 net1428 VGND VGND VPWR VPWR booth_b34_m61 sky130_fd_sc_hd__xor2_1
XU$$1713 t$5280 net1470 VGND VGND VPWR VPWR booth_b24_m31 sky130_fd_sc_hd__xor2_1
XU$$1724 net965 net604 net957 net877 VGND VGND VPWR VPWR t$5286 sky130_fd_sc_hd__a22o_1
XU$$2469 net1408 notblock$5665\[1\] VGND VGND VPWR VPWR t$5666 sky130_fd_sc_hd__and2_1
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_26_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_16
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1735 t$5291 net1470 VGND VGND VPWR VPWR booth_b24_m42 sky130_fd_sc_hd__xor2_1
XU$$1746 net1697 net607 net1689 net880 VGND VGND VPWR VPWR t$5297 sky130_fd_sc_hd__a22o_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1757 t$5302 net1474 VGND VGND VPWR VPWR booth_b24_m53 sky130_fd_sc_hd__xor2_1
XU$$4461_1851 VGND VGND VPWR VPWR U$$4461_1851/HI net1851 sky130_fd_sc_hd__conb_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1768 net1588 net608 net1579 net881 VGND VGND VPWR VPWR t$5308 sky130_fd_sc_hd__a22o_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1779 t$5313 net1474 VGND VGND VPWR VPWR booth_b24_m64 sky130_fd_sc_hd__xor2_1
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1860_ clknet_leaf_80_clk booth_b12_m39 VGND VGND VPWR VPWR pp_row51_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_30_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0811_ clknet_leaf_97_clk booth_b60_m31 VGND VGND VPWR VPWR pp_row91_17 sky130_fd_sc_hd__dfxtp_1
Xinput12 a[1] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_2
X_1791_ clknet_leaf_222_clk net1338 VGND VGND VPWR VPWR pp_row48_25 sky130_fd_sc_hd__dfxtp_1
XFILLER_156_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput23 a[2] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_4
Xinput34 a[3] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_2
Xinput45 a[4] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_4
X_0742_ clknet_leaf_166_clk booth_b64_m24 VGND VGND VPWR VPWR pp_row88_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_156_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput56 a[5] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_2
Xinput67 b[11] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_4
Xinput78 b[21] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__buf_4
Xinput89 b[31] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0673_ clknet_leaf_175_clk booth_b30_m56 VGND VGND VPWR VPWR pp_row86_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_192_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2412_ clknet_leaf_84_clk booth_b8_m59 VGND VGND VPWR VPWR pp_row67_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_170_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2343_ clknet_leaf_87_clk booth_b18_m47 VGND VGND VPWR VPWR pp_row65_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_111_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_62_2 c$556 c$558 c$560 VGND VGND VPWR VPWR c$1474 s$1475 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$409 final_adder.p_new$410 final_adder.g_new$415 final_adder.g_new$411
+ VGND VGND VPWR VPWR final_adder.g_new$537 sky130_fd_sc_hd__a21o_1
X_2274_ clknet_leaf_209_clk booth_b26_m37 VGND VGND VPWR VPWR pp_row63_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_42_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_55_1 c$424 c$426 c$428 VGND VGND VPWR VPWR c$1388 s$1389 sky130_fd_sc_hd__fa_2
XFILLER_81_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1225_ clknet_leaf_48_clk booth_b18_m5 VGND VGND VPWR VPWR pp_row23_9 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_32_0 c$2876 c$2878 c$2880 VGND VGND VPWR VPWR c$3524 s$3525 sky130_fd_sc_hd__fa_1
XU$$4350 t$6627 net1256 VGND VGND VPWR VPWR booth_b62_m48 sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_48_0 pp_row48_23 pp_row48_24 pp_row48_25 VGND VGND VPWR VPWR c$1302 s$1303
+ sky130_fd_sc_hd__fa_1
XU$$4361 net1636 net424 net1625 net706 VGND VGND VPWR VPWR t$6633 sky130_fd_sc_hd__a22o_1
XU$$4372 t$6638 net1255 VGND VGND VPWR VPWR booth_b62_m59 sky130_fd_sc_hd__xor2_1
XFILLER_77_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4383 net1257 VGND VGND VPWR VPWR notsign$6644 sky130_fd_sc_hd__inv_1
X_1156_ clknet_leaf_15_clk booth_b18_m0 VGND VGND VPWR VPWR pp_row18_9 sky130_fd_sc_hd__dfxtp_1
XU$$4394 net76 sel_0$6647 net1038 net698 VGND VGND VPWR VPWR t$6651 sky130_fd_sc_hd__a22o_1
XU$$3660 net1717 sel_0$6227 net1708 sel_1$6228 VGND VGND VPWR VPWR t$6275 sky130_fd_sc_hd__a22o_1
XU$$3671 t$6280 net1326 VGND VGND VPWR VPWR booth_b52_m51 sky130_fd_sc_hd__xor2_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3682 net1608 net483 net1600 net756 VGND VGND VPWR VPWR t$6286 sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_17_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_16
XU$$3693 t$6291 net1327 VGND VGND VPWR VPWR booth_b52_m62 sky130_fd_sc_hd__xor2_1
X_1087_ clknet_leaf_58_clk booth_b6_m6 VGND VGND VPWR VPWR pp_row12_3 sky130_fd_sc_hd__dfxtp_1
XU$$2970 t$5922 net1369 VGND VGND VPWR VPWR booth_b42_m43 sky130_fd_sc_hd__xor2_1
XFILLER_179_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_9_1 pp_row9_5 c$2750 s$2753 VGND VGND VPWR VPWR c$3434 s$3435 sky130_fd_sc_hd__fa_1
XU$$2981 net1692 net525 net1685 net798 VGND VGND VPWR VPWR t$5928 sky130_fd_sc_hd__a22o_1
XU$$2992 t$5933 net1373 VGND VGND VPWR VPWR booth_b42_m54 sky130_fd_sc_hd__xor2_1
XFILLER_119_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1989_ clknet_leaf_81_clk booth_b16_m39 VGND VGND VPWR VPWR pp_row55_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_193_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_77_2 s$2457 s$2459 s$2461 VGND VGND VPWR VPWR c$3156 s$3157 sky130_fd_sc_hd__fa_1
XFILLER_115_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_47_0 s$3587 c$3988 s$3991 VGND VGND VPWR VPWR c$4246 s$4247 sky130_fd_sc_hd__fa_2
XFILLER_75_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$910 final_adder.$signal$1192 final_adder.g_new$989 final_adder.$signal$206
+ VGND VGND VPWR VPWR final_adder.g_new$1038 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$921 final_adder.$signal$1170 final_adder.g_new$1011 final_adder.$signal$162
+ VGND VGND VPWR VPWR final_adder.g_new$1049 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$932 final_adder.$signal$1148 final_adder.g_new$937 final_adder.$signal$118
+ VGND VGND VPWR VPWR final_adder.g_new$1060 sky130_fd_sc_hd__a21o_1
XFILLER_21_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_50_0 pp_row50_0 pp_row50_1 pp_row50_2 VGND VGND VPWR VPWR c$348 s$349
+ sky130_fd_sc_hd__fa_2
XFILLER_56_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$943 final_adder.$signal$1126 final_adder.g_new$959 final_adder.$signal$74
+ VGND VGND VPWR VPWR final_adder.g_new$1071 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$954 final_adder.$signal$1104 final_adder.g_new$749 final_adder.$signal$30
+ VGND VGND VPWR VPWR final_adder.g_new$1082 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$965 final_adder.$signal$1094 final_adder.g_new$509 VGND VGND VPWR
+ VPWR net329 sky130_fd_sc_hd__xor2_2
XFILLER_21_1137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$804 t$4815 net1419 VGND VGND VPWR VPWR booth_b10_m56 sky130_fd_sc_hd__xor2_1
XU$$815 net1543 net403 net1535 net669 VGND VGND VPWR VPWR t$4821 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$976 final_adder.$signal$1105 final_adder.g_new$1082 VGND VGND VPWR
+ VPWR net291 sky130_fd_sc_hd__xor2_2
XU$$826 notblock$4825\[2\] net4 net1417 t$4826 notblock$4825\[0\] VGND VGND VPWR VPWR
+ sel_0$4827 sky130_fd_sc_hd__a32o_1
Xfinal_adder.U$$987 final_adder.$signal$1116 final_adder.g_new$857 VGND VGND VPWR
+ VPWR net303 sky130_fd_sc_hd__xor2_2
XFILLER_16_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$837 t$4833 net1310 VGND VGND VPWR VPWR booth_b12_m4 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$998 final_adder.$signal$1127 final_adder.g_new$1071 VGND VGND VPWR
+ VPWR net315 sky130_fd_sc_hd__xor2_2
XU$$848 net1496 net396 net1221 net662 VGND VGND VPWR VPWR t$4839 sky130_fd_sc_hd__a22o_1
XU$$859 t$4844 net1310 VGND VGND VPWR VPWR booth_b12_m15 sky130_fd_sc_hd__xor2_1
XU$$1009 net1108 net388 net1100 net654 VGND VGND VPWR VPWR t$4921 sky130_fd_sc_hd__a22o_1
XFILLER_44_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_936 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_885 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4491_1866 VGND VGND VPWR VPWR U$$4491_1866/HI net1866 sky130_fd_sc_hd__conb_1
XFILLER_180_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_72_1 c$1582 c$1584 c$1586 VGND VGND VPWR VPWR c$2416 s$2417 sky130_fd_sc_hd__fa_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1110 net78 VGND VGND VPWR VPWR net1110 sky130_fd_sc_hd__buf_6
Xdadda_fa_3_65_0 s$635 c$1494 c$1496 VGND VGND VPWR VPWR c$2358 s$2359 sky130_fd_sc_hd__fa_1
Xfanout1121 net77 VGND VGND VPWR VPWR net1121 sky130_fd_sc_hd__buf_4
Xfanout1132 net75 VGND VGND VPWR VPWR net1132 sky130_fd_sc_hd__buf_6
XFILLER_78_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1143 net1145 VGND VGND VPWR VPWR net1143 sky130_fd_sc_hd__buf_4
Xfanout1154 net73 VGND VGND VPWR VPWR net1154 sky130_fd_sc_hd__buf_4
Xfanout1165 net1167 VGND VGND VPWR VPWR net1165 sky130_fd_sc_hd__buf_2
XFILLER_120_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1176 net1182 VGND VGND VPWR VPWR net1176 sky130_fd_sc_hd__clkbuf_4
XFILLER_19_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1187 net7 VGND VGND VPWR VPWR net1187 sky130_fd_sc_hd__buf_6
XFILLER_187_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1198 net1200 VGND VGND VPWR VPWR net1198 sky130_fd_sc_hd__buf_6
X_1010_ clknet_leaf_129_clk booth_b60_m62 VGND VGND VPWR VPWR pp_row122_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_47_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2200 net1230 net571 net1126 net844 VGND VGND VPWR VPWR t$5530 sky130_fd_sc_hd__a22o_1
XU$$2211 t$5535 net1430 VGND VGND VPWR VPWR booth_b32_m6 sky130_fd_sc_hd__xor2_1
XFILLER_47_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_101_1 c$2642 c$2644 s$2647 VGND VGND VPWR VPWR c$3298 s$3299 sky130_fd_sc_hd__fa_1
XFILLER_74_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2222 net1212 net569 net1204 net842 VGND VGND VPWR VPWR t$5541 sky130_fd_sc_hd__a22o_1
XFILLER_62_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2233 t$5546 net1431 VGND VGND VPWR VPWR booth_b32_m17 sky130_fd_sc_hd__xor2_1
XU$$2244 net1101 net571 net1092 net844 VGND VGND VPWR VPWR t$5552 sky130_fd_sc_hd__a22o_1
XU$$1510 net1481 notblock$5175\[1\] VGND VGND VPWR VPWR t$5176 sky130_fd_sc_hd__and2_1
XFILLER_23_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2255 t$5557 net1431 VGND VGND VPWR VPWR booth_b32_m28 sky130_fd_sc_hd__xor2_1
XU$$1521 net932 net610 net1671 net883 VGND VGND VPWR VPWR t$5183 sky130_fd_sc_hd__a22o_1
XU$$2266 net993 net572 net989 net845 VGND VGND VPWR VPWR t$5563 sky130_fd_sc_hd__a22o_1
XU$$1532 t$5188 net1476 VGND VGND VPWR VPWR booth_b22_m9 sky130_fd_sc_hd__xor2_1
XU$$2277 t$5568 net1434 VGND VGND VPWR VPWR booth_b32_m39 sky130_fd_sc_hd__xor2_1
XU$$2288 net1721 net573 net1712 net846 VGND VGND VPWR VPWR t$5574 sky130_fd_sc_hd__a22o_1
XU$$1543 net1179 net613 net1170 net886 VGND VGND VPWR VPWR t$5194 sky130_fd_sc_hd__a22o_1
XU$$2299 t$5579 net1434 VGND VGND VPWR VPWR booth_b32_m50 sky130_fd_sc_hd__xor2_1
XU$$1554 t$5199 net1475 VGND VGND VPWR VPWR booth_b22_m20 sky130_fd_sc_hd__xor2_1
XU$$1565 net1073 net612 net1064 net885 VGND VGND VPWR VPWR t$5205 sky130_fd_sc_hd__a22o_1
XU$$1576 t$5210 net1479 VGND VGND VPWR VPWR booth_b22_m31 sky130_fd_sc_hd__xor2_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1587 net965 net615 net957 net888 VGND VGND VPWR VPWR t$5216 sky130_fd_sc_hd__a22o_1
X_1912_ clknet_leaf_31_clk booth_b52_m0 VGND VGND VPWR VPWR pp_row52_26 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_7_122_0 s$3887 c$4138 s$4141 VGND VGND VPWR VPWR c$4396 s$4397 sky130_fd_sc_hd__fa_1
XFILLER_176_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1598 t$5221 net1484 VGND VGND VPWR VPWR booth_b22_m42 sky130_fd_sc_hd__xor2_1
XFILLER_30_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1843_ clknet_leaf_71_clk booth_b36_m14 VGND VGND VPWR VPWR pp_row50_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_129_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1774_ clknet_leaf_238_clk booth_b18_m30 VGND VGND VPWR VPWR pp_row48_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_144_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_87_1 s$3213 s$3215 s$3217 VGND VGND VPWR VPWR c$3746 s$3747 sky130_fd_sc_hd__fa_1
X_0725_ clknet_leaf_135_clk booth_b32_m56 VGND VGND VPWR VPWR pp_row88_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_144_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0656_ clknet_leaf_178_clk booth_b44_m41 VGND VGND VPWR VPWR pp_row85_12 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_6_clk clknet_5_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_170_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0587_ clknet_leaf_186_clk notsign$5104 VGND VGND VPWR VPWR pp_row83_0 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_79_8 pp_row79_24 pp_row79_25 pp_row79_26 VGND VGND VPWR VPWR c$886 s$887
+ sky130_fd_sc_hd__fa_2
XFILLER_97_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2326_ clknet_leaf_74_clk booth_b54_m10 VGND VGND VPWR VPWR pp_row64_27 sky130_fd_sc_hd__dfxtp_1
XFILLER_170_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$206 final_adder.$signal$1138 final_adder.$signal$101 VGND VGND VPWR
+ VPWR final_adder.p_new$334 sky130_fd_sc_hd__and2_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$217 final_adder.$signal$1129 final_adder.$signal$78 final_adder.$signal$80
+ VGND VGND VPWR VPWR final_adder.g_new$345 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$228 final_adder.$signal$1116 final_adder.$signal$1117 VGND VGND VPWR
+ VPWR final_adder.p_new$356 sky130_fd_sc_hd__and2_1
X_2257_ clknet_leaf_227_clk net1254 VGND VGND VPWR VPWR pp_row62_32 sky130_fd_sc_hd__dfxtp_1
XFILLER_111_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$239 final_adder.$signal$1107 final_adder.$signal$34 final_adder.$signal$36
+ VGND VGND VPWR VPWR final_adder.g_new$367 sky130_fd_sc_hd__a21o_1
XFILLER_27_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1208_ clknet_leaf_47_clk booth_b14_m8 VGND VGND VPWR VPWR pp_row22_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_150_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2188_ clknet_leaf_227_clk booth_b2_m59 VGND VGND VPWR VPWR pp_row61_1 sky130_fd_sc_hd__dfxtp_1
XU$$4180 net1021 net441 net1004 net723 VGND VGND VPWR VPWR t$6541 sky130_fd_sc_hd__a22o_1
XU$$4191 t$6546 net1272 VGND VGND VPWR VPWR booth_b60_m37 sky130_fd_sc_hd__xor2_1
XFILLER_38_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1139_ clknet_leaf_16_clk booth_b6_m11 VGND VGND VPWR VPWR pp_row17_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_81_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3490 t$6188 net1331 VGND VGND VPWR VPWR booth_b50_m29 sky130_fd_sc_hd__xor2_1
XFILLER_41_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_82_0 s$1721 c$2486 c$2488 VGND VGND VPWR VPWR c$3182 s$3183 sky130_fd_sc_hd__fa_1
XFILLER_190_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_103_3 c$1948 s$1951 s$1953 VGND VGND VPWR VPWR c$2668 s$2669 sky130_fd_sc_hd__fa_1
XFILLER_150_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput202 c[50] VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_1
Xinput213 c[60] VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_1
XFILLER_68_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput224 c[70] VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput235 c[80] VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_5_26__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_5_26__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xinput246 c[90] VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__clkbuf_1
XFILLER_124_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$740 final_adder.p_new$788 final_adder.p_new$756 VGND VGND VPWR VPWR
+ final_adder.p_new$868 sky130_fd_sc_hd__and2_1
XFILLER_25_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$751 final_adder.p_new$766 final_adder.g_new$799 final_adder.g_new$767
+ VGND VGND VPWR VPWR final_adder.g_new$879 sky130_fd_sc_hd__a21o_1
XFILLER_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$762 final_adder.p_new$810 final_adder.p_new$778 VGND VGND VPWR VPWR
+ final_adder.p_new$890 sky130_fd_sc_hd__and2_1
XU$$601 t$4712 net1236 VGND VGND VPWR VPWR booth_b8_m23 sky130_fd_sc_hd__xor2_1
XFILLER_99_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_883 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$612 net1049 net415 net1041 net681 VGND VGND VPWR VPWR t$4718 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$773 final_adder.p_new$788 final_adder.g_new$821 final_adder.g_new$789
+ VGND VGND VPWR VPWR final_adder.g_new$901 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$784 final_adder.p_new$832 final_adder.p_new$800 VGND VGND VPWR VPWR
+ final_adder.p_new$912 sky130_fd_sc_hd__and2_1
XU$$623 t$4723 net1235 VGND VGND VPWR VPWR booth_b8_m34 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$795 final_adder.p_new$810 final_adder.g_new$843 final_adder.g_new$811
+ VGND VGND VPWR VPWR final_adder.g_new$923 sky130_fd_sc_hd__a21o_1
XU$$634 net940 net411 net924 net677 VGND VGND VPWR VPWR t$4729 sky130_fd_sc_hd__a22o_1
XFILLER_186_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$645 t$4734 net1242 VGND VGND VPWR VPWR booth_b8_m45 sky130_fd_sc_hd__xor2_1
XFILLER_189_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$656 net1654 net411 net1646 net677 VGND VGND VPWR VPWR t$4740 sky130_fd_sc_hd__a22o_1
XU$$667 t$4745 net1237 VGND VGND VPWR VPWR booth_b8_m56 sky130_fd_sc_hd__xor2_1
XU$$678 net1547 net416 net1539 net682 VGND VGND VPWR VPWR t$4751 sky130_fd_sc_hd__a22o_1
XFILLER_17_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$689 notblock$4755\[2\] net2 net1238 t$4756 notblock$4755\[0\] VGND VGND VPWR VPWR
+ sel_0$4757 sky130_fd_sc_hd__a32o_1
XFILLER_140_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_97_0 c$3780 c$3782 s$3785 VGND VGND VPWR VPWR c$4090 s$4091 sky130_fd_sc_hd__fa_1
XFILLER_157_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0510_ clknet_leaf_173_clk booth_b30_m50 VGND VGND VPWR VPWR pp_row80_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1490_ clknet_leaf_44_clk booth_b18_m19 VGND VGND VPWR VPWR pp_row37_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_126_899 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0441_ clknet_leaf_197_clk net231 VGND VGND VPWR VPWR pp_row77_27 sky130_fd_sc_hd__dfxtp_1
X_0372_ clknet_leaf_203_clk booth_b54_m21 VGND VGND VPWR VPWR pp_row75_22 sky130_fd_sc_hd__dfxtp_1
Xdadda_ha_2_33_5 pp_row33_15 pp_row33_16 VGND VGND VPWR VPWR c$1132 s$1133 sky130_fd_sc_hd__ha_1
X_2111_ clknet_leaf_85_clk booth_b56_m2 VGND VGND VPWR VPWR pp_row58_28 sky130_fd_sc_hd__dfxtp_1
XFILLER_66_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2042_ clknet_leaf_82_clk booth_b54_m2 VGND VGND VPWR VPWR pp_row56_27 sky130_fd_sc_hd__dfxtp_1
XFILLER_66_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_32_3 pp_row32_9 pp_row32_10 pp_row32_11 VGND VGND VPWR VPWR c$1116 s$1117
+ sky130_fd_sc_hd__fa_1
XU$$2030 net1639 net590 net1631 net863 VGND VGND VPWR VPWR t$5442 sky130_fd_sc_hd__a22o_1
XU$$2041 t$5447 net1453 VGND VGND VPWR VPWR booth_b28_m58 sky130_fd_sc_hd__xor2_1
XU$$2052 net1532 net591 net1770 net864 VGND VGND VPWR VPWR t$5453 sky130_fd_sc_hd__a22o_1
XU$$2063 net1227 net576 net1122 net849 VGND VGND VPWR VPWR t$5460 sky130_fd_sc_hd__a22o_1
XU$$2074 t$5465 net1441 VGND VGND VPWR VPWR booth_b30_m6 sky130_fd_sc_hd__xor2_1
XU$$1340 t$5089 net1670 VGND VGND VPWR VPWR booth_b18_m50 sky130_fd_sc_hd__xor2_1
XU$$2085 net1210 net576 net1201 net849 VGND VGND VPWR VPWR t$5471 sky130_fd_sc_hd__a22o_1
XU$$2096 t$5476 net1440 VGND VGND VPWR VPWR booth_b30_m17 sky130_fd_sc_hd__xor2_1
XU$$1351 net1612 net640 net1604 net913 VGND VGND VPWR VPWR t$5095 sky130_fd_sc_hd__a22o_1
XFILLER_16_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1362 t$5100 net1668 VGND VGND VPWR VPWR booth_b18_m61 sky130_fd_sc_hd__xor2_1
XFILLER_149_914 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1373 net1491 notblock$5105\[1\] VGND VGND VPWR VPWR t$5106 sky130_fd_sc_hd__and2_1
XU$$1384 net933 net627 net1672 net900 VGND VGND VPWR VPWR t$5113 sky130_fd_sc_hd__a22o_1
XU$$1395 t$5118 net1485 VGND VGND VPWR VPWR booth_b20_m9 sky130_fd_sc_hd__xor2_1
XFILLER_128_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1826_ clknet_leaf_234_clk booth_b8_m42 VGND VGND VPWR VPWR pp_row50_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_159_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1757_ clknet_leaf_239_clk booth_b38_m9 VGND VGND VPWR VPWR pp_row47_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0708_ clknet_leaf_168_clk booth_b48_m39 VGND VGND VPWR VPWR pp_row87_13 sky130_fd_sc_hd__dfxtp_1
X_1688_ clknet_leaf_18_clk booth_b14_m31 VGND VGND VPWR VPWR pp_row45_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_116_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout903 net904 VGND VGND VPWR VPWR net903 sky130_fd_sc_hd__buf_6
XFILLER_132_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0639_ clknet_leaf_188_clk booth_b62_m22 VGND VGND VPWR VPWR pp_row84_22 sky130_fd_sc_hd__dfxtp_1
Xfanout914 net915 VGND VGND VPWR VPWR net914 sky130_fd_sc_hd__clkbuf_4
Xfanout925 net931 VGND VGND VPWR VPWR net925 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_77_5 pp_row77_18 pp_row77_19 pp_row77_20 VGND VGND VPWR VPWR c$844 s$845
+ sky130_fd_sc_hd__fa_1
Xfanout936 net939 VGND VGND VPWR VPWR net936 sky130_fd_sc_hd__buf_4
Xfanout947 net97 VGND VGND VPWR VPWR net947 sky130_fd_sc_hd__buf_12
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout958 net959 VGND VGND VPWR VPWR net958 sky130_fd_sc_hd__buf_6
XTAP_4008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout969 net972 VGND VGND VPWR VPWR net969 sky130_fd_sc_hd__buf_4
XTAP_4019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2309_ clknet_leaf_91_clk booth_b22_m42 VGND VGND VPWR VPWR pp_row64_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_161_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_307 net450 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_318 net588 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_329 net683 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$80 c$4310 s$4313 VGND VGND VPWR VPWR final_adder.$signal$162 final_adder.$signal$1170
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$91 c$4332 s$4335 VGND VGND VPWR VPWR final_adder.$signal$184 final_adder.$signal$1181
+ sky130_fd_sc_hd__ha_2
XFILLER_80_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_101_0 pp_row101_12 pp_row101_13 pp_row101_14 VGND VGND VPWR VPWR c$2646
+ s$2647 sky130_fd_sc_hd__fa_1
XFILLER_107_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_65_3 pp_row65_9 pp_row65_10 pp_row65_11 VGND VGND VPWR VPWR c$102 s$103
+ sky130_fd_sc_hd__fa_1
XFILLER_114_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_42_2 c$1228 s$1231 s$1233 VGND VGND VPWR VPWR c$2178 s$2179 sky130_fd_sc_hd__fa_1
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_0_58_2 pp_row58_6 pp_row58_7 pp_row58_8 VGND VGND VPWR VPWR c$28 s$29 sky130_fd_sc_hd__fa_1
XTAP_3830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$570 final_adder.p_new$582 final_adder.p_new$574 VGND VGND VPWR VPWR
+ final_adder.p_new$698 sky130_fd_sc_hd__and2_1
Xdadda_fa_3_35_1 c$1138 c$1140 c$1142 VGND VGND VPWR VPWR c$2120 s$2121 sky130_fd_sc_hd__fa_1
XTAP_3852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$420 t$4620 net1248 VGND VGND VPWR VPWR booth_b6_m1 sky130_fd_sc_hd__xor2_1
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$581 final_adder.p_new$584 final_adder.g_new$593 final_adder.g_new$585
+ VGND VGND VPWR VPWR final_adder.g_new$709 sky130_fd_sc_hd__a21o_1
XTAP_3863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$592 final_adder.p_new$604 final_adder.p_new$596 VGND VGND VPWR VPWR
+ final_adder.p_new$720 sky130_fd_sc_hd__and2_1
XU$$431 net1523 net429 net1515 net711 VGND VGND VPWR VPWR t$4626 sky130_fd_sc_hd__a22o_1
XTAP_3874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$442 t$4631 net1250 VGND VGND VPWR VPWR booth_b6_m12 sky130_fd_sc_hd__xor2_1
XTAP_3885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$453 net1147 net427 net1139 net709 VGND VGND VPWR VPWR t$4637 sky130_fd_sc_hd__a22o_1
Xdadda_fa_6_12_0 c$3440 c$3442 s$3445 VGND VGND VPWR VPWR c$3920 s$3921 sky130_fd_sc_hd__fa_1
XTAP_3896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$464 t$4642 net1244 VGND VGND VPWR VPWR booth_b6_m23 sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_28_0 pp_row28_11 pp_row28_12 pp_row28_13 VGND VGND VPWR VPWR c$2062 s$2063
+ sky130_fd_sc_hd__fa_1
XFILLER_189_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$475 net1050 net429 net1042 net711 VGND VGND VPWR VPWR t$4648 sky130_fd_sc_hd__a22o_1
XU$$486 t$4653 net1245 VGND VGND VPWR VPWR booth_b6_m34 sky130_fd_sc_hd__xor2_1
XU$$497 net940 net427 net924 net709 VGND VGND VPWR VPWR t$4659 sky130_fd_sc_hd__a22o_1
XFILLER_44_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0990_ clknet_leaf_118_clk booth_b54_m46 VGND VGND VPWR VPWR pp_row100_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_9_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1611_ clknet_leaf_239_clk booth_b20_m22 VGND VGND VPWR VPWR pp_row42_10 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_94_5 c$1038 c$1040 s$1043 VGND VGND VPWR VPWR c$1864 s$1865 sky130_fd_sc_hd__fa_1
X_1542_ clknet_leaf_12_clk booth_b26_m13 VGND VGND VPWR VPWR pp_row39_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_114_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_87_4 c$986 c$988 s$991 VGND VGND VPWR VPWR c$1778 s$1779 sky130_fd_sc_hd__fa_1
XFILLER_99_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1473_ clknet_leaf_39_clk booth_b28_m8 VGND VGND VPWR VPWR pp_row36_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_68_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0424_ clknet_leaf_211_clk booth_b34_m43 VGND VGND VPWR VPWR pp_row77_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_95_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0355_ clknet_leaf_125_clk booth_b54_m60 VGND VGND VPWR VPWR pp_row114_3 sky130_fd_sc_hd__dfxtp_1
Xdadda_ha_2_24_1 pp_row24_3 pp_row24_4 VGND VGND VPWR VPWR c$1056 s$1057 sky130_fd_sc_hd__ha_1
Xclkbuf_leaf_230_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_230_clk
+ sky130_fd_sc_hd__clkbuf_16
X_0286_ clknet_leaf_203_clk booth_b14_m59 VGND VGND VPWR VPWR pp_row73_3 sky130_fd_sc_hd__dfxtp_1
X_2025_ clknet_leaf_36_clk booth_b24_m32 VGND VGND VPWR VPWR pp_row56_12 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_30_0 pp_row30_0 pp_row30_1 pp_row30_2 VGND VGND VPWR VPWR c$1090 s$1091
+ sky130_fd_sc_hd__fa_1
XFILLER_36_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_103_2 pp_row103_6 pp_row103_7 pp_row103_8 VGND VGND VPWR VPWR c$1954 s$1955
+ sky130_fd_sc_hd__fa_1
XFILLER_23_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1170 net990 net645 net983 net918 VGND VGND VPWR VPWR t$5003 sky130_fd_sc_hd__a22o_1
XU$$1181 t$5008 net1010 VGND VGND VPWR VPWR booth_b16_m39 sky130_fd_sc_hd__xor2_1
XU$$1192 net1720 net648 net1711 net921 VGND VGND VPWR VPWR t$5014 sky130_fd_sc_hd__a22o_1
XFILLER_108_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_117_0 c$3386 c$3388 c$3390 VGND VGND VPWR VPWR c$3864 s$3865 sky130_fd_sc_hd__fa_1
XFILLER_163_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1809_ clknet_leaf_24_clk booth_b28_m21 VGND VGND VPWR VPWR pp_row49_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_82_3 pp_row82_9 pp_row82_10 pp_row82_11 VGND VGND VPWR VPWR c$928 s$929
+ sky130_fd_sc_hd__fa_1
XFILLER_172_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout700 net703 VGND VGND VPWR VPWR net700 sky130_fd_sc_hd__clkbuf_8
XFILLER_172_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1709 net1710 VGND VGND VPWR VPWR net1709 sky130_fd_sc_hd__clkbuf_2
Xfanout711 net712 VGND VGND VPWR VPWR net711 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_75_2 pp_row75_12 pp_row75_13 pp_row75_14 VGND VGND VPWR VPWR c$802 s$803
+ sky130_fd_sc_hd__fa_1
Xfanout722 net723 VGND VGND VPWR VPWR net722 sky130_fd_sc_hd__buf_4
Xfanout733 net734 VGND VGND VPWR VPWR net733 sky130_fd_sc_hd__buf_4
XFILLER_132_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout744 sel_1$6298 VGND VGND VPWR VPWR net744 sky130_fd_sc_hd__clkbuf_4
Xfanout755 net756 VGND VGND VPWR VPWR net755 sky130_fd_sc_hd__buf_4
XFILLER_98_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_52_1 c$2250 c$2252 s$2255 VGND VGND VPWR VPWR c$3004 s$3005 sky130_fd_sc_hd__fa_1
Xdadda_fa_1_68_1 pp_row68_20 pp_row68_21 pp_row68_22 VGND VGND VPWR VPWR c$674 s$675
+ sky130_fd_sc_hd__fa_1
Xfanout766 net769 VGND VGND VPWR VPWR net766 sky130_fd_sc_hd__buf_4
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_967 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout777 net782 VGND VGND VPWR VPWR net777 sky130_fd_sc_hd__clkbuf_4
Xfanout788 net789 VGND VGND VPWR VPWR net788 sky130_fd_sc_hd__buf_4
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout799 sel_1$5878 VGND VGND VPWR VPWR net799 sky130_fd_sc_hd__clkbuf_8
Xdadda_fa_4_45_0 s$1277 c$2190 c$2192 VGND VGND VPWR VPWR c$2960 s$2961 sky130_fd_sc_hd__fa_1
Xclkbuf_leaf_221_clk clknet_5_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_221_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_85_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_104 net575 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_115 net631 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 net683 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_137 net740 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_148 net791 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_159 net848 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_97_3 s$1895 s$1897 s$1899 VGND VGND VPWR VPWR c$2620 s$2621 sky130_fd_sc_hd__fa_1
XFILLER_6_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_0_70_1 pp_row70_3 pp_row70_4 pp_row70_5 VGND VGND VPWR VPWR c$156 s$157
+ sky130_fd_sc_hd__fa_1
XFILLER_7_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_0_63_0 pp_row63_0 pp_row63_1 pp_row63_2 VGND VGND VPWR VPWR c$72 s$73 sky130_fd_sc_hd__fa_1
Xclkbuf_leaf_212_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_212_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_65_926 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$250 t$4532 net1392 VGND VGND VPWR VPWR booth_b2_m53 sky130_fd_sc_hd__xor2_1
XTAP_3693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$261 net1586 net621 net1578 net894 VGND VGND VPWR VPWR t$4538 sky130_fd_sc_hd__a22o_1
XU$$272 t$4543 net1392 VGND VGND VPWR VPWR booth_b2_m64 sky130_fd_sc_hd__xor2_1
XU$$283 t$4550 net1277 VGND VGND VPWR VPWR booth_b4_m1 sky130_fd_sc_hd__xor2_1
XTAP_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4425_1833 VGND VGND VPWR VPWR U$$4425_1833/HI net1833 sky130_fd_sc_hd__conb_1
XTAP_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$294 net1523 net531 net1515 net804 VGND VGND VPWR VPWR t$4556 sky130_fd_sc_hd__a22o_1
XFILLER_177_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0973_ clknet_leaf_117_clk booth_b56_m43 VGND VGND VPWR VPWR pp_row99_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_146_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$0 net1753 VGND VGND VPWR VPWR notblock\[0\] sky130_fd_sc_hd__inv_1
XFILLER_69_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$8 c$4166 s$4169 VGND VGND VPWR VPWR final_adder.$signal$18 final_adder.$signal$1098
+ sky130_fd_sc_hd__ha_1
XFILLER_69_1018 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput303 net303 VGND VGND VPWR VPWR o[26] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_92_2 pp_row92_14 pp_row92_15 pp_row92_16 VGND VGND VPWR VPWR c$1834 s$1835
+ sky130_fd_sc_hd__fa_1
Xoutput314 net314 VGND VGND VPWR VPWR o[36] sky130_fd_sc_hd__buf_2
XFILLER_145_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput325 net325 VGND VGND VPWR VPWR o[46] sky130_fd_sc_hd__buf_2
XFILLER_160_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput336 net336 VGND VGND VPWR VPWR o[56] sky130_fd_sc_hd__buf_2
XFILLER_99_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput347 net347 VGND VGND VPWR VPWR o[66] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_85_1 pp_row85_21 pp_row85_22 pp_row85_23 VGND VGND VPWR VPWR c$1748 s$1749
+ sky130_fd_sc_hd__fa_1
XFILLER_126_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput358 net358 VGND VGND VPWR VPWR o[76] sky130_fd_sc_hd__buf_2
Xoutput369 net369 VGND VGND VPWR VPWR o[86] sky130_fd_sc_hd__buf_2
X_1525_ clknet_leaf_241_clk net1394 VGND VGND VPWR VPWR pp_row38_20 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_62_0 c$3056 c$3058 c$3060 VGND VGND VPWR VPWR c$3644 s$3645 sky130_fd_sc_hd__fa_1
Xdadda_fa_2_78_0 s$203 c$834 c$836 VGND VGND VPWR VPWR c$1662 s$1663 sky130_fd_sc_hd__fa_1
XFILLER_113_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1456_ clknet_leaf_244_clk net185 VGND VGND VPWR VPWR pp_row35_18 sky130_fd_sc_hd__dfxtp_2
Xdadda_fa_1_61_8 s$53 s$55 s$57 VGND VGND VPWR VPWR c$562 s$563 sky130_fd_sc_hd__fa_2
X_0407_ clknet_leaf_205_clk booth_b60_m16 VGND VGND VPWR VPWR pp_row76_25 sky130_fd_sc_hd__dfxtp_1
X_1387_ clknet_leaf_42_clk booth_b28_m4 VGND VGND VPWR VPWR pp_row32_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_45_1095 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_775 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_203_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_203_clk
+ sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_1_54_7 pp_row54_26 pp_row54_27 pp_row54_28 VGND VGND VPWR VPWR c$434 s$435
+ sky130_fd_sc_hd__fa_1
X_0338_ clknet_leaf_225_clk booth_b50_m24 VGND VGND VPWR VPWR pp_row74_21 sky130_fd_sc_hd__dfxtp_1
X_0269_ clknet_leaf_217_clk booth_b44_m28 VGND VGND VPWR VPWR pp_row72_19 sky130_fd_sc_hd__dfxtp_1
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2008_ clknet_leaf_72_clk booth_b50_m5 VGND VGND VPWR VPWR pp_row55_25 sky130_fd_sc_hd__dfxtp_1
XFILLER_42_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_77_0 s$3707 c$4048 s$4051 VGND VGND VPWR VPWR c$4306 s$4307 sky130_fd_sc_hd__fa_2
XFILLER_191_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_80_0 net1896 pp_row80_1 pp_row80_2 VGND VGND VPWR VPWR c$888 s$889 sky130_fd_sc_hd__fa_1
Xfanout1506 net1507 VGND VGND VPWR VPWR net1506 sky130_fd_sc_hd__clkbuf_4
XFILLER_105_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1517 net1518 VGND VGND VPWR VPWR net1517 sky130_fd_sc_hd__buf_4
Xfanout530 sel_0$4547 VGND VGND VPWR VPWR net530 sky130_fd_sc_hd__buf_6
Xfanout1528 net1530 VGND VGND VPWR VPWR net1528 sky130_fd_sc_hd__buf_4
XFILLER_132_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1539 net123 VGND VGND VPWR VPWR net1539 sky130_fd_sc_hd__buf_4
Xfanout541 net542 VGND VGND VPWR VPWR net541 sky130_fd_sc_hd__clkbuf_4
Xfanout552 net553 VGND VGND VPWR VPWR net552 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4009 net1177 net451 net1168 net724 VGND VGND VPWR VPWR t$6454 sky130_fd_sc_hd__a22o_1
Xfanout563 net564 VGND VGND VPWR VPWR net563 sky130_fd_sc_hd__buf_4
Xfanout574 net575 VGND VGND VPWR VPWR net574 sky130_fd_sc_hd__buf_4
XFILLER_150_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout585 net586 VGND VGND VPWR VPWR net585 sky130_fd_sc_hd__clkbuf_4
XFILLER_74_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout596 net597 VGND VGND VPWR VPWR net596 sky130_fd_sc_hd__buf_4
XU$$3308 net1525 net497 net1517 net770 VGND VGND VPWR VPWR t$6096 sky130_fd_sc_hd__a22o_1
XFILLER_150_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3319 t$6101 net1338 VGND VGND VPWR VPWR booth_b48_m12 sky130_fd_sc_hd__xor2_1
XFILLER_73_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2607 notblock$5735\[2\] net32 net1408 t$5736 notblock$5735\[0\] VGND VGND VPWR
+ VPWR sel_0$5737 sky130_fd_sc_hd__a32o_1
XU$$2618 t$5743 net1394 VGND VGND VPWR VPWR booth_b38_m4 sky130_fd_sc_hd__xor2_1
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2629 net1495 net543 net1220 net816 VGND VGND VPWR VPWR t$5749 sky130_fd_sc_hd__a22o_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1906 t$5378 net1463 VGND VGND VPWR VPWR booth_b26_m59 sky130_fd_sc_hd__xor2_1
XFILLER_73_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_992 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1917 net20 VGND VGND VPWR VPWR notsign$5384 sky130_fd_sc_hd__inv_1
XU$$1928 net1122 net584 net1031 net857 VGND VGND VPWR VPWR t$5391 sky130_fd_sc_hd__a22o_1
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1939 t$5396 net1451 VGND VGND VPWR VPWR booth_b28_m7 sky130_fd_sc_hd__xor2_1
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_95_0 s$1047 c$1854 c$1856 VGND VGND VPWR VPWR c$2598 s$2599 sky130_fd_sc_hd__fa_1
XFILLER_6_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4455_1848 VGND VGND VPWR VPWR U$$4455_1848/HI net1848 sky130_fd_sc_hd__conb_1
XFILLER_182_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1310_ clknet_leaf_2_clk booth_b24_m4 VGND VGND VPWR VPWR pp_row28_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_97_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2290_ clknet_leaf_216_clk booth_b54_m9 VGND VGND VPWR VPWR pp_row63_27 sky130_fd_sc_hd__dfxtp_1
XFILLER_173_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1241_ clknet_leaf_13_clk booth_b20_m4 VGND VGND VPWR VPWR pp_row24_10 sky130_fd_sc_hd__dfxtp_1
XU$$6_1883 VGND VGND VPWR VPWR U$$6_1883/HI net1883 sky130_fd_sc_hd__conb_1
XFILLER_77_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4510 net1580 sel_0$6647 net1554 net695 VGND VGND VPWR VPWR t$6709 sky130_fd_sc_hd__a22o_1
XFILLER_49_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_57_5 s$485 s$487 s$489 VGND VGND VPWR VPWR c$1420 s$1421 sky130_fd_sc_hd__fa_2
X_1172_ clknet_leaf_129_clk booth_b64_m58 VGND VGND VPWR VPWR pp_row122_4 sky130_fd_sc_hd__dfxtp_1
XU$$13 t$4413 net1573 VGND VGND VPWR VPWR booth_b0_m3 sky130_fd_sc_hd__xor2_1
XFILLER_37_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$24 net1508 net446 net1499 net688 VGND VGND VPWR VPWR t$4419 sky130_fd_sc_hd__a22o_1
XU$$35 t$4424 net1575 VGND VGND VPWR VPWR booth_b0_m14 sky130_fd_sc_hd__xor2_1
XU$$3820 t$6356 net1306 VGND VGND VPWR VPWR booth_b54_m57 sky130_fd_sc_hd__xor2_1
XU$$3831 net1537 net469 net1529 net742 VGND VGND VPWR VPWR t$6362 sky130_fd_sc_hd__a22o_1
XU$$46 net1133 net448 net1117 net690 VGND VGND VPWR VPWR t$4430 sky130_fd_sc_hd__a22o_1
XTAP_4180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$57 t$4435 net1569 VGND VGND VPWR VPWR booth_b0_m25 sky130_fd_sc_hd__xor2_1
XU$$3842 net1799 net464 net1233 net737 VGND VGND VPWR VPWR t$6369 sky130_fd_sc_hd__a22o_1
XTAP_4191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3853 t$6374 net1291 VGND VGND VPWR VPWR booth_b56_m5 sky130_fd_sc_hd__xor2_1
XU$$3864 net1226 net467 net1217 net740 VGND VGND VPWR VPWR t$6380 sky130_fd_sc_hd__a22o_1
XU$$68 net1023 net442 net1015 net684 VGND VGND VPWR VPWR t$4441 sky130_fd_sc_hd__a22o_1
XFILLER_24_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$79 t$4446 net1575 VGND VGND VPWR VPWR booth_b0_m36 sky130_fd_sc_hd__xor2_1
XU$$3875 t$6385 net1291 VGND VGND VPWR VPWR booth_b56_m16 sky130_fd_sc_hd__xor2_1
XFILLER_92_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3886 net1111 net461 net1102 net734 VGND VGND VPWR VPWR t$6391 sky130_fd_sc_hd__a22o_1
XFILLER_52_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3897 t$6396 net1294 VGND VGND VPWR VPWR booth_b56_m27 sky130_fd_sc_hd__xor2_1
XFILLER_21_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_15 s$4405 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_26 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_37 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_59 net392 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0956_ clknet_leaf_116_clk booth_b58_m40 VGND VGND VPWR VPWR pp_row98_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_107_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0887_ clknet_leaf_100_clk booth_b42_m53 VGND VGND VPWR VPWR pp_row95_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1508_ clknet_leaf_16_clk booth_b8_m30 VGND VGND VPWR VPWR pp_row38_4 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_5_7__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_5_7__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_101_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2488_ clknet_leaf_90_clk booth_b18_m51 VGND VGND VPWR VPWR pp_row69_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_134_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1439_ clknet_leaf_121_clk booth_b58_m46 VGND VGND VPWR VPWR pp_row104_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_52_4 pp_row52_14 pp_row52_15 pp_row52_16 VGND VGND VPWR VPWR c$392 s$393
+ sky130_fd_sc_hd__fa_1
XFILLER_29_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_45_3 pp_row45_9 pp_row45_10 pp_row45_11 VGND VGND VPWR VPWR c$282 s$283
+ sky130_fd_sc_hd__fa_1
XFILLER_71_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_22_2 s$2017 s$2019 s$2021 VGND VGND VPWR VPWR c$2826 s$2827 sky130_fd_sc_hd__fa_1
Xdadda_fa_4_15_1 pp_row15_5 pp_row15_6 pp_row15_7 VGND VGND VPWR VPWR c$2782 s$2783
+ sky130_fd_sc_hd__fa_1
XFILLER_178_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$1007 final_adder.$signal$1136 final_adder.g_new$949 VGND VGND VPWR
+ VPWR net325 sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$1018 final_adder.$signal$1147 final_adder.g_new$1061 VGND VGND VPWR
+ VPWR net337 sky130_fd_sc_hd__xor2_1
XFILLER_137_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1029 final_adder.$signal$1158 final_adder.g_new$1023 VGND VGND VPWR
+ VPWR net349 sky130_fd_sc_hd__xor2_2
XFILLER_164_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1303 net1309 VGND VGND VPWR VPWR net1303 sky130_fd_sc_hd__buf_6
Xfanout1314 net1315 VGND VGND VPWR VPWR net1314 sky130_fd_sc_hd__buf_6
Xfanout1325 net1328 VGND VGND VPWR VPWR net1325 sky130_fd_sc_hd__buf_4
XFILLER_121_967 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1336 net1337 VGND VGND VPWR VPWR net1336 sky130_fd_sc_hd__clkbuf_4
Xfanout1347 net44 VGND VGND VPWR VPWR net1347 sky130_fd_sc_hd__buf_4
XFILLER_28_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1358 net1366 VGND VGND VPWR VPWR net1358 sky130_fd_sc_hd__buf_6
Xfanout1369 net1370 VGND VGND VPWR VPWR net1369 sky130_fd_sc_hd__buf_4
XFILLER_120_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout393 net394 VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__buf_4
XFILLER_4_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3105 t$5991 net1361 VGND VGND VPWR VPWR booth_b44_m42 sky130_fd_sc_hd__xor2_1
XU$$3116 net1700 net515 net1693 net788 VGND VGND VPWR VPWR t$5997 sky130_fd_sc_hd__a22o_1
XU$$3127 t$6002 net1364 VGND VGND VPWR VPWR booth_b44_m53 sky130_fd_sc_hd__xor2_1
XFILLER_98_1055 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3138 net1590 net513 net1582 net786 VGND VGND VPWR VPWR t$6008 sky130_fd_sc_hd__a22o_1
XU$$2404 t$5633 net1428 VGND VGND VPWR VPWR booth_b34_m34 sky130_fd_sc_hd__xor2_1
XU$$3149 t$6013 net1360 VGND VGND VPWR VPWR booth_b44_m64 sky130_fd_sc_hd__xor2_1
XU$$2415 net941 net562 net925 net835 VGND VGND VPWR VPWR t$5639 sky130_fd_sc_hd__a22o_1
XU$$2426 t$5644 net1425 VGND VGND VPWR VPWR booth_b34_m45 sky130_fd_sc_hd__xor2_1
XU$$2437 net1656 net566 net1648 net839 VGND VGND VPWR VPWR t$5650 sky130_fd_sc_hd__a22o_1
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1703 t$5275 net1468 VGND VGND VPWR VPWR booth_b24_m26 sky130_fd_sc_hd__xor2_1
XU$$2448 t$5655 net1427 VGND VGND VPWR VPWR booth_b34_m56 sky130_fd_sc_hd__xor2_1
XU$$2459 net1547 net567 net123 net840 VGND VGND VPWR VPWR t$5661 sky130_fd_sc_hd__a22o_1
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1714 net1017 net606 net1000 net879 VGND VGND VPWR VPWR t$5281 sky130_fd_sc_hd__a22o_1
XU$$1725 t$5286 net1468 VGND VGND VPWR VPWR booth_b24_m37 sky130_fd_sc_hd__xor2_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1736 net1743 net609 net1735 net882 VGND VGND VPWR VPWR t$5292 sky130_fd_sc_hd__a22o_1
XU$$1747 t$5297 net1473 VGND VGND VPWR VPWR booth_b24_m48 sky130_fd_sc_hd__xor2_1
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1758 net1630 net607 net1621 net880 VGND VGND VPWR VPWR t$5303 sky130_fd_sc_hd__a22o_1
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1769 t$5308 net1471 VGND VGND VPWR VPWR booth_b24_m59 sky130_fd_sc_hd__xor2_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0810_ clknet_leaf_132_clk booth_b58_m61 VGND VGND VPWR VPWR pp_row119_2 sky130_fd_sc_hd__dfxtp_1
Xinput13 a[20] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_2
X_1790_ clknet_leaf_221_clk booth_b48_m0 VGND VGND VPWR VPWR pp_row48_24 sky130_fd_sc_hd__dfxtp_1
Xinput24 a[30] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput35 a[40] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dlymetal6s2s_1
X_0741_ clknet_leaf_171_clk booth_b62_m26 VGND VGND VPWR VPWR pp_row88_20 sky130_fd_sc_hd__dfxtp_1
Xinput46 a[50] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_2
Xinput57 a[60] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput68 b[12] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_2
XFILLER_171_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput79 b[22] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__buf_4
X_0672_ clknet_leaf_175_clk booth_b28_m58 VGND VGND VPWR VPWR pp_row86_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_192_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2411_ clknet_leaf_77_clk booth_b6_m61 VGND VGND VPWR VPWR pp_row67_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_124_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2342_ clknet_leaf_89_clk booth_b16_m49 VGND VGND VPWR VPWR pp_row65_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_62_3 c$562 s$565 s$567 VGND VGND VPWR VPWR c$1476 s$1477 sky130_fd_sc_hd__fa_1
X_2273_ clknet_leaf_216_clk booth_b24_m39 VGND VGND VPWR VPWR pp_row63_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_78_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_55_2 c$430 c$432 c$434 VGND VGND VPWR VPWR c$1390 s$1391 sky130_fd_sc_hd__fa_1
XFILLER_37_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1224_ clknet_leaf_48_clk booth_b16_m7 VGND VGND VPWR VPWR pp_row23_8 sky130_fd_sc_hd__dfxtp_1
XU$$4340 t$6622 net1262 VGND VGND VPWR VPWR booth_b62_m43 sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_32_1 s$2883 s$2885 s$2887 VGND VGND VPWR VPWR c$3526 s$3527 sky130_fd_sc_hd__fa_1
XU$$4351 net1692 net423 net1685 net705 VGND VGND VPWR VPWR t$6628 sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_48_1 pp_row48_26 c$302 c$304 VGND VGND VPWR VPWR c$1304 s$1305 sky130_fd_sc_hd__fa_1
XU$$4362 t$6633 net1262 VGND VGND VPWR VPWR booth_b62_m54 sky130_fd_sc_hd__xor2_1
XU$$4373 net1584 net423 net1557 net705 VGND VGND VPWR VPWR t$6639 sky130_fd_sc_hd__a22o_1
XFILLER_77_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1155_ clknet_leaf_15_clk booth_b16_m2 VGND VGND VPWR VPWR pp_row18_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_37_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_25_0 c$2834 c$2836 c$2838 VGND VGND VPWR VPWR c$3496 s$3497 sky130_fd_sc_hd__fa_1
XU$$4384 net1260 VGND VGND VPWR VPWR notblock$6645\[0\] sky130_fd_sc_hd__inv_1
XU$$4395 t$6651 net1818 VGND VGND VPWR VPWR booth_b64_m2 sky130_fd_sc_hd__xor2_1
XU$$3650 net930 net478 net1751 net751 VGND VGND VPWR VPWR t$6270 sky130_fd_sc_hd__a22o_1
XU$$3661 t$6275 net1326 VGND VGND VPWR VPWR booth_b52_m46 sky130_fd_sc_hd__xor2_1
XU$$3672 net1652 net482 net1644 net755 VGND VGND VPWR VPWR t$6281 sky130_fd_sc_hd__a22o_1
X_1086_ clknet_leaf_58_clk booth_b4_m8 VGND VGND VPWR VPWR pp_row12_2 sky130_fd_sc_hd__dfxtp_1
XU$$3683 t$6286 net1327 VGND VGND VPWR VPWR booth_b52_m57 sky130_fd_sc_hd__xor2_1
XU$$3694 net1537 net477 net1529 net750 VGND VGND VPWR VPWR t$6292 sky130_fd_sc_hd__a22o_1
XU$$2960 t$5917 net1371 VGND VGND VPWR VPWR booth_b42_m38 sky130_fd_sc_hd__xor2_1
XU$$2971 net1731 net521 net1722 net794 VGND VGND VPWR VPWR t$5923 sky130_fd_sc_hd__a22o_1
XU$$2982 t$5928 net1374 VGND VGND VPWR VPWR booth_b42_m49 sky130_fd_sc_hd__xor2_1
XU$$2993 net1626 net524 net1618 net797 VGND VGND VPWR VPWR t$5934 sky130_fd_sc_hd__a22o_1
XFILLER_33_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_691 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1988_ clknet_leaf_38_clk booth_b14_m41 VGND VGND VPWR VPWR pp_row55_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_165_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0939_ clknet_leaf_114_clk booth_b64_m33 VGND VGND VPWR VPWR pp_row97_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$900 final_adder.$signal$1212 final_adder.g_new$969 final_adder.$signal$246
+ VGND VGND VPWR VPWR final_adder.g_new$1028 sky130_fd_sc_hd__a21o_1
Xdadda_ha_1_37_1 pp_row37_3 pp_row37_4 VGND VGND VPWR VPWR c$214 s$215 sky130_fd_sc_hd__ha_1
XFILLER_102_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$911 final_adder.$signal$1190 final_adder.g_new$991 final_adder.$signal$202
+ VGND VGND VPWR VPWR final_adder.g_new$1039 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$922 final_adder.$signal$1168 final_adder.g_new$1013 final_adder.$signal$158
+ VGND VGND VPWR VPWR final_adder.g_new$1050 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$933 final_adder.$signal$1146 final_adder.g_new$939 final_adder.$signal$114
+ VGND VGND VPWR VPWR final_adder.g_new$1061 sky130_fd_sc_hd__a21o_1
Xdadda_fa_1_50_1 pp_row50_3 pp_row50_4 pp_row50_5 VGND VGND VPWR VPWR c$350 s$351
+ sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$944 final_adder.$signal$1124 final_adder.g_new$961 final_adder.$signal$70
+ VGND VGND VPWR VPWR final_adder.g_new$1072 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$955 final_adder.$signal$1102 final_adder.g_new$751 final_adder.$signal$26
+ VGND VGND VPWR VPWR final_adder.g_new$1083 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$966 final_adder.$signal$1095 final_adder.g_new$1087 VGND VGND VPWR
+ VPWR net340 sky130_fd_sc_hd__xor2_1
XU$$805 net1607 net407 net1599 net673 VGND VGND VPWR VPWR t$4816 sky130_fd_sc_hd__a22o_1
XFILLER_21_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$816 t$4821 net1418 VGND VGND VPWR VPWR booth_b10_m62 sky130_fd_sc_hd__xor2_1
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$977 final_adder.$signal$1106 final_adder.g_new$747 VGND VGND VPWR
+ VPWR net292 sky130_fd_sc_hd__xor2_2
XU$$827 net4 net1417 VGND VGND VPWR VPWR sel_1$4828 sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_43_0 pp_row43_0 pp_row43_1 pp_row43_2 VGND VGND VPWR VPWR c$254 s$255
+ sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$988 final_adder.$signal$1117 final_adder.g_new$1076 VGND VGND VPWR
+ VPWR net304 sky130_fd_sc_hd__xor2_2
XU$$838 net1672 net394 net1561 net660 VGND VGND VPWR VPWR t$4834 sky130_fd_sc_hd__a22o_1
XFILLER_83_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$999 final_adder.$signal$1128 final_adder.g_new$957 VGND VGND VPWR
+ VPWR net316 sky130_fd_sc_hd__xor2_2
XFILLER_71_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$849 t$4839 net1312 VGND VGND VPWR VPWR booth_b12_m10 sky130_fd_sc_hd__xor2_1
XFILLER_189_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_72_2 c$1588 s$1591 s$1593 VGND VGND VPWR VPWR c$2418 s$2419 sky130_fd_sc_hd__fa_1
XFILLER_106_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1100 net1101 VGND VGND VPWR VPWR net1100 sky130_fd_sc_hd__clkbuf_8
XFILLER_79_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1111 net1113 VGND VGND VPWR VPWR net1111 sky130_fd_sc_hd__buf_4
Xdadda_fa_3_65_1 c$1498 c$1500 c$1502 VGND VGND VPWR VPWR c$2360 s$2361 sky130_fd_sc_hd__fa_1
XFILLER_152_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1122 net1124 VGND VGND VPWR VPWR net1122 sky130_fd_sc_hd__buf_4
XFILLER_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1133 net1134 VGND VGND VPWR VPWR net1133 sky130_fd_sc_hd__buf_4
Xfanout1144 net1145 VGND VGND VPWR VPWR net1144 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_6_42_0 c$3560 c$3562 s$3565 VGND VGND VPWR VPWR c$3980 s$3981 sky130_fd_sc_hd__fa_1
XFILLER_66_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_58_0 s$509 c$1410 c$1412 VGND VGND VPWR VPWR c$2302 s$2303 sky130_fd_sc_hd__fa_1
Xfanout1155 net1158 VGND VGND VPWR VPWR net1155 sky130_fd_sc_hd__buf_4
Xfanout1166 net1167 VGND VGND VPWR VPWR net1166 sky130_fd_sc_hd__buf_4
Xfanout1177 net1182 VGND VGND VPWR VPWR net1177 sky130_fd_sc_hd__buf_4
Xfanout1188 net1189 VGND VGND VPWR VPWR net1188 sky130_fd_sc_hd__buf_6
Xfanout1199 net1200 VGND VGND VPWR VPWR net1199 sky130_fd_sc_hd__clkbuf_4
XFILLER_93_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2201 t$5530 net1432 VGND VGND VPWR VPWR booth_b32_m1 sky130_fd_sc_hd__xor2_1
XU$$2212 net1521 net569 net1513 net842 VGND VGND VPWR VPWR t$5536 sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_101_2 s$2649 s$2651 s$2653 VGND VGND VPWR VPWR c$3300 s$3301 sky130_fd_sc_hd__fa_1
XFILLER_35_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2223 t$5541 net1430 VGND VGND VPWR VPWR booth_b32_m12 sky130_fd_sc_hd__xor2_1
XU$$2234 net1150 net571 net1144 net844 VGND VGND VPWR VPWR t$5547 sky130_fd_sc_hd__a22o_1
XU$$2245 t$5552 net1433 VGND VGND VPWR VPWR booth_b32_m23 sky130_fd_sc_hd__xor2_1
XU$$1500 net1544 net633 net1536 net906 VGND VGND VPWR VPWR t$5171 sky130_fd_sc_hd__a22o_1
XU$$1511 notblock$5175\[2\] net15 net1491 t$5176 notblock$5175\[0\] VGND VGND VPWR
+ VPWR sel_0$5177 sky130_fd_sc_hd__a32o_4
XU$$2256 net1050 net572 net1042 net845 VGND VGND VPWR VPWR t$5558 sky130_fd_sc_hd__a22o_1
XU$$2267 t$5563 net1433 VGND VGND VPWR VPWR booth_b32_m34 sky130_fd_sc_hd__xor2_1
XU$$1522 t$5183 net1475 VGND VGND VPWR VPWR booth_b22_m4 sky130_fd_sc_hd__xor2_1
XU$$2278 net941 net570 net925 net843 VGND VGND VPWR VPWR t$5569 sky130_fd_sc_hd__a22o_1
XU$$1533 net1497 net613 net1221 net886 VGND VGND VPWR VPWR t$5189 sky130_fd_sc_hd__a22o_1
XFILLER_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1544 t$5194 net1478 VGND VGND VPWR VPWR booth_b22_m15 sky130_fd_sc_hd__xor2_1
XFILLER_15_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2289 t$5574 net1434 VGND VGND VPWR VPWR booth_b32_m45 sky130_fd_sc_hd__xor2_1
XU$$1555 net1114 net610 net1105 net883 VGND VGND VPWR VPWR t$5200 sky130_fd_sc_hd__a22o_1
XU$$1566 t$5205 net1477 VGND VGND VPWR VPWR booth_b22_m26 sky130_fd_sc_hd__xor2_1
Xdadda_ha_3_116_0 net1918 pp_row116_1 VGND VGND VPWR VPWR c$2748 s$2749 sky130_fd_sc_hd__ha_1
X_1911_ clknet_leaf_70_clk booth_b50_m2 VGND VGND VPWR VPWR pp_row52_25 sky130_fd_sc_hd__dfxtp_1
XU$$1577 net1018 net614 net1001 net887 VGND VGND VPWR VPWR t$5211 sky130_fd_sc_hd__a22o_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1588 t$5216 net1480 VGND VGND VPWR VPWR booth_b22_m37 sky130_fd_sc_hd__xor2_1
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1599 net1741 net615 net1733 net888 VGND VGND VPWR VPWR t$5222 sky130_fd_sc_hd__a22o_1
XFILLER_176_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1842_ clknet_leaf_62_clk booth_b34_m16 VGND VGND VPWR VPWR pp_row50_17 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_7_115_0 s$3859 c$4124 s$4127 VGND VGND VPWR VPWR c$4382 s$4383 sky130_fd_sc_hd__fa_1
XFILLER_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1773_ clknet_leaf_238_clk booth_b16_m32 VGND VGND VPWR VPWR pp_row48_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_8_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0724_ clknet_leaf_135_clk booth_b30_m58 VGND VGND VPWR VPWR pp_row88_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_183_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0655_ clknet_leaf_131_clk booth_b58_m59 VGND VGND VPWR VPWR pp_row117_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_131_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0586_ clknet_leaf_194_clk net237 VGND VGND VPWR VPWR pp_row82_25 sky130_fd_sc_hd__dfxtp_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2325_ clknet_leaf_74_clk booth_b52_m12 VGND VGND VPWR VPWR pp_row64_26 sky130_fd_sc_hd__dfxtp_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_2_60_0 s$49 c$510 c$512 VGND VGND VPWR VPWR c$1446 s$1447 sky130_fd_sc_hd__fa_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$207 final_adder.$signal$101 final_adder.$signal$98 final_adder.$signal$100
+ VGND VGND VPWR VPWR final_adder.g_new$335 sky130_fd_sc_hd__a21o_1
XFILLER_85_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$218 final_adder.$signal$1126 final_adder.$signal$1127 VGND VGND VPWR
+ VPWR final_adder.p_new$346 sky130_fd_sc_hd__and2_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$229 final_adder.$signal$1117 final_adder.$signal$54 final_adder.$signal$56
+ VGND VGND VPWR VPWR final_adder.g_new$357 sky130_fd_sc_hd__a21o_1
X_2256_ clknet_leaf_149_clk booth_b62_m0 VGND VGND VPWR VPWR pp_row62_31 sky130_fd_sc_hd__dfxtp_1
XFILLER_100_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1207_ clknet_leaf_47_clk booth_b12_m10 VGND VGND VPWR VPWR pp_row22_6 sky130_fd_sc_hd__dfxtp_1
X_2187_ clknet_leaf_227_clk booth_b0_m61 VGND VGND VPWR VPWR pp_row61_0 sky130_fd_sc_hd__dfxtp_1
XU$$4170 net1069 net435 net1061 net717 VGND VGND VPWR VPWR t$6536 sky130_fd_sc_hd__a22o_1
XU$$4181 t$6541 net1269 VGND VGND VPWR VPWR booth_b60_m32 sky130_fd_sc_hd__xor2_1
XFILLER_65_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4192 net962 net440 net953 net722 VGND VGND VPWR VPWR t$6547 sky130_fd_sc_hd__a22o_1
X_1138_ clknet_leaf_119_clk booth_b62_m40 VGND VGND VPWR VPWR pp_row102_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_92_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3480 t$6183 net1329 VGND VGND VPWR VPWR booth_b50_m24 sky130_fd_sc_hd__xor2_1
XU$$3491 net1043 net486 net1027 net759 VGND VGND VPWR VPWR t$6189 sky130_fd_sc_hd__a22o_1
XFILLER_41_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1069_ clknet_leaf_51_clk booth_b4_m6 VGND VGND VPWR VPWR pp_row10_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_129_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2790 net1110 net536 net1099 net809 VGND VGND VPWR VPWR t$5831 sky130_fd_sc_hd__a22o_1
XFILLER_193_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_82_1 c$2490 c$2492 s$2495 VGND VGND VPWR VPWR c$3184 s$3185 sky130_fd_sc_hd__fa_1
XFILLER_190_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_75_0 s$1637 c$2430 c$2432 VGND VGND VPWR VPWR c$3140 s$3141 sky130_fd_sc_hd__fa_1
XFILLER_134_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput203 c[51] VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_1
Xinput214 c[61] VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__clkbuf_1
Xinput225 c[71] VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__clkbuf_1
Xinput236 c[81] VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__clkbuf_1
Xinput247 c[91] VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$741 final_adder.p_new$756 final_adder.g_new$789 final_adder.g_new$757
+ VGND VGND VPWR VPWR final_adder.g_new$869 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$752 final_adder.p_new$800 final_adder.p_new$768 VGND VGND VPWR VPWR
+ final_adder.p_new$880 sky130_fd_sc_hd__and2_1
XFILLER_5_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$763 final_adder.p_new$778 final_adder.g_new$811 final_adder.g_new$779
+ VGND VGND VPWR VPWR final_adder.g_new$891 sky130_fd_sc_hd__a21o_1
XU$$602 net1089 net410 net1081 net676 VGND VGND VPWR VPWR t$4713 sky130_fd_sc_hd__a22o_1
XFILLER_44_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$613 t$4718 net1241 VGND VGND VPWR VPWR booth_b8_m29 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$774 final_adder.p_new$822 final_adder.p_new$790 VGND VGND VPWR VPWR
+ final_adder.p_new$902 sky130_fd_sc_hd__and2_1
XFILLER_57_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$785 final_adder.p_new$800 final_adder.g_new$833 final_adder.g_new$801
+ VGND VGND VPWR VPWR final_adder.g_new$913 sky130_fd_sc_hd__a21o_1
XU$$624 net982 net409 net973 net675 VGND VGND VPWR VPWR t$4724 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$796 final_adder.p_new$844 final_adder.p_new$812 VGND VGND VPWR VPWR
+ final_adder.p_new$924 sky130_fd_sc_hd__and2_1
XU$$635 t$4729 net1237 VGND VGND VPWR VPWR booth_b8_m40 sky130_fd_sc_hd__xor2_1
XU$$646 net1716 net414 net1707 net680 VGND VGND VPWR VPWR t$4735 sky130_fd_sc_hd__a22o_1
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$657 t$4740 net1238 VGND VGND VPWR VPWR booth_b8_m51 sky130_fd_sc_hd__xor2_1
XFILLER_189_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$668 net1607 net417 net1599 net683 VGND VGND VPWR VPWR t$4746 sky130_fd_sc_hd__a22o_1
XFILLER_182_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_876 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$679 t$4751 net1242 VGND VGND VPWR VPWR booth_b8_m62 sky130_fd_sc_hd__xor2_1
XFILLER_44_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0440_ clknet_leaf_161_clk booth_b64_m13 VGND VGND VPWR VPWR pp_row77_26 sky130_fd_sc_hd__dfxtp_1
XFILLER_79_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0371_ clknet_leaf_203_clk booth_b52_m23 VGND VGND VPWR VPWR pp_row75_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_67_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2110_ clknet_leaf_86_clk booth_b54_m4 VGND VGND VPWR VPWR pp_row58_27 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4387_1812 VGND VGND VPWR VPWR U$$4387_1812/HI net1812 sky130_fd_sc_hd__conb_1
XFILLER_181_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2041_ clknet_leaf_82_clk booth_b52_m4 VGND VGND VPWR VPWR pp_row56_26 sky130_fd_sc_hd__dfxtp_1
XFILLER_82_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2020 net1695 net589 net1687 net862 VGND VGND VPWR VPWR t$5437 sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_32_4 pp_row32_12 pp_row32_13 pp_row32_14 VGND VGND VPWR VPWR c$1118 s$1119
+ sky130_fd_sc_hd__fa_1
XU$$2031 t$5442 net1453 VGND VGND VPWR VPWR booth_b28_m53 sky130_fd_sc_hd__xor2_1
XU$$2042 net1588 net589 net1579 net862 VGND VGND VPWR VPWR t$5448 sky130_fd_sc_hd__a22o_1
XFILLER_62_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2053 t$5453 net1455 VGND VGND VPWR VPWR booth_b28_m64 sky130_fd_sc_hd__xor2_1
XU$$2064 t$5460 net1439 VGND VGND VPWR VPWR booth_b30_m1 sky130_fd_sc_hd__xor2_1
XU$$1330 t$5084 net1669 VGND VGND VPWR VPWR booth_b18_m45 sky130_fd_sc_hd__xor2_1
XU$$2075 net1521 net581 net1515 net854 VGND VGND VPWR VPWR t$5466 sky130_fd_sc_hd__a22o_1
XU$$2086 t$5471 net1439 VGND VGND VPWR VPWR booth_b30_m12 sky130_fd_sc_hd__xor2_1
XU$$1341 net1657 net642 net1649 net915 VGND VGND VPWR VPWR t$5090 sky130_fd_sc_hd__a22o_1
XU$$1352 t$5095 net1669 VGND VGND VPWR VPWR booth_b18_m56 sky130_fd_sc_hd__xor2_1
XU$$2097 net1148 net576 net1140 net849 VGND VGND VPWR VPWR t$5477 sky130_fd_sc_hd__a22o_1
XU$$1363 net1544 net641 net1536 net914 VGND VGND VPWR VPWR t$5101 sky130_fd_sc_hd__a22o_1
XU$$1374 notblock$5105\[2\] net13 net1668 t$5106 notblock$5105\[0\] VGND VGND VPWR
+ VPWR sel_0$5107 sky130_fd_sc_hd__a32o_2
XFILLER_149_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1385 t$5113 net1485 VGND VGND VPWR VPWR booth_b20_m4 sky130_fd_sc_hd__xor2_1
XFILLER_176_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1396 net1494 net627 net1219 net900 VGND VGND VPWR VPWR t$5119 sky130_fd_sc_hd__a22o_1
X_1825_ clknet_leaf_234_clk booth_b6_m44 VGND VGND VPWR VPWR pp_row50_3 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_92_0 c$3236 c$3238 c$3240 VGND VGND VPWR VPWR c$3764 s$3765 sky130_fd_sc_hd__fa_1
X_1756_ clknet_leaf_239_clk booth_b36_m11 VGND VGND VPWR VPWR pp_row47_18 sky130_fd_sc_hd__dfxtp_1
X_0707_ clknet_leaf_167_clk booth_b46_m41 VGND VGND VPWR VPWR pp_row87_12 sky130_fd_sc_hd__dfxtp_1
X_1687_ clknet_leaf_25_clk booth_b12_m33 VGND VGND VPWR VPWR pp_row45_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_144_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0638_ clknet_leaf_188_clk booth_b60_m24 VGND VGND VPWR VPWR pp_row84_21 sky130_fd_sc_hd__dfxtp_1
Xfanout904 sel_1$5108 VGND VGND VPWR VPWR net904 sky130_fd_sc_hd__buf_4
Xfanout915 sel_1$5038 VGND VGND VPWR VPWR net915 sky130_fd_sc_hd__buf_6
XFILLER_131_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout926 net931 VGND VGND VPWR VPWR net926 sky130_fd_sc_hd__clkbuf_8
Xdadda_fa_1_77_6 pp_row77_21 pp_row77_22 pp_row77_23 VGND VGND VPWR VPWR c$846 s$847
+ sky130_fd_sc_hd__fa_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout937 net939 VGND VGND VPWR VPWR net937 sky130_fd_sc_hd__clkbuf_4
Xfanout948 net949 VGND VGND VPWR VPWR net948 sky130_fd_sc_hd__buf_4
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0569_ clknet_leaf_188_clk booth_b34_m48 VGND VGND VPWR VPWR pp_row82_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_98_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout959 net960 VGND VGND VPWR VPWR net959 sky130_fd_sc_hd__buf_6
XTAP_4009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_892 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2308_ clknet_leaf_90_clk booth_b20_m44 VGND VGND VPWR VPWR pp_row64_10 sky130_fd_sc_hd__dfxtp_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2239_ clknet_leaf_230_clk booth_b30_m32 VGND VGND VPWR VPWR pp_row62_15 sky130_fd_sc_hd__dfxtp_1
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_308 net450 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_319 net592 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$70 c$4290 s$4293 VGND VGND VPWR VPWR final_adder.$signal$142 final_adder.$signal$1160
+ sky130_fd_sc_hd__ha_1
XFILLER_0_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$81 c$4312 s$4315 VGND VGND VPWR VPWR final_adder.$signal$164 final_adder.$signal$1171
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$92 c$4334 s$4337 VGND VGND VPWR VPWR final_adder.$signal$186 final_adder.$signal$1182
+ sky130_fd_sc_hd__ha_1
XFILLER_179_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_101_1 pp_row101_15 c$1924 c$1926 VGND VGND VPWR VPWR c$2648 s$2649 sky130_fd_sc_hd__fa_1
XFILLER_102_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_122_0 c$3880 c$3882 s$3885 VGND VGND VPWR VPWR c$4140 s$4141 sky130_fd_sc_hd__fa_1
Xdadda_fa_0_65_4 pp_row65_12 pp_row65_13 pp_row65_14 VGND VGND VPWR VPWR c$104 s$105
+ sky130_fd_sc_hd__fa_1
XFILLER_36_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_42_3 s$1235 s$1237 s$1239 VGND VGND VPWR VPWR c$2180 s$2181 sky130_fd_sc_hd__fa_1
XTAP_3820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$560 final_adder.p_new$572 final_adder.p_new$564 VGND VGND VPWR VPWR
+ final_adder.p_new$688 sky130_fd_sc_hd__and2_1
XTAP_3842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$410 net1280 VGND VGND VPWR VPWR notsign$4614 sky130_fd_sc_hd__inv_1
Xfinal_adder.U$$571 final_adder.p_new$574 final_adder.g_new$583 final_adder.g_new$575
+ VGND VGND VPWR VPWR final_adder.g_new$699 sky130_fd_sc_hd__a21o_1
XTAP_3853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$421 net1127 net430 net1035 net712 VGND VGND VPWR VPWR t$4621 sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_35_2 c$1144 s$1147 s$1149 VGND VGND VPWR VPWR c$2122 s$2123 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$582 final_adder.p_new$594 final_adder.p_new$586 VGND VGND VPWR VPWR
+ final_adder.p_new$710 sky130_fd_sc_hd__and2_1
XTAP_3864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$593 final_adder.p_new$596 final_adder.g_new$605 final_adder.g_new$597
+ VGND VGND VPWR VPWR final_adder.g_new$721 sky130_fd_sc_hd__a21o_1
XU$$432 t$4626 net1248 VGND VGND VPWR VPWR booth_b6_m7 sky130_fd_sc_hd__xor2_1
XFILLER_45_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$443 net1206 net431 net1198 net713 VGND VGND VPWR VPWR t$4632 sky130_fd_sc_hd__a22o_1
XTAP_3886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$454 t$4637 net1245 VGND VGND VPWR VPWR booth_b6_m18 sky130_fd_sc_hd__xor2_1
XTAP_3897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$465 net1088 net426 net1080 net708 VGND VGND VPWR VPWR t$4643 sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_28_1 pp_row28_14 pp_row28_15 pp_row28_16 VGND VGND VPWR VPWR c$2064 s$2065
+ sky130_fd_sc_hd__fa_2
XFILLER_60_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$476 t$4648 net1249 VGND VGND VPWR VPWR booth_b6_m29 sky130_fd_sc_hd__xor2_1
XFILLER_32_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$487 net982 net426 net973 net708 VGND VGND VPWR VPWR t$4654 sky130_fd_sc_hd__a22o_1
XU$$498 t$4659 net1244 VGND VGND VPWR VPWR booth_b6_m40 sky130_fd_sc_hd__xor2_1
XFILLER_44_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_992 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1610_ clknet_leaf_239_clk booth_b18_m24 VGND VGND VPWR VPWR pp_row42_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_154_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1541_ clknet_leaf_8_clk booth_b24_m15 VGND VGND VPWR VPWR pp_row39_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_141_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_87_5 s$993 s$995 s$997 VGND VGND VPWR VPWR c$1780 s$1781 sky130_fd_sc_hd__fa_2
XFILLER_113_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1472_ clknet_leaf_110_clk booth_b64_m40 VGND VGND VPWR VPWR pp_row104_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_140_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0423_ clknet_leaf_207_clk booth_b32_m45 VGND VGND VPWR VPWR pp_row77_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_79_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0354_ clknet_leaf_196_clk booth_b22_m53 VGND VGND VPWR VPWR pp_row75_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_83_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0285_ clknet_leaf_202_clk booth_b12_m61 VGND VGND VPWR VPWR pp_row73_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_82_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2024_ clknet_leaf_35_clk booth_b22_m34 VGND VGND VPWR VPWR pp_row56_11 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_30_1 pp_row30_3 pp_row30_4 pp_row30_5 VGND VGND VPWR VPWR c$1092 s$1093
+ sky130_fd_sc_hd__fa_1
XFILLER_47_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1160 net1047 net644 net1039 net917 VGND VGND VPWR VPWR t$4998 sky130_fd_sc_hd__a22o_1
XU$$1171 t$5003 net1010 VGND VGND VPWR VPWR booth_b16_m34 sky130_fd_sc_hd__xor2_1
XFILLER_149_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1182 net944 net645 net928 net918 VGND VGND VPWR VPWR t$5009 sky130_fd_sc_hd__a22o_1
XFILLER_10_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1193 t$5014 net1007 VGND VGND VPWR VPWR booth_b16_m45 sky130_fd_sc_hd__xor2_1
XFILLER_137_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_117_1 s$3393 s$3395 s$3397 VGND VGND VPWR VPWR c$3866 s$3867 sky130_fd_sc_hd__fa_2
XFILLER_40_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1808_ clknet_leaf_24_clk booth_b26_m23 VGND VGND VPWR VPWR pp_row49_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_145_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1739_ clknet_leaf_122_clk booth_b58_m48 VGND VGND VPWR VPWR pp_row106_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_172_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_82_4 pp_row82_12 pp_row82_13 pp_row82_14 VGND VGND VPWR VPWR c$930 s$931
+ sky130_fd_sc_hd__fa_1
Xfanout701 net703 VGND VGND VPWR VPWR net701 sky130_fd_sc_hd__buf_4
XFILLER_131_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout712 net713 VGND VGND VPWR VPWR net712 sky130_fd_sc_hd__buf_4
Xfanout723 sel_1$6508 VGND VGND VPWR VPWR net723 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_1_75_3 pp_row75_15 pp_row75_16 pp_row75_17 VGND VGND VPWR VPWR c$804 s$805
+ sky130_fd_sc_hd__fa_1
Xfanout734 sel_1$6368 VGND VGND VPWR VPWR net734 sky130_fd_sc_hd__clkbuf_4
XFILLER_131_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout745 net748 VGND VGND VPWR VPWR net745 sky130_fd_sc_hd__buf_6
Xdadda_fa_4_52_2 s$2257 s$2259 s$2261 VGND VGND VPWR VPWR c$3006 s$3007 sky130_fd_sc_hd__fa_1
Xfanout756 sel_1$6228 VGND VGND VPWR VPWR net756 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_68_2 pp_row68_23 pp_row68_24 pp_row68_25 VGND VGND VPWR VPWR c$676 s$677
+ sky130_fd_sc_hd__fa_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout767 net768 VGND VGND VPWR VPWR net767 sky130_fd_sc_hd__buf_4
XFILLER_86_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout778 net779 VGND VGND VPWR VPWR net778 sky130_fd_sc_hd__buf_4
XFILLER_100_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout789 net790 VGND VGND VPWR VPWR net789 sky130_fd_sc_hd__buf_4
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_45_1 c$2194 c$2196 s$2199 VGND VGND VPWR VPWR c$2962 s$2963 sky130_fd_sc_hd__fa_1
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_22_0 s$3487 c$3938 s$3941 VGND VGND VPWR VPWR c$4196 s$4197 sky130_fd_sc_hd__fa_1
XTAP_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_38_0 s$1193 c$2134 c$2136 VGND VGND VPWR VPWR c$2918 s$2919 sky130_fd_sc_hd__fa_1
XTAP_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_105 net581 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_116 net644 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_127 net683 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 net740 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_149 net791 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_748 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_0_57_2 pp_row57_6 pp_row57_7 VGND VGND VPWR VPWR c$22 s$23 sky130_fd_sc_hd__ha_1
XFILLER_190_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_0_70_2 pp_row70_6 pp_row70_7 pp_row70_8 VGND VGND VPWR VPWR c$158 s$159
+ sky130_fd_sc_hd__fa_1
XFILLER_49_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_0_63_1 pp_row63_3 pp_row63_4 pp_row63_5 VGND VGND VPWR VPWR c$74 s$75 sky130_fd_sc_hd__fa_1
XFILLER_76_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_938 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_40_0 s$235 c$1194 c$1196 VGND VGND VPWR VPWR c$2158 s$2159 sky130_fd_sc_hd__fa_1
XTAP_4362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_56_0 pp_row56_0 pp_row56_1 pp_row56_2 VGND VGND VPWR VPWR c$12 s$13 sky130_fd_sc_hd__fa_1
XTAP_4373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$390 final_adder.p_new$396 final_adder.p_new$392 VGND VGND VPWR VPWR
+ final_adder.p_new$518 sky130_fd_sc_hd__and2_1
XFILLER_18_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$240 t$4527 net1387 VGND VGND VPWR VPWR booth_b2_m48 sky130_fd_sc_hd__xor2_1
XTAP_3683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$251 net1633 sel_0$4477 net1623 sel_1$4478 VGND VGND VPWR VPWR t$4533 sky130_fd_sc_hd__a22o_1
XFILLER_189_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$262 t$4538 net1387 VGND VGND VPWR VPWR booth_b2_m59 sky130_fd_sc_hd__xor2_1
XFILLER_17_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$273 net1393 VGND VGND VPWR VPWR notsign$4544 sky130_fd_sc_hd__inv_1
XU$$284 net1128 net534 net1035 net807 VGND VGND VPWR VPWR t$4551 sky130_fd_sc_hd__a22o_1
XTAP_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$295 t$4556 net1277 VGND VGND VPWR VPWR booth_b4_m7 sky130_fd_sc_hd__xor2_1
XTAP_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0972_ clknet_leaf_117_clk booth_b54_m45 VGND VGND VPWR VPWR pp_row99_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_158_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1 net1 VGND VGND VPWR VPWR notblock\[1\] sky130_fd_sc_hd__inv_1
XFILLER_145_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$9 c$4168 s$4171 VGND VGND VPWR VPWR final_adder.$signal$20 final_adder.$signal$1099
+ sky130_fd_sc_hd__ha_1
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput304 net304 VGND VGND VPWR VPWR o[27] sky130_fd_sc_hd__buf_2
XFILLER_161_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_92_3 pp_row92_17 pp_row92_18 pp_row92_19 VGND VGND VPWR VPWR c$1836 s$1837
+ sky130_fd_sc_hd__fa_1
Xoutput315 net315 VGND VGND VPWR VPWR o[37] sky130_fd_sc_hd__buf_2
XFILLER_99_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput326 net326 VGND VGND VPWR VPWR o[47] sky130_fd_sc_hd__buf_2
Xoutput337 net337 VGND VGND VPWR VPWR o[57] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_85_2 c$952 c$954 c$956 VGND VGND VPWR VPWR c$1750 s$1751 sky130_fd_sc_hd__fa_1
XFILLER_142_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput348 net348 VGND VGND VPWR VPWR o[67] sky130_fd_sc_hd__buf_2
X_1524_ clknet_leaf_242_clk booth_b38_m0 VGND VGND VPWR VPWR pp_row38_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_113_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput359 net359 VGND VGND VPWR VPWR o[77] sky130_fd_sc_hd__buf_2
Xdadda_fa_5_62_1 s$3063 s$3065 s$3067 VGND VGND VPWR VPWR c$3646 s$3647 sky130_fd_sc_hd__fa_1
Xdadda_fa_2_78_1 c$838 c$840 c$842 VGND VGND VPWR VPWR c$1664 s$1665 sky130_fd_sc_hd__fa_1
XFILLER_87_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1455_ clknet_leaf_40_clk booth_b34_m1 VGND VGND VPWR VPWR pp_row35_17 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_55_0 c$3014 c$3016 c$3018 VGND VGND VPWR VPWR c$3616 s$3617 sky130_fd_sc_hd__fa_1
XFILLER_171_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0406_ clknet_leaf_206_clk booth_b58_m18 VGND VGND VPWR VPWR pp_row76_24 sky130_fd_sc_hd__dfxtp_1
X_1386_ clknet_leaf_42_clk booth_b26_m6 VGND VGND VPWR VPWR pp_row32_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_67_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_54_8 pp_row54_29 c$2 s$5 VGND VGND VPWR VPWR c$436 s$437 sky130_fd_sc_hd__fa_1
X_0337_ clknet_leaf_226_clk booth_b48_m26 VGND VGND VPWR VPWR pp_row74_20 sky130_fd_sc_hd__dfxtp_1
XFILLER_67_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0268_ clknet_leaf_209_clk booth_b42_m30 VGND VGND VPWR VPWR pp_row72_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_71_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2007_ clknet_leaf_72_clk booth_b48_m7 VGND VGND VPWR VPWR pp_row55_24 sky130_fd_sc_hd__dfxtp_1
XFILLER_70_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_101_0 pp_row101_0 pp_row101_1 pp_row101_2 VGND VGND VPWR VPWR c$1934 s$1935
+ sky130_fd_sc_hd__fa_1
X_0199_ clknet_leaf_153_clk booth_b40_m30 VGND VGND VPWR VPWR pp_row70_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_50_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4107_1804 VGND VGND VPWR VPWR U$$4107_1804/HI net1804 sky130_fd_sc_hd__conb_1
XFILLER_91_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_80_1 pp_row80_3 pp_row80_4 pp_row80_5 VGND VGND VPWR VPWR c$890 s$891
+ sky130_fd_sc_hd__fa_1
Xfanout1507 net127 VGND VGND VPWR VPWR net1507 sky130_fd_sc_hd__buf_6
XFILLER_132_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_73_0 pp_row73_9 pp_row73_10 pp_row73_11 VGND VGND VPWR VPWR c$762 s$763
+ sky130_fd_sc_hd__fa_1
Xfanout520 sel_0$5877 VGND VGND VPWR VPWR net520 sky130_fd_sc_hd__buf_4
Xfanout1518 net126 VGND VGND VPWR VPWR net1518 sky130_fd_sc_hd__buf_8
Xfanout1529 net1530 VGND VGND VPWR VPWR net1529 sky130_fd_sc_hd__buf_2
XFILLER_99_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout531 net532 VGND VGND VPWR VPWR net531 sky130_fd_sc_hd__buf_4
Xfanout542 sel_0$5807 VGND VGND VPWR VPWR net542 sky130_fd_sc_hd__buf_8
Xfanout553 net559 VGND VGND VPWR VPWR net553 sky130_fd_sc_hd__buf_4
XFILLER_150_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout564 net568 VGND VGND VPWR VPWR net564 sky130_fd_sc_hd__buf_4
Xfanout575 sel_0$5527 VGND VGND VPWR VPWR net575 sky130_fd_sc_hd__buf_6
XFILLER_24_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout586 net592 VGND VGND VPWR VPWR net586 sky130_fd_sc_hd__buf_4
Xfanout597 net601 VGND VGND VPWR VPWR net597 sky130_fd_sc_hd__buf_6
XFILLER_47_938 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3309 t$6096 net1343 VGND VGND VPWR VPWR booth_b48_m7 sky130_fd_sc_hd__xor2_1
XFILLER_18_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2608 net32 net1411 VGND VGND VPWR VPWR sel_1$5738 sky130_fd_sc_hd__xor2_1
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2619 net1673 net543 net1562 net816 VGND VGND VPWR VPWR t$5744 sky130_fd_sc_hd__a22o_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1907 net1579 net599 net1553 net872 VGND VGND VPWR VPWR t$5379 sky130_fd_sc_hd__a22o_1
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1918 net1463 VGND VGND VPWR VPWR notblock$5385\[0\] sky130_fd_sc_hd__inv_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1929 t$5391 net1448 VGND VGND VPWR VPWR booth_b28_m2 sky130_fd_sc_hd__xor2_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_130_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_130_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_183_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_95_1 c$1858 c$1860 c$1862 VGND VGND VPWR VPWR c$2600 s$2601 sky130_fd_sc_hd__fa_2
XFILLER_6_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_72_0 c$3680 c$3682 s$3685 VGND VGND VPWR VPWR c$4040 s$4041 sky130_fd_sc_hd__fa_1
Xdadda_fa_3_88_0 s$1009 c$1770 c$1772 VGND VGND VPWR VPWR c$2542 s$2543 sky130_fd_sc_hd__fa_1
XFILLER_170_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1240_ clknet_leaf_13_clk booth_b18_m6 VGND VGND VPWR VPWR pp_row24_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_1_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4500 net1625 sel_0$6647 net1617 net699 VGND VGND VPWR VPWR t$6704 sky130_fd_sc_hd__a22o_1
XU$$4511 t$6709 net1876 VGND VGND VPWR VPWR booth_b64_m60 sky130_fd_sc_hd__xor2_1
XFILLER_65_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_197_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_197_clk
+ sky130_fd_sc_hd__clkbuf_16
X_1171_ clknet_leaf_125_clk notsign$5804 VGND VGND VPWR VPWR pp_row103_0 sky130_fd_sc_hd__dfxtp_1
XU$$14 net937 net447 net1675 net689 VGND VGND VPWR VPWR t$4414 sky130_fd_sc_hd__a22o_1
XU$$25 t$4419 net1573 VGND VGND VPWR VPWR booth_b0_m9 sky130_fd_sc_hd__xor2_1
XU$$3810 t$6351 net1306 VGND VGND VPWR VPWR booth_b54_m52 sky130_fd_sc_hd__xor2_1
XFILLER_49_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_117_0 pp_row117_0 pp_row117_1 pp_row117_2 VGND VGND VPWR VPWR c$3392 s$3393
+ sky130_fd_sc_hd__fa_1
XU$$3821 net1600 net473 net1591 net746 VGND VGND VPWR VPWR t$6357 sky130_fd_sc_hd__a22o_1
XTAP_4170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$36 net1175 net443 net1166 net685 VGND VGND VPWR VPWR t$4425 sky130_fd_sc_hd__a22o_1
XU$$3832 t$6362 net1302 VGND VGND VPWR VPWR booth_b54_m63 sky130_fd_sc_hd__xor2_1
XTAP_4181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$47 t$4430 net1575 VGND VGND VPWR VPWR booth_b0_m20 sky130_fd_sc_hd__xor2_1
XTAP_4192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$58 net1071 net442 net1063 net684 VGND VGND VPWR VPWR t$4436 sky130_fd_sc_hd__a22o_1
XU$$3843 t$6369 net1296 VGND VGND VPWR VPWR booth_b56_m0 sky130_fd_sc_hd__xor2_1
XU$$69 t$4441 net1568 VGND VGND VPWR VPWR booth_b0_m31 sky130_fd_sc_hd__xor2_1
XU$$3854 net1563 net461 net1522 net734 VGND VGND VPWR VPWR t$6375 sky130_fd_sc_hd__a22o_1
XU$$3865 t$6380 net1296 VGND VGND VPWR VPWR booth_b56_m11 sky130_fd_sc_hd__xor2_1
Xdadda_ha_5_4_0 pp_row4_0 pp_row4_1 VGND VGND VPWR VPWR c$3416 s$3417 sky130_fd_sc_hd__ha_1
XU$$3876 net1159 net460 net1151 net733 VGND VGND VPWR VPWR t$6386 sky130_fd_sc_hd__a22o_1
XTAP_3480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3887 t$6391 net1291 VGND VGND VPWR VPWR booth_b56_m22 sky130_fd_sc_hd__xor2_1
XTAP_3491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3898 net1061 net463 net1052 net736 VGND VGND VPWR VPWR t$6397 sky130_fd_sc_hd__a22o_1
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_16 sel_0$4477 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_27 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_38 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_49 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0955_ clknet_leaf_131_clk booth_b60_m61 VGND VGND VPWR VPWR pp_row121_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_186_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_121_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_121_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_146_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0886_ clknet_leaf_100_clk booth_b40_m55 VGND VGND VPWR VPWR pp_row95_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_173_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_90_0 pp_row90_11 pp_row90_12 pp_row90_13 VGND VGND VPWR VPWR c$1806 s$1807
+ sky130_fd_sc_hd__fa_1
XFILLER_161_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1507_ clknet_leaf_16_clk booth_b6_m32 VGND VGND VPWR VPWR pp_row38_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_141_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2487_ clknet_leaf_90_clk booth_b16_m53 VGND VGND VPWR VPWR pp_row69_6 sky130_fd_sc_hd__dfxtp_1
Xdadda_ha_1_46_6 pp_row46_18 pp_row46_19 VGND VGND VPWR VPWR c$300 s$301 sky130_fd_sc_hd__ha_1
XFILLER_114_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1438_ clknet_leaf_55_clk booth_b4_m31 VGND VGND VPWR VPWR pp_row35_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_130_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_188_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_188_clk
+ sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_1_52_5 pp_row52_17 pp_row52_18 pp_row52_19 VGND VGND VPWR VPWR c$394 s$395
+ sky130_fd_sc_hd__fa_1
X_1369_ clknet_leaf_4_clk booth_b30_m1 VGND VGND VPWR VPWR pp_row31_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_56_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_45_4 pp_row45_12 pp_row45_13 pp_row45_14 VGND VGND VPWR VPWR c$284 s$285
+ sky130_fd_sc_hd__fa_1
XFILLER_110_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_15_2 pp_row15_8 c$1974 s$1977 VGND VGND VPWR VPWR c$2784 s$2785 sky130_fd_sc_hd__fa_1
XFILLER_169_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$1008 final_adder.$signal$1137 final_adder.g_new$1066 VGND VGND VPWR
+ VPWR net326 sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$1019 final_adder.$signal$1148 final_adder.g_new$937 VGND VGND VPWR
+ VPWR net338 sky130_fd_sc_hd__xor2_2
XFILLER_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_112_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_112_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_165_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_913 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1304 net1305 VGND VGND VPWR VPWR net1304 sky130_fd_sc_hd__clkbuf_8
Xfanout1315 net5 VGND VGND VPWR VPWR net1315 sky130_fd_sc_hd__buf_4
Xfanout1326 net1327 VGND VGND VPWR VPWR net1326 sky130_fd_sc_hd__buf_6
XFILLER_8_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1337 net47 VGND VGND VPWR VPWR net1337 sky130_fd_sc_hd__buf_6
Xfanout1348 net1349 VGND VGND VPWR VPWR net1348 sky130_fd_sc_hd__buf_6
XFILLER_121_979 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1359 net1361 VGND VGND VPWR VPWR net1359 sky130_fd_sc_hd__buf_6
XFILLER_93_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_179_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_179_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_120_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout394 net400 VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__buf_6
XU$$3106 net1740 net512 net1732 net785 VGND VGND VPWR VPWR t$5992 sky130_fd_sc_hd__a22o_1
XFILLER_86_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3117 t$5997 net1364 VGND VGND VPWR VPWR booth_b44_m48 sky130_fd_sc_hd__xor2_1
XFILLER_4_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3128 net1635 net516 net1626 net789 VGND VGND VPWR VPWR t$6003 sky130_fd_sc_hd__a22o_1
XU$$3139 t$6008 net1360 VGND VGND VPWR VPWR booth_b44_m59 sky130_fd_sc_hd__xor2_1
XU$$2405 net988 net567 net979 net840 VGND VGND VPWR VPWR t$5634 sky130_fd_sc_hd__a22o_1
XFILLER_98_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2416 t$5639 net1422 VGND VGND VPWR VPWR booth_b34_m40 sky130_fd_sc_hd__xor2_1
XU$$2427 net1713 net565 net1704 net838 VGND VGND VPWR VPWR t$5645 sky130_fd_sc_hd__a22o_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2438 t$5650 net1427 VGND VGND VPWR VPWR booth_b34_m51 sky130_fd_sc_hd__xor2_1
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1704 net1066 net605 net1057 net878 VGND VGND VPWR VPWR t$5276 sky130_fd_sc_hd__a22o_1
XU$$2449 net1608 net567 net1600 net840 VGND VGND VPWR VPWR t$5656 sky130_fd_sc_hd__a22o_1
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1715 t$5281 net1470 VGND VGND VPWR VPWR booth_b24_m32 sky130_fd_sc_hd__xor2_1
XFILLER_27_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1726 net957 net604 net948 net877 VGND VGND VPWR VPWR t$5287 sky130_fd_sc_hd__a22o_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1737 t$5292 net1474 VGND VGND VPWR VPWR booth_b24_m43 sky130_fd_sc_hd__xor2_1
XU$$1748 net1687 net607 net1679 net880 VGND VGND VPWR VPWR t$5298 sky130_fd_sc_hd__a22o_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1759 t$5303 net1473 VGND VGND VPWR VPWR booth_b24_m54 sky130_fd_sc_hd__xor2_1
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput14 a[21] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_4
XFILLER_174_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput25 a[31] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_103_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_103_clk
+ sky130_fd_sc_hd__clkbuf_16
Xinput36 a[41] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
X_0740_ clknet_leaf_163_clk booth_b60_m28 VGND VGND VPWR VPWR pp_row88_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_7_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput47 a[51] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_2
Xinput58 a[61] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_4
Xinput69 b[13] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_4
XFILLER_155_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0671_ clknet_leaf_175_clk booth_b26_m60 VGND VGND VPWR VPWR pp_row86_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_7_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2410_ clknet_leaf_84_clk booth_b4_m63 VGND VGND VPWR VPWR pp_row67_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_143_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2341_ clknet_leaf_89_clk booth_b14_m51 VGND VGND VPWR VPWR pp_row65_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2272_ clknet_leaf_210_clk booth_b22_m41 VGND VGND VPWR VPWR pp_row63_11 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_62_4 s$569 s$571 s$573 VGND VGND VPWR VPWR c$1478 s$1479 sky130_fd_sc_hd__fa_1
XFILLER_78_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_819 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1223_ clknet_leaf_48_clk booth_b14_m9 VGND VGND VPWR VPWR pp_row23_7 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_55_3 c$436 s$439 s$441 VGND VGND VPWR VPWR c$1392 s$1393 sky130_fd_sc_hd__fa_1
XFILLER_84_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4330 t$6617 net1261 VGND VGND VPWR VPWR booth_b62_m38 sky130_fd_sc_hd__xor2_1
XFILLER_65_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4341 net1731 net419 net1722 net701 VGND VGND VPWR VPWR t$6623 sky130_fd_sc_hd__a22o_1
XFILLER_77_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_48_2 c$306 c$308 c$310 VGND VGND VPWR VPWR c$1306 s$1307 sky130_fd_sc_hd__fa_1
XU$$4352 t$6628 net1260 VGND VGND VPWR VPWR booth_b62_m49 sky130_fd_sc_hd__xor2_1
X_1154_ clknet_leaf_47_clk booth_b14_m4 VGND VGND VPWR VPWR pp_row18_7 sky130_fd_sc_hd__dfxtp_1
XU$$4363 net1628 net420 net1617 net702 VGND VGND VPWR VPWR t$6634 sky130_fd_sc_hd__a22o_1
XU$$4374 t$6639 net1261 VGND VGND VPWR VPWR booth_b62_m60 sky130_fd_sc_hd__xor2_1
XFILLER_92_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3640 net979 net478 net970 net751 VGND VGND VPWR VPWR t$6265 sky130_fd_sc_hd__a22o_1
XU$$4385 net1810 VGND VGND VPWR VPWR notblock$6645\[1\] sky130_fd_sc_hd__inv_1
XU$$4396 net1038 sel_0$6647 net939 net698 VGND VGND VPWR VPWR t$6652 sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_25_1 s$2841 s$2843 s$2845 VGND VGND VPWR VPWR c$3498 s$3499 sky130_fd_sc_hd__fa_2
XU$$3651 t$6270 net1322 VGND VGND VPWR VPWR booth_b52_m41 sky130_fd_sc_hd__xor2_1
XFILLER_37_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_587 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3662 net1708 net482 net1700 net755 VGND VGND VPWR VPWR t$6276 sky130_fd_sc_hd__a22o_1
XU$$3673 t$6281 net1326 VGND VGND VPWR VPWR booth_b52_m52 sky130_fd_sc_hd__xor2_1
X_1085_ clknet_leaf_58_clk booth_b2_m10 VGND VGND VPWR VPWR pp_row12_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_18_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_18_0 c$2792 c$2794 c$2796 VGND VGND VPWR VPWR c$3468 s$3469 sky130_fd_sc_hd__fa_1
XU$$3684 net1600 net483 net1591 net756 VGND VGND VPWR VPWR t$6287 sky130_fd_sc_hd__a22o_1
XU$$2950 t$5912 net1370 VGND VGND VPWR VPWR booth_b42_m33 sky130_fd_sc_hd__xor2_1
XU$$3695 t$6292 net1321 VGND VGND VPWR VPWR booth_b52_m63 sky130_fd_sc_hd__xor2_1
XFILLER_34_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2961 net951 net521 net943 net794 VGND VGND VPWR VPWR t$5918 sky130_fd_sc_hd__a22o_1
XU$$2972 t$5923 net1369 VGND VGND VPWR VPWR booth_b42_m44 sky130_fd_sc_hd__xor2_1
XFILLER_34_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2983 net1684 net524 net1660 net797 VGND VGND VPWR VPWR t$5929 sky130_fd_sc_hd__a22o_1
XU$$2994 t$5934 net1373 VGND VGND VPWR VPWR booth_b42_m55 sky130_fd_sc_hd__xor2_1
XFILLER_33_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1987_ clknet_leaf_81_clk booth_b12_m43 VGND VGND VPWR VPWR pp_row55_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_193_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0938_ clknet_leaf_113_clk booth_b62_m35 VGND VGND VPWR VPWR pp_row97_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_180_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0869_ clknet_leaf_104_clk booth_b46_m48 VGND VGND VPWR VPWR pp_row94_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_134_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$901 final_adder.$signal$1210 final_adder.g_new$971 final_adder.$signal$242
+ VGND VGND VPWR VPWR final_adder.g_new$1029 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$912 final_adder.$signal$1188 final_adder.g_new$993 final_adder.$signal$198
+ VGND VGND VPWR VPWR final_adder.g_new$1040 sky130_fd_sc_hd__a21o_1
XFILLER_102_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$923 final_adder.$signal$1166 final_adder.g_new$1015 final_adder.$signal$154
+ VGND VGND VPWR VPWR final_adder.g_new$1051 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$934 final_adder.$signal$111 final_adder.g_new$941 final_adder.$signal$110
+ VGND VGND VPWR VPWR final_adder.g_new$1062 sky130_fd_sc_hd__a21o_1
XFILLER_68_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_50_2 pp_row50_6 pp_row50_7 pp_row50_8 VGND VGND VPWR VPWR c$352 s$353
+ sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$945 final_adder.$signal$1122 final_adder.g_new$851 final_adder.$signal$66
+ VGND VGND VPWR VPWR final_adder.g_new$1073 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$956 final_adder.$signal$1100 final_adder.g_new$753 final_adder.$signal$22
+ VGND VGND VPWR VPWR final_adder.g_new$1084 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$967 final_adder.$signal$1096 final_adder.g_new$633 VGND VGND VPWR
+ VPWR net351 sky130_fd_sc_hd__xor2_2
XU$$806 t$4816 net1419 VGND VGND VPWR VPWR booth_b10_m57 sky130_fd_sc_hd__xor2_1
XU$$817 net1535 net403 net1527 net669 VGND VGND VPWR VPWR t$4822 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$978 final_adder.$signal$1107 final_adder.g_new$1081 VGND VGND VPWR
+ VPWR net293 sky130_fd_sc_hd__xor2_2
Xdadda_fa_1_43_1 pp_row43_3 pp_row43_4 pp_row43_5 VGND VGND VPWR VPWR c$256 s$257
+ sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$989 final_adder.$signal$1118 final_adder.g_new$855 VGND VGND VPWR
+ VPWR net305 sky130_fd_sc_hd__xor2_2
XU$$828 net1887 net397 net1231 net663 VGND VGND VPWR VPWR t$4829 sky130_fd_sc_hd__a22o_1
XU$$839 t$4834 net1310 VGND VGND VPWR VPWR booth_b12_m5 sky130_fd_sc_hd__xor2_1
XFILLER_56_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_20_0 pp_row20_11 pp_row20_12 c$1992 VGND VGND VPWR VPWR c$2810 s$2811
+ sky130_fd_sc_hd__fa_1
XFILLER_189_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1082 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_36_0 pp_row36_0 pp_row36_1 pp_row36_2 VGND VGND VPWR VPWR c$208 s$209
+ sky130_fd_sc_hd__fa_1
XFILLER_188_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_72_3 s$1595 s$1597 s$1599 VGND VGND VPWR VPWR c$2420 s$2421 sky130_fd_sc_hd__fa_1
XFILLER_191_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1101 net79 VGND VGND VPWR VPWR net1101 sky130_fd_sc_hd__buf_6
XFILLER_78_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1112 net1113 VGND VGND VPWR VPWR net1112 sky130_fd_sc_hd__buf_4
Xdadda_fa_3_65_2 c$1504 s$1507 s$1509 VGND VGND VPWR VPWR c$2362 s$2363 sky130_fd_sc_hd__fa_1
XFILLER_79_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1123 net1124 VGND VGND VPWR VPWR net1123 sky130_fd_sc_hd__buf_4
Xfanout1134 net75 VGND VGND VPWR VPWR net1134 sky130_fd_sc_hd__buf_4
Xfanout1145 net74 VGND VGND VPWR VPWR net1145 sky130_fd_sc_hd__buf_4
XFILLER_113_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1156 net1158 VGND VGND VPWR VPWR net1156 sky130_fd_sc_hd__buf_2
Xdadda_fa_3_58_1 c$1414 c$1416 c$1418 VGND VGND VPWR VPWR c$2304 s$2305 sky130_fd_sc_hd__fa_1
Xfanout1167 net71 VGND VGND VPWR VPWR net1167 sky130_fd_sc_hd__buf_4
Xfanout1178 net1182 VGND VGND VPWR VPWR net1178 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_6_35_0 c$3532 c$3534 s$3537 VGND VGND VPWR VPWR c$3966 s$3967 sky130_fd_sc_hd__fa_1
Xfanout1189 net1190 VGND VGND VPWR VPWR net1189 sky130_fd_sc_hd__clkbuf_4
XFILLER_75_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2202 net1128 net572 net1035 net845 VGND VGND VPWR VPWR t$5531 sky130_fd_sc_hd__a22o_1
XFILLER_170_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2213 t$5536 net1430 VGND VGND VPWR VPWR booth_b32_m7 sky130_fd_sc_hd__xor2_1
XU$$2224 net1203 net570 net1194 net843 VGND VGND VPWR VPWR t$5542 sky130_fd_sc_hd__a22o_1
XU$$2235 t$5547 net1432 VGND VGND VPWR VPWR booth_b32_m18 sky130_fd_sc_hd__xor2_1
XFILLER_28_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2246 net1092 net572 net1084 net845 VGND VGND VPWR VPWR t$5553 sky130_fd_sc_hd__a22o_1
XU$$1501 t$5171 net1491 VGND VGND VPWR VPWR booth_b20_m62 sky130_fd_sc_hd__xor2_1
XU$$1512 net15 net1491 VGND VGND VPWR VPWR sel_1$5178 sky130_fd_sc_hd__xor2_4
XU$$2257 t$5558 net1433 VGND VGND VPWR VPWR booth_b32_m29 sky130_fd_sc_hd__xor2_1
XU$$2268 net989 net572 net978 net845 VGND VGND VPWR VPWR t$5564 sky130_fd_sc_hd__a22o_1
XU$$1523 net1671 net610 net1560 net883 VGND VGND VPWR VPWR t$5184 sky130_fd_sc_hd__a22o_1
XFILLER_37_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2279 t$5569 net1431 VGND VGND VPWR VPWR booth_b32_m40 sky130_fd_sc_hd__xor2_1
XU$$1534 t$5189 net1478 VGND VGND VPWR VPWR booth_b22_m10 sky130_fd_sc_hd__xor2_1
XFILLER_31_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1545 net1166 net613 net1157 net886 VGND VGND VPWR VPWR t$5195 sky130_fd_sc_hd__a22o_1
XU$$1556 t$5200 net1475 VGND VGND VPWR VPWR booth_b22_m21 sky130_fd_sc_hd__xor2_1
X_1910_ clknet_leaf_70_clk booth_b48_m4 VGND VGND VPWR VPWR pp_row52_24 sky130_fd_sc_hd__dfxtp_1
XFILLER_163_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1567 net1064 net612 net1056 net885 VGND VGND VPWR VPWR t$5206 sky130_fd_sc_hd__a22o_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1578 t$5211 net1479 VGND VGND VPWR VPWR booth_b22_m32 sky130_fd_sc_hd__xor2_1
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1589 net957 net612 net949 net885 VGND VGND VPWR VPWR t$5217 sky130_fd_sc_hd__a22o_1
XFILLER_179_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1841_ clknet_leaf_62_clk booth_b32_m18 VGND VGND VPWR VPWR pp_row50_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1772_ clknet_leaf_187_clk booth_b64_m42 VGND VGND VPWR VPWR pp_row106_12 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_7_108_0 s$3831 c$4110 s$4113 VGND VGND VPWR VPWR c$4368 s$4369 sky130_fd_sc_hd__fa_1
XFILLER_144_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0723_ clknet_leaf_135_clk booth_b28_m60 VGND VGND VPWR VPWR pp_row88_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_116_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0654_ clknet_leaf_169_clk booth_b42_m43 VGND VGND VPWR VPWR pp_row85_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_170_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0585_ clknet_leaf_188_clk booth_b64_m18 VGND VGND VPWR VPWR pp_row82_24 sky130_fd_sc_hd__dfxtp_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2324_ clknet_leaf_74_clk booth_b50_m14 VGND VGND VPWR VPWR pp_row64_25 sky130_fd_sc_hd__dfxtp_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_2_60_1 c$514 c$516 c$518 VGND VGND VPWR VPWR c$1448 s$1449 sky130_fd_sc_hd__fa_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_84_0_1898 VGND VGND VPWR VPWR net1898 dadda_fa_1_84_0_1898/LO sky130_fd_sc_hd__conb_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$208 final_adder.$signal$1136 final_adder.$signal$1137 VGND VGND VPWR
+ VPWR final_adder.p_new$336 sky130_fd_sc_hd__and2_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2255_ clknet_leaf_149_clk booth_b60_m2 VGND VGND VPWR VPWR pp_row62_30 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$219 final_adder.$signal$1127 final_adder.$signal$74 final_adder.$signal$76
+ VGND VGND VPWR VPWR final_adder.g_new$347 sky130_fd_sc_hd__a21o_1
Xdadda_fa_2_53_0 s$3 c$384 c$386 VGND VGND VPWR VPWR c$1362 s$1363 sky130_fd_sc_hd__fa_1
XFILLER_84_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1206_ clknet_leaf_47_clk booth_b10_m12 VGND VGND VPWR VPWR pp_row22_5 sky130_fd_sc_hd__dfxtp_1
Xfanout1690 net107 VGND VGND VPWR VPWR net1690 sky130_fd_sc_hd__buf_4
XFILLER_38_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2186_ clknet_leaf_231_clk net213 VGND VGND VPWR VPWR pp_row60_32 sky130_fd_sc_hd__dfxtp_1
XU$$4160 net1112 net436 net1103 net718 VGND VGND VPWR VPWR t$6531 sky130_fd_sc_hd__a22o_1
XU$$4171 t$6536 net1266 VGND VGND VPWR VPWR booth_b60_m27 sky130_fd_sc_hd__xor2_1
XU$$4182 net1004 net437 net996 net719 VGND VGND VPWR VPWR t$6542 sky130_fd_sc_hd__a22o_1
XU$$4193 t$6547 net1271 VGND VGND VPWR VPWR booth_b60_m38 sky130_fd_sc_hd__xor2_1
X_1137_ clknet_leaf_16_clk booth_b4_m13 VGND VGND VPWR VPWR pp_row17_2 sky130_fd_sc_hd__dfxtp_1
XU$$3470 t$6178 net1333 VGND VGND VPWR VPWR booth_b50_m19 sky130_fd_sc_hd__xor2_1
XFILLER_20_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3481 net1086 net485 net1076 net758 VGND VGND VPWR VPWR t$6184 sky130_fd_sc_hd__a22o_1
XFILLER_80_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3492 t$6189 net1330 VGND VGND VPWR VPWR booth_b50_m30 sky130_fd_sc_hd__xor2_1
XFILLER_80_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1068_ clknet_leaf_51_clk booth_b2_m8 VGND VGND VPWR VPWR pp_row10_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_7_0 pp_row7_0 pp_row7_1 pp_row7_2 VGND VGND VPWR VPWR c$3424 s$3425 sky130_fd_sc_hd__fa_1
XU$$2780 net1161 net542 net1150 net815 VGND VGND VPWR VPWR t$5826 sky130_fd_sc_hd__a22o_1
XU$$2791 t$5831 net1377 VGND VGND VPWR VPWR booth_b40_m22 sky130_fd_sc_hd__xor2_1
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_908 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_82_2 s$2497 s$2499 s$2501 VGND VGND VPWR VPWR c$3186 s$3187 sky130_fd_sc_hd__fa_1
XU$$1787_1767 VGND VGND VPWR VPWR U$$1787_1767/HI net1767 sky130_fd_sc_hd__conb_1
Xdadda_fa_4_75_1 c$2434 c$2436 s$2439 VGND VGND VPWR VPWR c$3142 s$3143 sky130_fd_sc_hd__fa_1
XFILLER_68_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_52_0 s$3607 c$3998 s$4001 VGND VGND VPWR VPWR c$4256 s$4257 sky130_fd_sc_hd__fa_1
XFILLER_191_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_68_0 s$1553 c$2374 c$2376 VGND VGND VPWR VPWR c$3098 s$3099 sky130_fd_sc_hd__fa_1
Xinput204 c[52] VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_1
Xinput215 c[62] VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput226 c[72] VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__clkbuf_1
Xinput237 c[82] VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput248 c[92] VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__clkbuf_1
Xfinal_adder.U$$720 final_adder.p_new$744 final_adder.p_new$728 VGND VGND VPWR VPWR
+ final_adder.p_new$848 sky130_fd_sc_hd__and2_1
XFILLER_29_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$731 final_adder.p_new$738 final_adder.g_new$631 final_adder.g_new$739
+ VGND VGND VPWR VPWR final_adder.g_new$859 sky130_fd_sc_hd__a21o_2
Xfinal_adder.U$$742 final_adder.p_new$790 final_adder.p_new$758 VGND VGND VPWR VPWR
+ final_adder.p_new$870 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$753 final_adder.p_new$768 final_adder.g_new$801 final_adder.g_new$769
+ VGND VGND VPWR VPWR final_adder.g_new$881 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$764 final_adder.p_new$812 final_adder.p_new$780 VGND VGND VPWR VPWR
+ final_adder.p_new$892 sky130_fd_sc_hd__and2_1
XU$$603 t$4713 net1236 VGND VGND VPWR VPWR booth_b8_m24 sky130_fd_sc_hd__xor2_1
XU$$614 net1040 net410 net1024 net676 VGND VGND VPWR VPWR t$4719 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$775 final_adder.p_new$790 final_adder.g_new$823 final_adder.g_new$791
+ VGND VGND VPWR VPWR final_adder.g_new$903 sky130_fd_sc_hd__a21o_1
XFILLER_17_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$625 t$4724 net1235 VGND VGND VPWR VPWR booth_b8_m35 sky130_fd_sc_hd__xor2_1
XFILLER_72_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$786 final_adder.p_new$834 final_adder.p_new$802 VGND VGND VPWR VPWR
+ final_adder.p_new$914 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$797 final_adder.p_new$812 final_adder.g_new$845 final_adder.g_new$813
+ VGND VGND VPWR VPWR final_adder.g_new$925 sky130_fd_sc_hd__a21o_1
XU$$636 net925 net412 net1746 net678 VGND VGND VPWR VPWR t$4730 sky130_fd_sc_hd__a22o_1
XU$$647 t$4735 net1241 VGND VGND VPWR VPWR booth_b8_m46 sky130_fd_sc_hd__xor2_1
XU$$658 net1648 net411 net1640 net677 VGND VGND VPWR VPWR t$4741 sky130_fd_sc_hd__a22o_1
XU$$669 t$4746 net1242 VGND VGND VPWR VPWR booth_b8_m57 sky130_fd_sc_hd__xor2_1
XFILLER_140_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2746_1782 VGND VGND VPWR VPWR U$$2746_1782/HI net1782 sky130_fd_sc_hd__conb_1
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_70_0 s$725 c$1554 c$1556 VGND VGND VPWR VPWR c$2398 s$2399 sky130_fd_sc_hd__fa_1
XFILLER_152_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0370_ clknet_leaf_205_clk booth_b50_m25 VGND VGND VPWR VPWR pp_row75_20 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_0_72_0_1893 VGND VGND VPWR VPWR net1893 dadda_fa_0_72_0_1893/LO sky130_fd_sc_hd__conb_1
XFILLER_121_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2040_ clknet_leaf_83_clk booth_b50_m6 VGND VGND VPWR VPWR pp_row56_25 sky130_fd_sc_hd__dfxtp_1
XFILLER_181_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2010 net1738 net589 net1730 net862 VGND VGND VPWR VPWR t$5432 sky130_fd_sc_hd__a22o_1
XU$$2021 t$5437 net1454 VGND VGND VPWR VPWR booth_b28_m48 sky130_fd_sc_hd__xor2_1
XU$$2032 net1631 net590 net1622 net863 VGND VGND VPWR VPWR t$5443 sky130_fd_sc_hd__a22o_1
XU$$2043 t$5448 net1453 VGND VGND VPWR VPWR booth_b28_m59 sky130_fd_sc_hd__xor2_1
XU$$2054 net1455 VGND VGND VPWR VPWR notsign$5454 sky130_fd_sc_hd__inv_1
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2065 net1126 net581 net1032 net854 VGND VGND VPWR VPWR t$5461 sky130_fd_sc_hd__a22o_1
XU$$1320 t$5079 net1666 VGND VGND VPWR VPWR booth_b18_m40 sky130_fd_sc_hd__xor2_1
XU$$1331 net1715 net642 net1706 net915 VGND VGND VPWR VPWR t$5085 sky130_fd_sc_hd__a22o_1
XU$$2076 t$5466 net1441 VGND VGND VPWR VPWR booth_b30_m7 sky130_fd_sc_hd__xor2_1
XU$$2087 net1201 net576 net1192 net849 VGND VGND VPWR VPWR t$5472 sky130_fd_sc_hd__a22o_1
XU$$1342 t$5090 net1670 VGND VGND VPWR VPWR booth_b18_m51 sky130_fd_sc_hd__xor2_1
XU$$1353 net1604 net640 net1595 net913 VGND VGND VPWR VPWR t$5096 sky130_fd_sc_hd__a22o_1
XU$$2098 t$5477 net1439 VGND VGND VPWR VPWR booth_b30_m18 sky130_fd_sc_hd__xor2_1
XFILLER_149_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1364 t$5101 net1670 VGND VGND VPWR VPWR booth_b18_m62 sky130_fd_sc_hd__xor2_1
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1375 net13 net1668 VGND VGND VPWR VPWR sel_1$5108 sky130_fd_sc_hd__xor2_4
XU$$1386 net1671 net628 net1560 net901 VGND VGND VPWR VPWR t$5114 sky130_fd_sc_hd__a22o_1
XU$$1397 t$5119 net1485 VGND VGND VPWR VPWR booth_b20_m10 sky130_fd_sc_hd__xor2_1
XFILLER_176_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_960 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1824_ clknet_leaf_234_clk booth_b4_m46 VGND VGND VPWR VPWR pp_row50_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_191_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_92_1 s$3243 s$3245 s$3247 VGND VGND VPWR VPWR c$3766 s$3767 sky130_fd_sc_hd__fa_1
XFILLER_163_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1755_ clknet_leaf_238_clk booth_b34_m13 VGND VGND VPWR VPWR pp_row47_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_8_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_790 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_85_0 c$3194 c$3196 c$3198 VGND VGND VPWR VPWR c$3736 s$3737 sky130_fd_sc_hd__fa_1
X_0706_ clknet_leaf_171_clk booth_b44_m43 VGND VGND VPWR VPWR pp_row87_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_116_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1686_ clknet_leaf_19_clk booth_b10_m35 VGND VGND VPWR VPWR pp_row45_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_143_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0637_ clknet_leaf_188_clk booth_b58_m26 VGND VGND VPWR VPWR pp_row84_20 sky130_fd_sc_hd__dfxtp_1
XFILLER_171_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout905 net907 VGND VGND VPWR VPWR net905 sky130_fd_sc_hd__buf_4
XFILLER_131_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout916 net917 VGND VGND VPWR VPWR net916 sky130_fd_sc_hd__buf_4
Xfanout927 net931 VGND VGND VPWR VPWR net927 sky130_fd_sc_hd__buf_4
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_77_7 pp_row77_24 pp_row77_25 pp_row77_26 VGND VGND VPWR VPWR c$848 s$849
+ sky130_fd_sc_hd__fa_1
XFILLER_174_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0568_ clknet_leaf_188_clk booth_b32_m50 VGND VGND VPWR VPWR pp_row82_8 sky130_fd_sc_hd__dfxtp_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout938 net939 VGND VGND VPWR VPWR net938 sky130_fd_sc_hd__buf_4
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout949 net952 VGND VGND VPWR VPWR net949 sky130_fd_sc_hd__buf_6
XFILLER_86_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2307_ clknet_leaf_91_clk booth_b18_m46 VGND VGND VPWR VPWR pp_row64_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_100_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0499_ clknet_leaf_126_clk booth_b62_m53 VGND VGND VPWR VPWR pp_row115_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_100_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2238_ clknet_leaf_136_clk booth_b52_m58 VGND VGND VPWR VPWR pp_row110_4 sky130_fd_sc_hd__dfxtp_1
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_309 net461 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2169_ clknet_leaf_215_clk booth_b36_m24 VGND VGND VPWR VPWR pp_row60_18 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_92_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_92_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$60 c$4270 s$4273 VGND VGND VPWR VPWR final_adder.$signal$122 final_adder.$signal$1150
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$71 c$4292 s$4295 VGND VGND VPWR VPWR final_adder.$signal$144 final_adder.$signal$1161
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$82 c$4314 s$4317 VGND VGND VPWR VPWR final_adder.$signal$166 final_adder.$signal$1172
+ sky130_fd_sc_hd__ha_1
XFILLER_80_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$93 c$4336 s$4339 VGND VGND VPWR VPWR final_adder.$signal$188 final_adder.$signal$1183
+ sky130_fd_sc_hd__ha_1
XFILLER_16_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_101_2 c$1928 c$1930 c$1932 VGND VGND VPWR VPWR c$2650 s$2651 sky130_fd_sc_hd__fa_1
XFILLER_190_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_0_65_5 pp_row65_15 pp_row65_16 pp_row65_17 VGND VGND VPWR VPWR c$106 s$107
+ sky130_fd_sc_hd__fa_2
Xdadda_fa_6_115_0 c$3852 c$3854 s$3857 VGND VGND VPWR VPWR c$4126 s$4127 sky130_fd_sc_hd__fa_1
XTAP_3810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$550 final_adder.p_new$562 final_adder.p_new$554 VGND VGND VPWR VPWR
+ final_adder.p_new$678 sky130_fd_sc_hd__and2_1
XTAP_3832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$561 final_adder.p_new$564 final_adder.g_new$573 final_adder.g_new$565
+ VGND VGND VPWR VPWR final_adder.g_new$689 sky130_fd_sc_hd__a21o_1
XU$$400 net1578 net529 net1551 net802 VGND VGND VPWR VPWR t$4609 sky130_fd_sc_hd__a22o_1
XFILLER_57_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$411 net1275 VGND VGND VPWR VPWR notblock$4615\[0\] sky130_fd_sc_hd__inv_1
Xfinal_adder.U$$572 final_adder.p_new$584 final_adder.p_new$576 VGND VGND VPWR VPWR
+ final_adder.p_new$700 sky130_fd_sc_hd__and2_1
XTAP_3854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$422 t$4621 net1248 VGND VGND VPWR VPWR booth_b6_m2 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$583 final_adder.p_new$586 final_adder.g_new$595 final_adder.g_new$587
+ VGND VGND VPWR VPWR final_adder.g_new$711 sky130_fd_sc_hd__a21o_1
Xdadda_fa_3_35_3 s$1151 s$1153 s$1155 VGND VGND VPWR VPWR c$2124 s$2125 sky130_fd_sc_hd__fa_1
XTAP_3865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$433 net1513 net431 net1505 net713 VGND VGND VPWR VPWR t$4627 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$594 final_adder.p_new$606 final_adder.p_new$598 VGND VGND VPWR VPWR
+ final_adder.p_new$722 sky130_fd_sc_hd__and2_1
XTAP_3876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$444 t$4632 net1250 VGND VGND VPWR VPWR booth_b6_m13 sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_83_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_83_clk sky130_fd_sc_hd__clkbuf_16
XTAP_3887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$455 net1139 net427 net1131 net709 VGND VGND VPWR VPWR t$4638 sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_28_2 c$1068 c$1070 c$1072 VGND VGND VPWR VPWR c$2066 s$2067 sky130_fd_sc_hd__fa_1
XTAP_3898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$466 t$4643 net1244 VGND VGND VPWR VPWR booth_b6_m24 sky130_fd_sc_hd__xor2_1
XFILLER_44_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$477 net1041 net431 net1025 net713 VGND VGND VPWR VPWR t$4649 sky130_fd_sc_hd__a22o_1
XFILLER_189_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$488 t$4654 net1244 VGND VGND VPWR VPWR booth_b6_m35 sky130_fd_sc_hd__xor2_1
XU$$499 net924 net426 net1745 net708 VGND VGND VPWR VPWR t$4660 sky130_fd_sc_hd__a22o_1
XFILLER_60_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1540_ clknet_leaf_12_clk booth_b22_m17 VGND VGND VPWR VPWR pp_row39_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_154_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1471_ clknet_leaf_39_clk booth_b26_m10 VGND VGND VPWR VPWR pp_row36_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_113_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0422_ clknet_leaf_181_clk net145 VGND VGND VPWR VPWR pp_row114_9 sky130_fd_sc_hd__dfxtp_2
XFILLER_68_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_ha_2_31_4 pp_row31_12 pp_row31_13 VGND VGND VPWR VPWR c$1108 s$1109 sky130_fd_sc_hd__ha_1
XFILLER_140_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0353_ clknet_leaf_200_clk booth_b20_m55 VGND VGND VPWR VPWR pp_row75_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_68_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0284_ clknet_leaf_202_clk booth_b10_m63 VGND VGND VPWR VPWR pp_row73_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_82_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_7_1_0 pp_row1_0 pp_row1_1 VGND VGND VPWR VPWR c$4154 s$4155 sky130_fd_sc_hd__ha_1
XFILLER_36_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2023_ clknet_leaf_34_clk booth_b20_m36 VGND VGND VPWR VPWR pp_row56_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_35_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_74_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_74_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_91_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_30_2 pp_row30_6 pp_row30_7 pp_row30_8 VGND VGND VPWR VPWR c$1094 s$1095
+ sky130_fd_sc_hd__fa_1
XFILLER_91_983 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1150 net1088 net643 net1080 net916 VGND VGND VPWR VPWR t$4993 sky130_fd_sc_hd__a22o_1
XFILLER_126_1019 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1161 t$4998 net1007 VGND VGND VPWR VPWR booth_b16_m29 sky130_fd_sc_hd__xor2_1
XU$$1172 net987 net647 net977 net920 VGND VGND VPWR VPWR t$5004 sky130_fd_sc_hd__a22o_1
XU$$1183 t$5009 net1011 VGND VGND VPWR VPWR booth_b16_m40 sky130_fd_sc_hd__xor2_1
XU$$1194 net1711 net648 net1703 net921 VGND VGND VPWR VPWR t$5015 sky130_fd_sc_hd__a22o_1
XFILLER_148_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1807_ clknet_leaf_24_clk booth_b24_m25 VGND VGND VPWR VPWR pp_row49_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1738_ clknet_leaf_236_clk booth_b4_m43 VGND VGND VPWR VPWR pp_row47_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_116_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_82_5 pp_row82_15 pp_row82_16 pp_row82_17 VGND VGND VPWR VPWR c$932 s$933
+ sky130_fd_sc_hd__fa_1
X_1669_ clknet_leaf_19_clk booth_b30_m14 VGND VGND VPWR VPWR pp_row44_15 sky130_fd_sc_hd__dfxtp_1
Xfanout702 net703 VGND VGND VPWR VPWR net702 sky130_fd_sc_hd__buf_4
XFILLER_160_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout713 net715 VGND VGND VPWR VPWR net713 sky130_fd_sc_hd__buf_4
XFILLER_172_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_75_4 pp_row75_18 pp_row75_19 pp_row75_20 VGND VGND VPWR VPWR c$806 s$807
+ sky130_fd_sc_hd__fa_1
Xfanout724 net732 VGND VGND VPWR VPWR net724 sky130_fd_sc_hd__buf_4
Xfanout735 net736 VGND VGND VPWR VPWR net735 sky130_fd_sc_hd__buf_4
Xfanout746 net748 VGND VGND VPWR VPWR net746 sky130_fd_sc_hd__buf_4
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout757 net760 VGND VGND VPWR VPWR net757 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_68_3 pp_row68_26 pp_row68_27 pp_row68_28 VGND VGND VPWR VPWR c$678 s$679
+ sky130_fd_sc_hd__fa_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout768 net769 VGND VGND VPWR VPWR net768 sky130_fd_sc_hd__clkbuf_8
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout779 net782 VGND VGND VPWR VPWR net779 sky130_fd_sc_hd__clkbuf_4
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_45_2 s$2201 s$2203 s$2205 VGND VGND VPWR VPWR c$2964 s$2965 sky130_fd_sc_hd__fa_1
XTAP_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_38_1 c$2138 c$2140 s$2143 VGND VGND VPWR VPWR c$2920 s$2921 sky130_fd_sc_hd__fa_1
XTAP_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_106 net581 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_65_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_65_clk sky130_fd_sc_hd__clkbuf_16
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_7_15_0 s$3459 c$3924 s$3927 VGND VGND VPWR VPWR c$4182 s$4183 sky130_fd_sc_hd__fa_1
XFILLER_54_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_117 net644 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_1102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_128 net703 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_139 net760 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_910 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2600_1778 VGND VGND VPWR VPWR U$$2600_1778/HI net1778 sky130_fd_sc_hd__conb_1
XFILLER_163_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_0_70_3 pp_row70_9 pp_row70_10 pp_row70_11 VGND VGND VPWR VPWR c$160 s$161
+ sky130_fd_sc_hd__fa_1
XFILLER_39_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_0_63_2 pp_row63_6 pp_row63_7 pp_row63_8 VGND VGND VPWR VPWR c$76 s$77 sky130_fd_sc_hd__fa_1
XTAP_4330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_40_1 c$1198 c$1200 c$1202 VGND VGND VPWR VPWR c$2160 s$2161 sky130_fd_sc_hd__fa_1
XTAP_4352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_56_1 pp_row56_3 pp_row56_4 pp_row56_5 VGND VGND VPWR VPWR c$14 s$15 sky130_fd_sc_hd__fa_1
XTAP_4374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_56_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_56_clk sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_3_33_0 pp_row33_17 c$1110 c$1112 VGND VGND VPWR VPWR c$2102 s$2103 sky130_fd_sc_hd__fa_2
XTAP_4396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$230 t$4522 net1388 VGND VGND VPWR VPWR booth_b2_m43 sky130_fd_sc_hd__xor2_1
XTAP_3662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$391 final_adder.p_new$392 final_adder.g_new$397 final_adder.g_new$393
+ VGND VGND VPWR VPWR final_adder.g_new$519 sky130_fd_sc_hd__a21o_1
XU$$241 net1691 net626 net1683 net899 VGND VGND VPWR VPWR t$4528 sky130_fd_sc_hd__a22o_1
XTAP_3673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$252 t$4533 net1393 VGND VGND VPWR VPWR booth_b2_m54 sky130_fd_sc_hd__xor2_1
XTAP_3695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$263 net1578 net621 net1551 net894 VGND VGND VPWR VPWR t$4539 sky130_fd_sc_hd__a22o_1
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$274 net1388 VGND VGND VPWR VPWR notblock$4545\[0\] sky130_fd_sc_hd__inv_1
XTAP_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$285 t$4551 net1277 VGND VGND VPWR VPWR booth_b4_m2 sky130_fd_sc_hd__xor2_1
XU$$296 net1516 net531 net1509 net804 VGND VGND VPWR VPWR t$4557 sky130_fd_sc_hd__a22o_1
XTAP_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0971_ clknet_leaf_117_clk booth_b52_m47 VGND VGND VPWR VPWR pp_row99_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_38_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2 net1571 VGND VGND VPWR VPWR notblock\[2\] sky130_fd_sc_hd__inv_1
XFILLER_69_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput305 net305 VGND VGND VPWR VPWR o[28] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_92_4 pp_row92_20 c$1026 c$1028 VGND VGND VPWR VPWR c$1838 s$1839 sky130_fd_sc_hd__fa_1
XFILLER_160_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput316 net316 VGND VGND VPWR VPWR o[38] sky130_fd_sc_hd__buf_2
Xoutput327 net327 VGND VGND VPWR VPWR o[48] sky130_fd_sc_hd__buf_2
XFILLER_114_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput338 net338 VGND VGND VPWR VPWR o[58] sky130_fd_sc_hd__buf_2
XFILLER_141_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput349 net349 VGND VGND VPWR VPWR o[68] sky130_fd_sc_hd__buf_2
X_1523_ clknet_leaf_242_clk booth_b36_m2 VGND VGND VPWR VPWR pp_row38_18 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_85_3 c$958 c$960 c$962 VGND VGND VPWR VPWR c$1752 s$1753 sky130_fd_sc_hd__fa_1
XFILLER_141_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1454_ clknet_leaf_64_clk booth_b32_m3 VGND VGND VPWR VPWR pp_row35_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_45_1020 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_78_2 c$844 c$846 c$848 VGND VGND VPWR VPWR c$1666 s$1667 sky130_fd_sc_hd__fa_1
XFILLER_141_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_55_1 s$3021 s$3023 s$3025 VGND VGND VPWR VPWR c$3618 s$3619 sky130_fd_sc_hd__fa_1
X_0405_ clknet_leaf_205_clk booth_b56_m20 VGND VGND VPWR VPWR pp_row76_23 sky130_fd_sc_hd__dfxtp_1
XFILLER_113_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1385_ clknet_leaf_42_clk booth_b24_m8 VGND VGND VPWR VPWR pp_row32_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_48_0 c$2972 c$2974 c$2976 VGND VGND VPWR VPWR c$3588 s$3589 sky130_fd_sc_hd__fa_1
X_0336_ clknet_leaf_225_clk booth_b46_m28 VGND VGND VPWR VPWR pp_row74_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_67_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_2_22_0 pp_row22_0 pp_row22_1 VGND VGND VPWR VPWR c$1050 s$1051 sky130_fd_sc_hd__ha_1
XFILLER_56_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0267_ clknet_leaf_209_clk booth_b40_m32 VGND VGND VPWR VPWR pp_row72_17 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_47_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_47_clk sky130_fd_sc_hd__clkbuf_16
X_2006_ clknet_leaf_72_clk booth_b46_m9 VGND VGND VPWR VPWR pp_row55_23 sky130_fd_sc_hd__dfxtp_1
X_0198_ clknet_leaf_153_clk booth_b38_m32 VGND VGND VPWR VPWR pp_row70_17 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_101_1 pp_row101_3 pp_row101_4 pp_row101_5 VGND VGND VPWR VPWR c$1936 s$1937
+ sky130_fd_sc_hd__fa_1
XFILLER_35_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_122_0 pp_row122_2 pp_row122_3 pp_row122_4 VGND VGND VPWR VPWR c$3884 s$3885
+ sky130_fd_sc_hd__fa_1
XFILLER_192_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_80_2 pp_row80_6 pp_row80_7 pp_row80_8 VGND VGND VPWR VPWR c$892 s$893
+ sky130_fd_sc_hd__fa_1
XFILLER_59_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout510 net518 VGND VGND VPWR VPWR net510 sky130_fd_sc_hd__buf_4
Xfanout1508 net1510 VGND VGND VPWR VPWR net1508 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_73_1 pp_row73_12 pp_row73_13 pp_row73_14 VGND VGND VPWR VPWR c$764 s$765
+ sky130_fd_sc_hd__fa_1
Xfanout521 net522 VGND VGND VPWR VPWR net521 sky130_fd_sc_hd__buf_4
Xfanout1519 net1521 VGND VGND VPWR VPWR net1519 sky130_fd_sc_hd__buf_4
Xfanout532 net534 VGND VGND VPWR VPWR net532 sky130_fd_sc_hd__buf_4
XFILLER_24_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout543 net544 VGND VGND VPWR VPWR net543 sky130_fd_sc_hd__buf_4
Xfanout554 net559 VGND VGND VPWR VPWR net554 sky130_fd_sc_hd__buf_4
Xdadda_fa_4_50_0 s$1337 c$2230 c$2232 VGND VGND VPWR VPWR c$2990 s$2991 sky130_fd_sc_hd__fa_1
Xfanout565 net568 VGND VGND VPWR VPWR net565 sky130_fd_sc_hd__clkbuf_8
Xdadda_fa_1_66_0 pp_row66_18 pp_row66_19 pp_row66_20 VGND VGND VPWR VPWR c$636 s$637
+ sky130_fd_sc_hd__fa_1
Xfanout576 net583 VGND VGND VPWR VPWR net576 sky130_fd_sc_hd__buf_4
XFILLER_19_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout587 net588 VGND VGND VPWR VPWR net587 sky130_fd_sc_hd__buf_4
Xfanout598 net600 VGND VGND VPWR VPWR net598 sky130_fd_sc_hd__buf_4
XFILLER_18_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2609 net1779 net543 net1227 net816 VGND VGND VPWR VPWR t$5739 sky130_fd_sc_hd__a22o_1
XFILLER_74_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_38_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_27_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1908 t$5379 net1463 VGND VGND VPWR VPWR booth_b26_m60 sky130_fd_sc_hd__xor2_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1919 net21 VGND VGND VPWR VPWR notblock$5385\[1\] sky130_fd_sc_hd__inv_1
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_791 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_95_2 c$1864 s$1867 s$1869 VGND VGND VPWR VPWR c$2602 s$2603 sky130_fd_sc_hd__fa_1
XFILLER_182_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_88_1 c$1774 c$1776 c$1778 VGND VGND VPWR VPWR c$2544 s$2545 sky130_fd_sc_hd__fa_2
XFILLER_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1513_1763 VGND VGND VPWR VPWR U$$1513_1763/HI net1763 sky130_fd_sc_hd__conb_1
Xdadda_fa_6_65_0 c$3652 c$3654 s$3657 VGND VGND VPWR VPWR c$4026 s$4027 sky130_fd_sc_hd__fa_2
XFILLER_124_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4501 t$6704 net1871 VGND VGND VPWR VPWR booth_b64_m55 sky130_fd_sc_hd__xor2_1
XU$$4512 net1553 sel_0$6647 net1544 net693 VGND VGND VPWR VPWR t$6710 sky130_fd_sc_hd__a22o_1
X_1170_ clknet_leaf_247_clk net167 VGND VGND VPWR VPWR pp_row19_10 sky130_fd_sc_hd__dfxtp_2
XU$$3800 t$6346 net1307 VGND VGND VPWR VPWR booth_b54_m47 sky130_fd_sc_hd__xor2_1
XFILLER_65_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$15 t$4414 net1573 VGND VGND VPWR VPWR booth_b0_m4 sky130_fd_sc_hd__xor2_1
XTAP_4160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3811 net1643 net470 net1634 net743 VGND VGND VPWR VPWR t$6352 sky130_fd_sc_hd__a22o_1
XU$$26 net1499 net446 net1224 net688 VGND VGND VPWR VPWR t$4420 sky130_fd_sc_hd__a22o_1
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$37 t$4425 net1568 VGND VGND VPWR VPWR booth_b0_m15 sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_117_1 pp_row117_3 pp_row117_4 pp_row117_5 VGND VGND VPWR VPWR c$3394 s$3395
+ sky130_fd_sc_hd__fa_1
XU$$3822 t$6357 net1306 VGND VGND VPWR VPWR booth_b54_m58 sky130_fd_sc_hd__xor2_1
XTAP_4171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_29_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_16
XU$$3833 net1533 net475 net1798 net748 VGND VGND VPWR VPWR t$6363 sky130_fd_sc_hd__a22o_1
XTAP_4182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$48 net1117 net448 net1108 net690 VGND VGND VPWR VPWR t$4431 sky130_fd_sc_hd__a22o_1
XU$$3844 net1233 net464 net1129 net737 VGND VGND VPWR VPWR t$6370 sky130_fd_sc_hd__a22o_1
XTAP_4193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$59 t$4436 net1568 VGND VGND VPWR VPWR booth_b0_m26 sky130_fd_sc_hd__xor2_1
XFILLER_64_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3855 t$6375 net1295 VGND VGND VPWR VPWR booth_b56_m6 sky130_fd_sc_hd__xor2_1
XFILLER_80_717 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3866 net1217 net464 net1208 net737 VGND VGND VPWR VPWR t$6381 sky130_fd_sc_hd__a22o_1
XTAP_3470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3877 t$6386 net1291 VGND VGND VPWR VPWR booth_b56_m17 sky130_fd_sc_hd__xor2_1
XTAP_3481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3888 net1102 net463 net1094 net736 VGND VGND VPWR VPWR t$6392 sky130_fd_sc_hd__a22o_1
XTAP_3492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3899 t$6397 net1294 VGND VGND VPWR VPWR booth_b56_m28 sky130_fd_sc_hd__xor2_1
XFILLER_33_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_17 sel_0$5107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_28 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_39 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0954_ clknet_leaf_116_clk booth_b56_m42 VGND VGND VPWR VPWR pp_row98_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_118_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0885_ clknet_leaf_100_clk booth_b38_m57 VGND VGND VPWR VPWR pp_row95_4 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_90_1 pp_row90_14 pp_row90_15 pp_row90_16 VGND VGND VPWR VPWR c$1808 s$1809
+ sky130_fd_sc_hd__fa_1
XFILLER_12_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_83_0 pp_row83_21 pp_row83_22 pp_row83_23 VGND VGND VPWR VPWR c$1722 s$1723
+ sky130_fd_sc_hd__fa_1
XFILLER_141_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1506_ clknet_leaf_164_clk booth_b60_m63 VGND VGND VPWR VPWR pp_row123_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_130_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2486_ clknet_leaf_146_clk booth_b14_m55 VGND VGND VPWR VPWR pp_row69_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_68_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1437_ clknet_leaf_53_clk booth_b2_m33 VGND VGND VPWR VPWR pp_row35_1 sky130_fd_sc_hd__dfxtp_1
X_1368_ clknet_leaf_4_clk booth_b28_m3 VGND VGND VPWR VPWR pp_row31_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_95_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_52_6 pp_row52_20 pp_row52_21 pp_row52_22 VGND VGND VPWR VPWR c$396 s$397
+ sky130_fd_sc_hd__fa_1
XFILLER_83_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0319_ clknet_leaf_200_clk booth_b16_m58 VGND VGND VPWR VPWR pp_row74_4 sky130_fd_sc_hd__dfxtp_1
X_1299_ clknet_leaf_250_clk booth_b4_m24 VGND VGND VPWR VPWR pp_row28_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_83_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_4_0 s$3417 c$3902 s$3905 VGND VGND VPWR VPWR c$4160 s$4161 sky130_fd_sc_hd__fa_1
XFILLER_12_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$1009 final_adder.$signal$1138 final_adder.g_new$947 VGND VGND VPWR
+ VPWR net327 sky130_fd_sc_hd__xor2_2
XFILLER_20_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_82_0 s$3727 c$4058 s$4061 VGND VGND VPWR VPWR c$4316 s$4317 sky130_fd_sc_hd__fa_2
Xdadda_fa_4_98_0 s$1913 c$2614 c$2616 VGND VGND VPWR VPWR c$3278 s$3279 sky130_fd_sc_hd__fa_1
XFILLER_180_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1305 net1308 VGND VGND VPWR VPWR net1305 sky130_fd_sc_hd__buf_4
Xfanout1316 net1317 VGND VGND VPWR VPWR net1316 sky130_fd_sc_hd__buf_4
Xfanout1327 net1328 VGND VGND VPWR VPWR net1327 sky130_fd_sc_hd__buf_8
Xfanout1338 net1347 VGND VGND VPWR VPWR net1338 sky130_fd_sc_hd__buf_6
Xfanout1349 net1352 VGND VGND VPWR VPWR net1349 sky130_fd_sc_hd__clkbuf_8
XFILLER_93_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout395 net400 VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__buf_4
XFILLER_46_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3107 t$5992 net1361 VGND VGND VPWR VPWR booth_b44_m43 sky130_fd_sc_hd__xor2_1
XFILLER_59_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3118 net1693 net515 net1684 net788 VGND VGND VPWR VPWR t$5998 sky130_fd_sc_hd__a22o_1
XFILLER_98_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3129 t$6003 net1364 VGND VGND VPWR VPWR booth_b44_m54 sky130_fd_sc_hd__xor2_1
XU$$2406 t$5634 net1428 VGND VGND VPWR VPWR booth_b34_m35 sky130_fd_sc_hd__xor2_1
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2417 net926 net565 net1747 net838 VGND VGND VPWR VPWR t$5640 sky130_fd_sc_hd__a22o_1
XFILLER_62_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2428 t$5645 net1425 VGND VGND VPWR VPWR booth_b34_m46 sky130_fd_sc_hd__xor2_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2439 net1647 net566 net1639 net839 VGND VGND VPWR VPWR t$5651 sky130_fd_sc_hd__a22o_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1705 t$5276 net1469 VGND VGND VPWR VPWR booth_b24_m27 sky130_fd_sc_hd__xor2_1
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1716 net1000 net605 net992 net878 VGND VGND VPWR VPWR t$5282 sky130_fd_sc_hd__a22o_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1727 t$5287 net1468 VGND VGND VPWR VPWR booth_b24_m38 sky130_fd_sc_hd__xor2_1
XFILLER_43_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1738 net1735 net609 net1727 net882 VGND VGND VPWR VPWR t$5293 sky130_fd_sc_hd__a22o_1
XU$$1749 t$5298 net1473 VGND VGND VPWR VPWR booth_b24_m49 sky130_fd_sc_hd__xor2_1
XFILLER_42_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput15 a[22] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_2
XFILLER_7_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput26 a[32] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_2
Xinput37 a[42] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_2
XFILLER_156_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput48 a[52] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput59 a[62] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dlymetal6s2s_1
X_0670_ clknet_leaf_180_clk booth_b24_m62 VGND VGND VPWR VPWR pp_row86_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_171_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2340_ clknet_leaf_89_clk booth_b12_m53 VGND VGND VPWR VPWR pp_row65_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_69_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2271_ clknet_leaf_129_clk booth_b58_m52 VGND VGND VPWR VPWR pp_row110_7 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_62_5 s$575 s$577 s$579 VGND VGND VPWR VPWR c$1480 s$1481 sky130_fd_sc_hd__fa_2
XFILLER_96_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1222_ clknet_leaf_48_clk booth_b12_m11 VGND VGND VPWR VPWR pp_row23_6 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_55_4 s$443 s$445 s$447 VGND VGND VPWR VPWR c$1394 s$1395 sky130_fd_sc_hd__fa_1
XU$$4320 t$6612 net1262 VGND VGND VPWR VPWR booth_b62_m33 sky130_fd_sc_hd__xor2_1
XU$$4331 net953 net424 net945 net706 VGND VGND VPWR VPWR t$6618 sky130_fd_sc_hd__a22o_1
XFILLER_42_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4342 t$6623 net1255 VGND VGND VPWR VPWR booth_b62_m44 sky130_fd_sc_hd__xor2_1
XFILLER_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4353 net1680 net419 net1655 net701 VGND VGND VPWR VPWR t$6629 sky130_fd_sc_hd__a22o_1
X_1153_ clknet_leaf_15_clk booth_b12_m6 VGND VGND VPWR VPWR pp_row18_6 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_48_3 c$312 c$314 s$317 VGND VGND VPWR VPWR c$1308 s$1309 sky130_fd_sc_hd__fa_1
XU$$4364 t$6634 net1256 VGND VGND VPWR VPWR booth_b62_m55 sky130_fd_sc_hd__xor2_1
XU$$3630 net1028 net477 net1020 net750 VGND VGND VPWR VPWR t$6260 sky130_fd_sc_hd__a22o_1
XU$$4375 net1554 net420 net1545 net702 VGND VGND VPWR VPWR t$6640 sky130_fd_sc_hd__a22o_1
XU$$3641 t$6265 net1321 VGND VGND VPWR VPWR booth_b52_m36 sky130_fd_sc_hd__xor2_1
XU$$4386 net1811 VGND VGND VPWR VPWR notblock$6645\[2\] sky130_fd_sc_hd__inv_1
XU$$4397 t$6652 net1819 VGND VGND VPWR VPWR booth_b64_m3 sky130_fd_sc_hd__xor2_1
XFILLER_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3652 net1751 net481 net1743 net754 VGND VGND VPWR VPWR t$6271 sky130_fd_sc_hd__a22o_1
XU$$3663 t$6276 net1326 VGND VGND VPWR VPWR booth_b52_m47 sky130_fd_sc_hd__xor2_1
X_1084_ clknet_leaf_58_clk booth_b0_m12 VGND VGND VPWR VPWR pp_row12_0 sky130_fd_sc_hd__dfxtp_1
XU$$3674 net1644 net482 net1635 net755 VGND VGND VPWR VPWR t$6282 sky130_fd_sc_hd__a22o_1
XFILLER_65_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2940 t$5907 net1371 VGND VGND VPWR VPWR booth_b42_m28 sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_18_1 s$2799 s$2801 s$2803 VGND VGND VPWR VPWR c$3470 s$3471 sky130_fd_sc_hd__fa_1
XU$$3685 t$6287 net1327 VGND VGND VPWR VPWR booth_b52_m58 sky130_fd_sc_hd__xor2_1
XU$$2951 net994 net521 net984 net794 VGND VGND VPWR VPWR t$5913 sky130_fd_sc_hd__a22o_1
XU$$3696 net1529 net477 net1796 net750 VGND VGND VPWR VPWR t$6293 sky130_fd_sc_hd__a22o_1
XU$$2962 t$5918 net1369 VGND VGND VPWR VPWR booth_b42_m39 sky130_fd_sc_hd__xor2_1
XU$$2973 net1723 net521 net1714 net794 VGND VGND VPWR VPWR t$5924 sky130_fd_sc_hd__a22o_1
XU$$2984 t$5929 net1373 VGND VGND VPWR VPWR booth_b42_m50 sky130_fd_sc_hd__xor2_1
XU$$2995 net1618 net524 net1609 net797 VGND VGND VPWR VPWR t$5935 sky130_fd_sc_hd__a22o_1
XFILLER_34_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1986_ clknet_leaf_81_clk booth_b10_m45 VGND VGND VPWR VPWR pp_row55_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_193_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0937_ clknet_leaf_104_clk booth_b60_m37 VGND VGND VPWR VPWR pp_row97_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_107_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_9_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_174_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0868_ clknet_leaf_111_clk booth_b44_m50 VGND VGND VPWR VPWR pp_row94_8 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_5_15__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_5_15__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_161_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0799_ clknet_leaf_132_clk booth_b56_m63 VGND VGND VPWR VPWR pp_row119_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_115_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2469_ clknet_leaf_124_clk booth_b52_m60 VGND VGND VPWR VPWR pp_row112_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_87_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$902 final_adder.$signal$1208 final_adder.g_new$973 final_adder.$signal$238
+ VGND VGND VPWR VPWR final_adder.g_new$1030 sky130_fd_sc_hd__a21o_1
XFILLER_180_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$913 final_adder.$signal$1186 final_adder.g_new$995 final_adder.$signal$194
+ VGND VGND VPWR VPWR final_adder.g_new$1041 sky130_fd_sc_hd__a21o_1
XFILLER_68_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$924 final_adder.$signal$1164 final_adder.g_new$1017 final_adder.$signal$150
+ VGND VGND VPWR VPWR final_adder.g_new$1052 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$935 final_adder.$signal$107 final_adder.g_new$943 final_adder.$signal$106
+ VGND VGND VPWR VPWR final_adder.g_new$1063 sky130_fd_sc_hd__a21o_1
Xdadda_fa_1_50_3 pp_row50_9 pp_row50_10 pp_row50_11 VGND VGND VPWR VPWR c$354 s$355
+ sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$946 final_adder.$signal$1120 final_adder.g_new$853 final_adder.$signal$62
+ VGND VGND VPWR VPWR final_adder.g_new$1074 sky130_fd_sc_hd__a21o_1
XFILLER_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$957 final_adder.$signal$1098 final_adder.g_new$631 final_adder.$signal$18
+ VGND VGND VPWR VPWR final_adder.g_new$1085 sky130_fd_sc_hd__a21o_1
XFILLER_110_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$968 final_adder.$signal$1097 final_adder.g_new$1086 VGND VGND VPWR
+ VPWR net362 sky130_fd_sc_hd__xor2_2
XU$$807 net1599 net407 net1590 net673 VGND VGND VPWR VPWR t$4817 sky130_fd_sc_hd__a22o_1
XU$$818 t$4822 net1417 VGND VGND VPWR VPWR booth_b10_m63 sky130_fd_sc_hd__xor2_1
XFILLER_113_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$979 final_adder.$signal$1108 final_adder.g_new$865 VGND VGND VPWR
+ VPWR net294 sky130_fd_sc_hd__xor2_2
Xdadda_fa_1_43_2 pp_row43_6 pp_row43_7 pp_row43_8 VGND VGND VPWR VPWR c$258 s$259
+ sky130_fd_sc_hd__fa_1
XFILLER_3_1050 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$829 t$4829 net1312 VGND VGND VPWR VPWR booth_b12_m0 sky130_fd_sc_hd__xor2_1
XFILLER_43_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_20_1 c$1994 c$1996 s$1999 VGND VGND VPWR VPWR c$2812 s$2813 sky130_fd_sc_hd__fa_1
XFILLER_3_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_13_0 pp_row13_0 pp_row13_1 pp_row13_2 VGND VGND VPWR VPWR c$2768 s$2769
+ sky130_fd_sc_hd__fa_1
XFILLER_169_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3833_1798 VGND VGND VPWR VPWR U$$3833_1798/HI net1798 sky130_fd_sc_hd__conb_1
XFILLER_184_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1102 net1104 VGND VGND VPWR VPWR net1102 sky130_fd_sc_hd__clkbuf_8
Xfanout1113 net78 VGND VGND VPWR VPWR net1113 sky130_fd_sc_hd__buf_4
Xdadda_fa_3_65_3 s$1511 s$1513 s$1515 VGND VGND VPWR VPWR c$2364 s$2365 sky130_fd_sc_hd__fa_1
Xfanout1124 net1125 VGND VGND VPWR VPWR net1124 sky130_fd_sc_hd__buf_2
Xfanout1135 net1136 VGND VGND VPWR VPWR net1135 sky130_fd_sc_hd__buf_6
Xfanout1146 net1147 VGND VGND VPWR VPWR net1146 sky130_fd_sc_hd__buf_4
Xfanout1157 net1158 VGND VGND VPWR VPWR net1157 sky130_fd_sc_hd__buf_4
Xdadda_fa_3_58_2 c$1420 s$1423 s$1425 VGND VGND VPWR VPWR c$2306 s$2307 sky130_fd_sc_hd__fa_1
Xfanout1168 net71 VGND VGND VPWR VPWR net1168 sky130_fd_sc_hd__clkbuf_8
Xfanout1179 net1181 VGND VGND VPWR VPWR net1179 sky130_fd_sc_hd__buf_6
XFILLER_59_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_28_0 c$3504 c$3506 s$3509 VGND VGND VPWR VPWR c$3952 s$3953 sky130_fd_sc_hd__fa_1
XU$$2203 t$5531 net1432 VGND VGND VPWR VPWR booth_b32_m2 sky130_fd_sc_hd__xor2_1
XU$$2214 net1511 net569 net1503 net842 VGND VGND VPWR VPWR t$5537 sky130_fd_sc_hd__a22o_1
XU$$2225 t$5542 net1431 VGND VGND VPWR VPWR booth_b32_m13 sky130_fd_sc_hd__xor2_1
XU$$2236 net1144 net571 net1134 net844 VGND VGND VPWR VPWR t$5548 sky130_fd_sc_hd__a22o_1
XU$$2247 t$5553 net1433 VGND VGND VPWR VPWR booth_b32_m24 sky130_fd_sc_hd__xor2_1
XU$$1502 net1536 net633 net1528 net906 VGND VGND VPWR VPWR t$5172 sky130_fd_sc_hd__a22o_1
XU$$2258 net1040 net570 net1024 net843 VGND VGND VPWR VPWR t$5559 sky130_fd_sc_hd__a22o_1
XU$$1513 net1763 net613 net1230 net886 VGND VGND VPWR VPWR t$5179 sky130_fd_sc_hd__a22o_1
XU$$2269 t$5564 net1438 VGND VGND VPWR VPWR booth_b32_m35 sky130_fd_sc_hd__xor2_1
XU$$1524 t$5184 net1475 VGND VGND VPWR VPWR booth_b22_m5 sky130_fd_sc_hd__xor2_1
XFILLER_37_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1535 net1224 net614 net1216 net887 VGND VGND VPWR VPWR t$5190 sky130_fd_sc_hd__a22o_1
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1546 t$5195 net1478 VGND VGND VPWR VPWR booth_b22_m16 sky130_fd_sc_hd__xor2_1
XU$$1557 net1107 net612 net1098 net885 VGND VGND VPWR VPWR t$5201 sky130_fd_sc_hd__a22o_1
XFILLER_188_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1568 t$5206 net1477 VGND VGND VPWR VPWR booth_b22_m27 sky130_fd_sc_hd__xor2_1
XU$$1579 net1001 net614 net993 net887 VGND VGND VPWR VPWR t$5212 sky130_fd_sc_hd__a22o_1
XFILLER_15_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1840_ clknet_leaf_62_clk booth_b30_m20 VGND VGND VPWR VPWR pp_row50_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1771_ clknet_leaf_238_clk booth_b14_m34 VGND VGND VPWR VPWR pp_row48_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0722_ clknet_leaf_181_clk net158 VGND VGND VPWR VPWR pp_row126_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_128_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0653_ clknet_leaf_169_clk booth_b40_m45 VGND VGND VPWR VPWR pp_row85_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_171_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0584_ clknet_leaf_174_clk booth_b62_m20 VGND VGND VPWR VPWR pp_row82_23 sky130_fd_sc_hd__dfxtp_1
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2323_ clknet_leaf_74_clk booth_b48_m16 VGND VGND VPWR VPWR pp_row64_24 sky130_fd_sc_hd__dfxtp_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_2_60_2 c$520 c$522 c$524 VGND VGND VPWR VPWR c$1450 s$1451 sky130_fd_sc_hd__fa_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$209 final_adder.$signal$1137 final_adder.$signal$94 final_adder.$signal$96
+ VGND VGND VPWR VPWR final_adder.g_new$337 sky130_fd_sc_hd__a21o_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2254_ clknet_leaf_148_clk booth_b58_m4 VGND VGND VPWR VPWR pp_row62_29 sky130_fd_sc_hd__dfxtp_1
XFILLER_111_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_53_1 c$388 c$390 c$392 VGND VGND VPWR VPWR c$1364 s$1365 sky130_fd_sc_hd__fa_1
XFILLER_38_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1680 net1681 VGND VGND VPWR VPWR net1680 sky130_fd_sc_hd__buf_6
X_1205_ clknet_leaf_143_clk booth_b44_m59 VGND VGND VPWR VPWR pp_row103_3 sky130_fd_sc_hd__dfxtp_1
Xfanout1691 net107 VGND VGND VPWR VPWR net1691 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_5_30_0 c$2864 c$2866 c$2868 VGND VGND VPWR VPWR c$3516 s$3517 sky130_fd_sc_hd__fa_1
X_2185_ clknet_leaf_216_clk net1263 VGND VGND VPWR VPWR pp_row60_31 sky130_fd_sc_hd__dfxtp_1
XU$$4150 net1160 net436 net1152 net718 VGND VGND VPWR VPWR t$6526 sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_46_0 pp_row46_20 pp_row46_21 pp_row46_22 VGND VGND VPWR VPWR c$1278 s$1279
+ sky130_fd_sc_hd__fa_1
XU$$4161 t$6531 net1268 VGND VGND VPWR VPWR booth_b60_m22 sky130_fd_sc_hd__xor2_1
XFILLER_81_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4172 net1062 net435 net1053 net717 VGND VGND VPWR VPWR t$6537 sky130_fd_sc_hd__a22o_1
XU$$4183 t$6542 net1272 VGND VGND VPWR VPWR booth_b60_m33 sky130_fd_sc_hd__xor2_1
XFILLER_26_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1136_ clknet_leaf_16_clk booth_b2_m15 VGND VGND VPWR VPWR pp_row17_1 sky130_fd_sc_hd__dfxtp_1
XU$$4194 net953 net440 net945 net722 VGND VGND VPWR VPWR t$6548 sky130_fd_sc_hd__a22o_1
XU$$3460 t$6173 net1333 VGND VGND VPWR VPWR booth_b50_m14 sky130_fd_sc_hd__xor2_1
XU$$3471 net1135 net486 net1119 net759 VGND VGND VPWR VPWR t$6179 sky130_fd_sc_hd__a22o_1
XU$$3482 t$6184 net1331 VGND VGND VPWR VPWR booth_b50_m25 sky130_fd_sc_hd__xor2_1
XU$$3493 net1027 net485 net1019 net758 VGND VGND VPWR VPWR t$6190 sky130_fd_sc_hd__a22o_1
X_1067_ clknet_leaf_51_clk booth_b0_m10 VGND VGND VPWR VPWR pp_row10_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_53_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_901 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2770 net1218 net539 net1207 net812 VGND VGND VPWR VPWR t$5821 sky130_fd_sc_hd__a22o_1
XU$$2781 t$5826 net1384 VGND VGND VPWR VPWR booth_b40_m17 sky130_fd_sc_hd__xor2_1
XFILLER_178_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2792 net1102 net538 net1094 net811 VGND VGND VPWR VPWR t$5832 sky130_fd_sc_hd__a22o_1
XFILLER_178_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1969_ clknet_leaf_72_clk booth_b40_m14 VGND VGND VPWR VPWR pp_row54_20 sky130_fd_sc_hd__dfxtp_1
XFILLER_147_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_814 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_75_2 s$2441 s$2443 s$2445 VGND VGND VPWR VPWR c$3144 s$3145 sky130_fd_sc_hd__fa_1
XFILLER_122_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_68_1 c$2378 c$2380 s$2383 VGND VGND VPWR VPWR c$3100 s$3101 sky130_fd_sc_hd__fa_1
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_755 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput205 c[53] VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__clkbuf_1
Xinput216 c[63] VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_7_45_0 s$3579 c$3984 s$3987 VGND VGND VPWR VPWR c$4242 s$4243 sky130_fd_sc_hd__fa_2
XFILLER_89_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_251_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_251_clk
+ sky130_fd_sc_hd__clkbuf_16
Xinput227 c[73] VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput238 c[83] VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__clkbuf_1
Xdadda_ha_1_35_0 pp_row35_0 pp_row35_1 VGND VGND VPWR VPWR c$206 s$207 sky130_fd_sc_hd__ha_1
Xinput249 c[93] VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__clkbuf_1
Xfinal_adder.U$$710 final_adder.p_new$734 final_adder.p_new$718 VGND VGND VPWR VPWR
+ final_adder.p_new$838 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$721 final_adder.p_new$728 final_adder.g_new$745 final_adder.g_new$729
+ VGND VGND VPWR VPWR final_adder.g_new$849 sky130_fd_sc_hd__a21o_1
XFILLER_5_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$743 final_adder.p_new$758 final_adder.g_new$791 final_adder.g_new$759
+ VGND VGND VPWR VPWR final_adder.g_new$871 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$754 final_adder.p_new$802 final_adder.p_new$770 VGND VGND VPWR VPWR
+ final_adder.p_new$882 sky130_fd_sc_hd__and2_1
XU$$604 net1083 net413 net1074 net679 VGND VGND VPWR VPWR t$4714 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$765 final_adder.p_new$780 final_adder.g_new$813 final_adder.g_new$781
+ VGND VGND VPWR VPWR final_adder.g_new$893 sky130_fd_sc_hd__a21o_1
XFILLER_1_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$776 final_adder.p_new$824 final_adder.p_new$792 VGND VGND VPWR VPWR
+ final_adder.p_new$904 sky130_fd_sc_hd__and2_1
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$615 t$4719 net1236 VGND VGND VPWR VPWR booth_b8_m30 sky130_fd_sc_hd__xor2_1
XU$$626 net973 net410 net964 net676 VGND VGND VPWR VPWR t$4725 sky130_fd_sc_hd__a22o_1
XFILLER_57_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1016 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$787 final_adder.p_new$802 final_adder.g_new$835 final_adder.g_new$803
+ VGND VGND VPWR VPWR final_adder.g_new$915 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$798 final_adder.p_new$846 final_adder.p_new$814 VGND VGND VPWR VPWR
+ final_adder.p_new$926 sky130_fd_sc_hd__and2_1
XU$$637 t$4730 net1238 VGND VGND VPWR VPWR booth_b8_m41 sky130_fd_sc_hd__xor2_1
XFILLER_112_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$648 net1707 net416 net1699 net682 VGND VGND VPWR VPWR t$4736 sky130_fd_sc_hd__a22o_1
XU$$659 t$4741 net1238 VGND VGND VPWR VPWR booth_b8_m52 sky130_fd_sc_hd__xor2_1
XFILLER_31_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_978 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_70_1 c$1558 c$1560 c$1562 VGND VGND VPWR VPWR c$2400 s$2401 sky130_fd_sc_hd__fa_1
XFILLER_79_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_63_0 s$599 c$1470 c$1472 VGND VGND VPWR VPWR c$2342 s$2343 sky130_fd_sc_hd__fa_1
Xclkbuf_leaf_242_clk clknet_5_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_242_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2000 net961 net588 net955 net861 VGND VGND VPWR VPWR t$5427 sky130_fd_sc_hd__a22o_1
XU$$2011 t$5432 net1454 VGND VGND VPWR VPWR booth_b28_m43 sky130_fd_sc_hd__xor2_1
XFILLER_63_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2022 net1692 net591 net1685 net864 VGND VGND VPWR VPWR t$5438 sky130_fd_sc_hd__a22o_1
XU$$2033 t$5443 net1454 VGND VGND VPWR VPWR booth_b28_m54 sky130_fd_sc_hd__xor2_1
XFILLER_74_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2044 net1580 net591 net1553 net864 VGND VGND VPWR VPWR t$5449 sky130_fd_sc_hd__a22o_1
XU$$1310 t$5074 net1666 VGND VGND VPWR VPWR booth_b18_m35 sky130_fd_sc_hd__xor2_1
XU$$2055 net1454 VGND VGND VPWR VPWR notblock$5455\[0\] sky130_fd_sc_hd__inv_1
XU$$1321 net925 net640 net1746 net913 VGND VGND VPWR VPWR t$5080 sky130_fd_sc_hd__a22o_1
XU$$2066 t$5461 net1441 VGND VGND VPWR VPWR booth_b30_m2 sky130_fd_sc_hd__xor2_1
XU$$2077 net1511 net576 net1503 net849 VGND VGND VPWR VPWR t$5467 sky130_fd_sc_hd__a22o_1
XU$$1332 t$5085 net1670 VGND VGND VPWR VPWR booth_b18_m46 sky130_fd_sc_hd__xor2_1
XU$$2088 t$5472 net1439 VGND VGND VPWR VPWR booth_b30_m13 sky130_fd_sc_hd__xor2_1
XU$$4244_1807 VGND VGND VPWR VPWR U$$4244_1807/HI net1807 sky130_fd_sc_hd__conb_1
XU$$1343 net1646 net642 net1640 net915 VGND VGND VPWR VPWR t$5091 sky130_fd_sc_hd__a22o_1
XU$$1354 t$5096 net1669 VGND VGND VPWR VPWR booth_b18_m57 sky130_fd_sc_hd__xor2_1
XU$$2099 net1139 net577 net1132 net850 VGND VGND VPWR VPWR t$5478 sky130_fd_sc_hd__a22o_1
XU$$1365 net1537 net641 net1528 net914 VGND VGND VPWR VPWR t$5102 sky130_fd_sc_hd__a22o_1
XU$$1376 net1760 net630 net1230 net903 VGND VGND VPWR VPWR t$5109 sky130_fd_sc_hd__a22o_1
XU$$1387 t$5114 net1485 VGND VGND VPWR VPWR booth_b20_m5 sky130_fd_sc_hd__xor2_1
XU$$1398 net1219 net627 net1210 net900 VGND VGND VPWR VPWR t$5120 sky130_fd_sc_hd__a22o_1
Xdadda_fa_7_120_0 s$3879 c$4134 s$4137 VGND VGND VPWR VPWR c$4392 s$4393 sky130_fd_sc_hd__fa_1
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1823_ clknet_leaf_234_clk booth_b2_m48 VGND VGND VPWR VPWR pp_row50_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_157_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1754_ clknet_leaf_238_clk booth_b32_m15 VGND VGND VPWR VPWR pp_row47_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_8_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_85_1 s$3201 s$3203 s$3205 VGND VGND VPWR VPWR c$3738 s$3739 sky130_fd_sc_hd__fa_1
XFILLER_156_493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0705_ clknet_leaf_172_clk booth_b42_m45 VGND VGND VPWR VPWR pp_row87_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_128_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1685_ clknet_leaf_19_clk booth_b8_m37 VGND VGND VPWR VPWR pp_row45_4 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_78_0 c$3152 c$3154 c$3156 VGND VGND VPWR VPWR c$3708 s$3709 sky130_fd_sc_hd__fa_1
X_0636_ clknet_leaf_174_clk booth_b56_m28 VGND VGND VPWR VPWR pp_row84_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_131_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout906 net907 VGND VGND VPWR VPWR net906 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout917 net920 VGND VGND VPWR VPWR net917 sky130_fd_sc_hd__buf_6
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout928 net931 VGND VGND VPWR VPWR net928 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_77_8 pp_row77_27 c$196 c$198 VGND VGND VPWR VPWR c$850 s$851 sky130_fd_sc_hd__fa_2
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0567_ clknet_leaf_188_clk booth_b30_m52 VGND VGND VPWR VPWR pp_row82_7 sky130_fd_sc_hd__dfxtp_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout939 net98 VGND VGND VPWR VPWR net939 sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_233_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_233_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2306_ clknet_leaf_84_clk booth_b16_m48 VGND VGND VPWR VPWR pp_row64_8 sky130_fd_sc_hd__dfxtp_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0498_ clknet_leaf_208_clk booth_b62_m17 VGND VGND VPWR VPWR pp_row79_24 sky130_fd_sc_hd__dfxtp_1
XFILLER_100_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2237_ clknet_leaf_228_clk booth_b28_m34 VGND VGND VPWR VPWR pp_row62_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_39_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2168_ clknet_leaf_28_clk booth_b34_m26 VGND VGND VPWR VPWR pp_row60_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_65_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1119_ clknet_leaf_48_clk booth_b10_m5 VGND VGND VPWR VPWR pp_row15_5 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$50 c$4250 s$4253 VGND VGND VPWR VPWR final_adder.$signal$102 final_adder.$signal$103
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$61 c$4272 s$4275 VGND VGND VPWR VPWR final_adder.$signal$124 final_adder.$signal$1151
+ sky130_fd_sc_hd__ha_1
XFILLER_0_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3290 net1340 VGND VGND VPWR VPWR notblock$6085\[2\] sky130_fd_sc_hd__inv_1
X_2099_ clknet_leaf_32_clk booth_b34_m24 VGND VGND VPWR VPWR pp_row58_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_81_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$72 c$4294 s$4297 VGND VGND VPWR VPWR final_adder.$signal$146 final_adder.$signal$1162
+ sky130_fd_sc_hd__ha_1
XFILLER_13_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$83 c$4316 s$4319 VGND VGND VPWR VPWR final_adder.$signal$168 final_adder.$signal$1173
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$94 c$4338 s$4341 VGND VGND VPWR VPWR final_adder.$signal$190 final_adder.$signal$1184
+ sky130_fd_sc_hd__ha_1
XFILLER_94_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1650_1765 VGND VGND VPWR VPWR U$$1650_1765/HI net1765 sky130_fd_sc_hd__conb_1
XFILLER_108_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_80_0 s$1697 c$2470 c$2472 VGND VGND VPWR VPWR c$3170 s$3171 sky130_fd_sc_hd__fa_1
Xdadda_fa_3_101_3 s$1935 s$1937 s$1939 VGND VGND VPWR VPWR c$2652 s$2653 sky130_fd_sc_hd__fa_1
XFILLER_123_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_224_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_224_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_49_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$540 final_adder.p_new$552 final_adder.p_new$544 VGND VGND VPWR VPWR
+ final_adder.p_new$668 sky130_fd_sc_hd__and2_1
XTAP_3822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$551 final_adder.p_new$554 final_adder.g_new$563 final_adder.g_new$555
+ VGND VGND VPWR VPWR final_adder.g_new$679 sky130_fd_sc_hd__a21o_1
XTAP_3833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$401 t$4609 net1275 VGND VGND VPWR VPWR booth_b4_m60 sky130_fd_sc_hd__xor2_1
Xdadda_fa_6_108_0 c$3824 c$3826 s$3829 VGND VGND VPWR VPWR c$4112 s$4113 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$562 final_adder.p_new$574 final_adder.p_new$566 VGND VGND VPWR VPWR
+ final_adder.p_new$690 sky130_fd_sc_hd__and2_1
XTAP_3844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$412 net61 VGND VGND VPWR VPWR notblock$4615\[1\] sky130_fd_sc_hd__inv_1
Xfinal_adder.U$$573 final_adder.p_new$576 final_adder.g_new$585 final_adder.g_new$577
+ VGND VGND VPWR VPWR final_adder.g_new$701 sky130_fd_sc_hd__a21o_1
XTAP_3855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$584 final_adder.p_new$596 final_adder.p_new$588 VGND VGND VPWR VPWR
+ final_adder.p_new$712 sky130_fd_sc_hd__and2_1
XU$$423 net1035 net430 net937 net712 VGND VGND VPWR VPWR t$4622 sky130_fd_sc_hd__a22o_1
XTAP_3866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$434 t$4627 net1250 VGND VGND VPWR VPWR booth_b6_m8 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$595 final_adder.p_new$598 final_adder.g_new$607 final_adder.g_new$599
+ VGND VGND VPWR VPWR final_adder.g_new$723 sky130_fd_sc_hd__a21o_1
XTAP_3877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$445 net1198 net429 net1179 net711 VGND VGND VPWR VPWR t$4633 sky130_fd_sc_hd__a22o_1
XFILLER_189_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$456 t$4638 net1245 VGND VGND VPWR VPWR booth_b6_m19 sky130_fd_sc_hd__xor2_1
XTAP_3899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_28_3 s$1075 s$1077 s$1079 VGND VGND VPWR VPWR c$2068 s$2069 sky130_fd_sc_hd__fa_1
XU$$467 net1080 net428 net1071 net710 VGND VGND VPWR VPWR t$4644 sky130_fd_sc_hd__a22o_1
XU$$478 t$4649 net1250 VGND VGND VPWR VPWR booth_b6_m30 sky130_fd_sc_hd__xor2_1
XU$$489 net973 net426 net964 net708 VGND VGND VPWR VPWR t$4655 sky130_fd_sc_hd__a22o_1
XFILLER_189_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_95_0 c$3772 c$3774 s$3777 VGND VGND VPWR VPWR c$4086 s$4087 sky130_fd_sc_hd__fa_1
XFILLER_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1470_ clknet_leaf_39_clk booth_b24_m12 VGND VGND VPWR VPWR pp_row36_12 sky130_fd_sc_hd__dfxtp_1
X_0421_ clknet_leaf_207_clk booth_b30_m47 VGND VGND VPWR VPWR pp_row77_9 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_215_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_215_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_122_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0352_ clknet_leaf_200_clk booth_b18_m57 VGND VGND VPWR VPWR pp_row75_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_95_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0283_ clknet_leaf_202_clk notsign$4754 VGND VGND VPWR VPWR pp_row73_0 sky130_fd_sc_hd__dfxtp_1
X_2022_ clknet_leaf_34_clk booth_b18_m38 VGND VGND VPWR VPWR pp_row56_9 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_30_3 pp_row30_9 pp_row30_10 pp_row30_11 VGND VGND VPWR VPWR c$1096 s$1097
+ sky130_fd_sc_hd__fa_1
XFILLER_39_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$990 t$4911 net1183 VGND VGND VPWR VPWR booth_b14_m12 sky130_fd_sc_hd__xor2_1
XU$$1140 net1144 net647 net1133 net920 VGND VGND VPWR VPWR t$4988 sky130_fd_sc_hd__a22o_1
XU$$1151 t$4993 net1006 VGND VGND VPWR VPWR booth_b16_m24 sky130_fd_sc_hd__xor2_1
XU$$1162 net1039 net644 net1023 net917 VGND VGND VPWR VPWR t$4999 sky130_fd_sc_hd__a22o_1
XU$$1173 t$5004 net1010 VGND VGND VPWR VPWR booth_b16_m35 sky130_fd_sc_hd__xor2_1
XU$$4441_1841 VGND VGND VPWR VPWR U$$4441_1841/HI net1841 sky130_fd_sc_hd__conb_1
XU$$1184 net928 net645 net1749 net918 VGND VGND VPWR VPWR t$5010 sky130_fd_sc_hd__a22o_1
XU$$1195 t$5015 net1007 VGND VGND VPWR VPWR booth_b16_m46 sky130_fd_sc_hd__xor2_1
XFILLER_176_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1806_ clknet_leaf_220_clk booth_b22_m27 VGND VGND VPWR VPWR pp_row49_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_145_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1737_ clknet_leaf_236_clk booth_b2_m45 VGND VGND VPWR VPWR pp_row47_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_105_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1668_ clknet_leaf_20_clk booth_b28_m16 VGND VGND VPWR VPWR pp_row44_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_131_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_82_6 pp_row82_18 pp_row82_19 pp_row82_20 VGND VGND VPWR VPWR c$934 s$935
+ sky130_fd_sc_hd__fa_1
XFILLER_104_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout703 sel_1$6578 VGND VGND VPWR VPWR net703 sky130_fd_sc_hd__buf_6
XFILLER_160_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0619_ clknet_leaf_187_clk booth_b26_m58 VGND VGND VPWR VPWR pp_row84_4 sky130_fd_sc_hd__dfxtp_1
Xfanout714 net715 VGND VGND VPWR VPWR net714 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_75_5 pp_row75_21 pp_row75_22 pp_row75_23 VGND VGND VPWR VPWR c$808 s$809
+ sky130_fd_sc_hd__fa_1
X_1599_ clknet_leaf_244_clk net192 VGND VGND VPWR VPWR pp_row41_21 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_206_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_206_clk
+ sky130_fd_sc_hd__clkbuf_16
Xfanout725 net732 VGND VGND VPWR VPWR net725 sky130_fd_sc_hd__buf_2
XFILLER_86_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout736 sel_1$6368 VGND VGND VPWR VPWR net736 sky130_fd_sc_hd__clkbuf_8
Xfanout747 net748 VGND VGND VPWR VPWR net747 sky130_fd_sc_hd__buf_4
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout758 net760 VGND VGND VPWR VPWR net758 sky130_fd_sc_hd__buf_4
XFILLER_140_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout769 sel_1$6088 VGND VGND VPWR VPWR net769 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_68_4 pp_row68_29 pp_row68_30 pp_row68_31 VGND VGND VPWR VPWR c$680 s$681
+ sky130_fd_sc_hd__fa_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_38_2 s$2145 s$2147 s$2149 VGND VGND VPWR VPWR c$2922 s$2923 sky130_fd_sc_hd__fa_1
XFILLER_96_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 net583 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 net644 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_129 net703 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_63_3 pp_row63_9 pp_row63_10 pp_row63_11 VGND VGND VPWR VPWR c$78 s$79
+ sky130_fd_sc_hd__fa_1
XTAP_4331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_40_2 c$1204 s$1207 s$1209 VGND VGND VPWR VPWR c$2162 s$2163 sky130_fd_sc_hd__fa_1
XTAP_4364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$370 final_adder.p_new$372 final_adder.p_new$370 VGND VGND VPWR VPWR
+ final_adder.p_new$498 sky130_fd_sc_hd__and2_1
XTAP_4397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$381 final_adder.p_new$380 final_adder.g_new$383 final_adder.g_new$381
+ VGND VGND VPWR VPWR final_adder.g_new$509 sky130_fd_sc_hd__a21o_4
XU$$220 t$4517 net1385 VGND VGND VPWR VPWR booth_b2_m38 sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_33_1 c$1114 c$1116 c$1118 VGND VGND VPWR VPWR c$2104 s$2105 sky130_fd_sc_hd__fa_1
XTAP_3663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$392 final_adder.p_new$398 final_adder.p_new$394 VGND VGND VPWR VPWR
+ final_adder.p_new$520 sky130_fd_sc_hd__and2_1
XFILLER_17_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$231 net1729 net621 net1720 net894 VGND VGND VPWR VPWR t$4523 sky130_fd_sc_hd__a22o_1
XFILLER_73_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$242 t$4528 net1392 VGND VGND VPWR VPWR booth_b2_m49 sky130_fd_sc_hd__xor2_1
XTAP_3674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_10_0 c$3432 c$3434 s$3437 VGND VGND VPWR VPWR c$3916 s$3917 sky130_fd_sc_hd__fa_1
XFILLER_189_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_26_0 pp_row26_8 pp_row26_9 pp_row26_10 VGND VGND VPWR VPWR c$2046 s$2047
+ sky130_fd_sc_hd__fa_1
XU$$253 net1623 net626 net1615 net899 VGND VGND VPWR VPWR t$4534 sky130_fd_sc_hd__a22o_1
XTAP_3696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$264 t$4539 net1387 VGND VGND VPWR VPWR booth_b2_m60 sky130_fd_sc_hd__xor2_1
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$275 net45 VGND VGND VPWR VPWR notblock$4545\[1\] sky130_fd_sc_hd__inv_1
XTAP_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$286 net1035 net531 net937 net804 VGND VGND VPWR VPWR t$4552 sky130_fd_sc_hd__a22o_1
XFILLER_33_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$297 t$4557 net1277 VGND VGND VPWR VPWR booth_b4_m8 sky130_fd_sc_hd__xor2_1
XTAP_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0970_ clknet_leaf_116_clk booth_b50_m49 VGND VGND VPWR VPWR pp_row99_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_41_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3 net1571 notblock\[1\] VGND VGND VPWR VPWR t sky130_fd_sc_hd__and2_1
Xoutput306 net306 VGND VGND VPWR VPWR o[29] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_92_5 c$1030 s$1033 s$1035 VGND VGND VPWR VPWR c$1840 s$1841 sky130_fd_sc_hd__fa_1
Xoutput317 net317 VGND VGND VPWR VPWR o[39] sky130_fd_sc_hd__buf_2
Xoutput328 net328 VGND VGND VPWR VPWR o[49] sky130_fd_sc_hd__buf_2
XFILLER_160_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1522_ clknet_leaf_242_clk booth_b34_m4 VGND VGND VPWR VPWR pp_row38_17 sky130_fd_sc_hd__dfxtp_1
Xoutput339 net339 VGND VGND VPWR VPWR o[59] sky130_fd_sc_hd__buf_2
XFILLER_181_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_85_4 c$964 s$967 s$969 VGND VGND VPWR VPWR c$1754 s$1755 sky130_fd_sc_hd__fa_1
XU$$4471_1856 VGND VGND VPWR VPWR U$$4471_1856/HI net1856 sky130_fd_sc_hd__conb_1
X_1453_ clknet_leaf_64_clk booth_b30_m5 VGND VGND VPWR VPWR pp_row35_15 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_78_3 c$850 s$853 s$855 VGND VGND VPWR VPWR c$1668 s$1669 sky130_fd_sc_hd__fa_1
XFILLER_68_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0404_ clknet_leaf_208_clk booth_b54_m22 VGND VGND VPWR VPWR pp_row76_22 sky130_fd_sc_hd__dfxtp_1
XFILLER_67_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1384_ clknet_leaf_44_clk booth_b22_m10 VGND VGND VPWR VPWR pp_row32_11 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_48_1 s$2979 s$2981 s$2983 VGND VGND VPWR VPWR c$3590 s$3591 sky130_fd_sc_hd__fa_1
XFILLER_132_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0335_ clknet_leaf_225_clk booth_b44_m30 VGND VGND VPWR VPWR pp_row74_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_110_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0266_ clknet_leaf_124_clk booth_b56_m57 VGND VGND VPWR VPWR pp_row113_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_36_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2005_ clknet_leaf_142_clk booth_b56_m52 VGND VGND VPWR VPWR pp_row108_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_64_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0197_ clknet_leaf_155_clk booth_b36_m34 VGND VGND VPWR VPWR pp_row70_16 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_101_2 pp_row101_6 pp_row101_7 pp_row101_8 VGND VGND VPWR VPWR c$1938 s$1939
+ sky130_fd_sc_hd__fa_1
XFILLER_63_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_122_1 pp_row122_5 c$3412 s$3415 VGND VGND VPWR VPWR c$3886 s$3887 sky130_fd_sc_hd__fa_1
XFILLER_13_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_115_0 c$3374 c$3376 c$3378 VGND VGND VPWR VPWR c$3856 s$3857 sky130_fd_sc_hd__fa_1
XFILLER_192_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_934 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_80_3 pp_row80_9 pp_row80_10 pp_row80_11 VGND VGND VPWR VPWR c$894 s$895
+ sky130_fd_sc_hd__fa_2
Xfanout500 sel_0$6087 VGND VGND VPWR VPWR net500 sky130_fd_sc_hd__buf_6
Xfanout1509 net1510 VGND VGND VPWR VPWR net1509 sky130_fd_sc_hd__buf_4
Xfanout511 net518 VGND VGND VPWR VPWR net511 sky130_fd_sc_hd__buf_4
XFILLER_132_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout522 sel_0$5877 VGND VGND VPWR VPWR net522 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_73_2 pp_row73_15 pp_row73_16 pp_row73_17 VGND VGND VPWR VPWR c$766 s$767
+ sky130_fd_sc_hd__fa_1
Xfanout533 net534 VGND VGND VPWR VPWR net533 sky130_fd_sc_hd__buf_4
Xfanout544 net550 VGND VGND VPWR VPWR net544 sky130_fd_sc_hd__buf_6
XFILLER_116_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout555 net556 VGND VGND VPWR VPWR net555 sky130_fd_sc_hd__buf_4
Xdadda_fa_4_50_1 c$2234 c$2236 s$2239 VGND VGND VPWR VPWR c$2992 s$2993 sky130_fd_sc_hd__fa_1
XFILLER_116_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_66_1 pp_row66_21 pp_row66_22 pp_row66_23 VGND VGND VPWR VPWR c$638 s$639
+ sky130_fd_sc_hd__fa_1
Xfanout566 net568 VGND VGND VPWR VPWR net566 sky130_fd_sc_hd__buf_4
Xdadda_ha_2_100_4 pp_row100_12 pp_row100_13 VGND VGND VPWR VPWR c$1932 s$1933 sky130_fd_sc_hd__ha_1
Xfanout577 net583 VGND VGND VPWR VPWR net577 sky130_fd_sc_hd__clkbuf_4
XFILLER_24_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_864 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout588 net592 VGND VGND VPWR VPWR net588 sky130_fd_sc_hd__buf_6
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_43_0 s$1253 c$2174 c$2176 VGND VGND VPWR VPWR c$2948 s$2949 sky130_fd_sc_hd__fa_1
XFILLER_86_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout599 net600 VGND VGND VPWR VPWR net599 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_1_59_0 pp_row59_11 pp_row59_12 pp_row59_13 VGND VGND VPWR VPWR c$510 s$511
+ sky130_fd_sc_hd__fa_1
XFILLER_111_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1909 net1553 net599 net1544 net872 VGND VGND VPWR VPWR t$5380 sky130_fd_sc_hd__a22o_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_95_3 s$1871 s$1873 s$1875 VGND VGND VPWR VPWR c$2604 s$2605 sky130_fd_sc_hd__fa_1
XFILLER_68_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_912 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_88_2 c$1780 s$1783 s$1785 VGND VGND VPWR VPWR c$2546 s$2547 sky130_fd_sc_hd__fa_1
XFILLER_151_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_0_55_1 pp_row55_3 pp_row55_4 VGND VGND VPWR VPWR c$10 s$11 sky130_fd_sc_hd__ha_1
XFILLER_111_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_58_0 c$3624 c$3626 s$3629 VGND VGND VPWR VPWR c$4012 s$4013 sky130_fd_sc_hd__fa_1
XFILLER_2_774 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4502 net1614 sel_0$6647 net1606 net699 VGND VGND VPWR VPWR t$6705 sky130_fd_sc_hd__a22o_1
XU$$4513 t$6710 net1877 VGND VGND VPWR VPWR booth_b64_m61 sky130_fd_sc_hd__xor2_1
Xdadda_fa_0_61_0 pp_row61_0 pp_row61_1 pp_row61_2 VGND VGND VPWR VPWR c$50 s$51 sky130_fd_sc_hd__fa_2
XU$$16 net1675 net446 net1565 net688 VGND VGND VPWR VPWR t$4415 sky130_fd_sc_hd__a22o_1
XU$$3801 net1701 net474 net1694 net747 VGND VGND VPWR VPWR t$6347 sky130_fd_sc_hd__a22o_1
XTAP_4150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3812 t$6352 net1301 VGND VGND VPWR VPWR booth_b54_m53 sky130_fd_sc_hd__xor2_1
XTAP_4161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_117_2 pp_row117_6 pp_row117_7 c$2748 VGND VGND VPWR VPWR c$3396 s$3397
+ sky130_fd_sc_hd__fa_1
XU$$27 t$4420 net1573 VGND VGND VPWR VPWR booth_b0_m10 sky130_fd_sc_hd__xor2_1
XU$$3823 net1591 net473 net1583 net746 VGND VGND VPWR VPWR t$6358 sky130_fd_sc_hd__a22o_1
XTAP_4172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$38 net1166 net443 net1157 net685 VGND VGND VPWR VPWR t$4426 sky130_fd_sc_hd__a22o_1
XTAP_4183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3834 t$6363 net1308 VGND VGND VPWR VPWR booth_b54_m64 sky130_fd_sc_hd__xor2_1
XU$$49 t$4431 net1575 VGND VGND VPWR VPWR booth_b0_m21 sky130_fd_sc_hd__xor2_1
XU$$3845 t$6370 net1296 VGND VGND VPWR VPWR booth_b56_m1 sky130_fd_sc_hd__xor2_1
XTAP_4194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3856 net1522 net460 net1518 net733 VGND VGND VPWR VPWR t$6376 sky130_fd_sc_hd__a22o_1
XU$$3867 t$6381 net1296 VGND VGND VPWR VPWR booth_b56_m12 sky130_fd_sc_hd__xor2_1
XTAP_3460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3878 net1151 net460 net1141 net733 VGND VGND VPWR VPWR t$6387 sky130_fd_sc_hd__a22o_1
XFILLER_80_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3889 t$6392 net1294 VGND VGND VPWR VPWR booth_b56_m23 sky130_fd_sc_hd__xor2_1
XFILLER_166_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_460 net1674 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_18 sel_0$5177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_29 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0953_ clknet_leaf_114_clk booth_b54_m44 VGND VGND VPWR VPWR pp_row98_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_119_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0884_ clknet_leaf_100_clk booth_b36_m59 VGND VGND VPWR VPWR pp_row95_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_185_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_90_2 pp_row90_17 pp_row90_18 pp_row90_19 VGND VGND VPWR VPWR c$1810 s$1811
+ sky130_fd_sc_hd__fa_1
XFILLER_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_83_1 pp_row83_24 c$922 c$924 VGND VGND VPWR VPWR c$1724 s$1725 sky130_fd_sc_hd__fa_1
XFILLER_47_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1505_ clknet_leaf_122_clk booth_b42_m63 VGND VGND VPWR VPWR pp_row105_1 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_60_0 c$3044 c$3046 c$3048 VGND VGND VPWR VPWR c$3636 s$3637 sky130_fd_sc_hd__fa_1
X_2485_ clknet_leaf_146_clk booth_b12_m57 VGND VGND VPWR VPWR pp_row69_4 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_76_0 s$199 c$798 c$800 VGND VGND VPWR VPWR c$1638 s$1639 sky130_fd_sc_hd__fa_1
XFILLER_114_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1436_ clknet_leaf_41_clk booth_b0_m35 VGND VGND VPWR VPWR pp_row35_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_96_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1367_ clknet_leaf_3_clk booth_b26_m5 VGND VGND VPWR VPWR pp_row31_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_83_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_52_7 pp_row52_23 pp_row52_24 pp_row52_25 VGND VGND VPWR VPWR c$398 s$399
+ sky130_fd_sc_hd__fa_1
X_0318_ clknet_leaf_200_clk booth_b14_m60 VGND VGND VPWR VPWR pp_row74_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1298_ clknet_leaf_251_clk booth_b2_m26 VGND VGND VPWR VPWR pp_row28_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_110_1130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0249_ clknet_leaf_209_clk booth_b8_m64 VGND VGND VPWR VPWR pp_row72_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_71_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2883_1785 VGND VGND VPWR VPWR U$$2883_1785/HI net1785 sky130_fd_sc_hd__conb_1
XFILLER_51_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_98_1 c$2618 c$2620 s$2623 VGND VGND VPWR VPWR c$3280 s$3281 sky130_fd_sc_hd__fa_1
Xdadda_fa_7_75_0 s$3699 c$4044 s$4047 VGND VGND VPWR VPWR c$4302 s$4303 sky130_fd_sc_hd__fa_2
XFILLER_164_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1306 net1308 VGND VGND VPWR VPWR net1306 sky130_fd_sc_hd__buf_6
Xfanout1317 net1318 VGND VGND VPWR VPWR net1317 sky130_fd_sc_hd__buf_6
Xfanout1328 net49 VGND VGND VPWR VPWR net1328 sky130_fd_sc_hd__buf_6
Xfanout1339 net1347 VGND VGND VPWR VPWR net1339 sky130_fd_sc_hd__clkbuf_4
Xfanout385 net386 VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__buf_4
XFILLER_59_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout396 net398 VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__buf_4
XFILLER_87_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3108 net1735 net513 net1727 net786 VGND VGND VPWR VPWR t$5993 sky130_fd_sc_hd__a22o_1
XU$$3119 t$5998 net1364 VGND VGND VPWR VPWR booth_b44_m49 sky130_fd_sc_hd__xor2_1
XFILLER_115_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2407 net975 net565 net966 net838 VGND VGND VPWR VPWR t$5635 sky130_fd_sc_hd__a22o_1
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2418 t$5640 net1425 VGND VGND VPWR VPWR booth_b34_m41 sky130_fd_sc_hd__xor2_1
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2429 net1705 net566 net1697 net839 VGND VGND VPWR VPWR t$5646 sky130_fd_sc_hd__a22o_1
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4381_1809 VGND VGND VPWR VPWR U$$4381_1809/HI net1809 sky130_fd_sc_hd__conb_1
XFILLER_15_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1706 net1057 net605 net1049 net878 VGND VGND VPWR VPWR t$5277 sky130_fd_sc_hd__a22o_1
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1717 t$5282 net1469 VGND VGND VPWR VPWR booth_b24_m33 sky130_fd_sc_hd__xor2_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1728 net949 net607 net941 net880 VGND VGND VPWR VPWR t$5288 sky130_fd_sc_hd__a22o_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1739 t$5293 net1474 VGND VGND VPWR VPWR booth_b24_m44 sky130_fd_sc_hd__xor2_1
XFILLER_188_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput16 a[23] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_8
XFILLER_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput27 a[33] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_1
XFILLER_11_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput38 a[43] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_4
Xinput49 a[53] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_1
XFILLER_182_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_93_0 s$1041 c$1830 c$1832 VGND VGND VPWR VPWR c$2582 s$2583 sky130_fd_sc_hd__fa_1
XFILLER_6_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_848 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2270_ clknet_leaf_210_clk booth_b20_m43 VGND VGND VPWR VPWR pp_row63_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1221_ clknet_leaf_48_clk booth_b10_m13 VGND VGND VPWR VPWR pp_row23_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_111_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4310 t$6607 net1260 VGND VGND VPWR VPWR booth_b62_m28 sky130_fd_sc_hd__xor2_1
XU$$4321 net996 net425 net989 net707 VGND VGND VPWR VPWR t$6613 sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_55_5 s$449 s$451 s$453 VGND VGND VPWR VPWR c$1396 s$1397 sky130_fd_sc_hd__fa_1
XU$$4332 t$6618 net1261 VGND VGND VPWR VPWR booth_b62_m39 sky130_fd_sc_hd__xor2_1
XFILLER_93_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1152_ clknet_leaf_15_clk booth_b10_m8 VGND VGND VPWR VPWR pp_row18_5 sky130_fd_sc_hd__dfxtp_1
XU$$4343 net1727 net423 net1719 net705 VGND VGND VPWR VPWR t$6624 sky130_fd_sc_hd__a22o_1
XU$$4354 t$6629 net1255 VGND VGND VPWR VPWR booth_b62_m50 sky130_fd_sc_hd__xor2_1
XFILLER_65_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_48_4 s$319 s$321 s$323 VGND VGND VPWR VPWR c$1310 s$1311 sky130_fd_sc_hd__fa_1
XU$$3620 net1076 net476 net1068 net749 VGND VGND VPWR VPWR t$6255 sky130_fd_sc_hd__a22o_1
XU$$4365 net1617 net420 net1610 net702 VGND VGND VPWR VPWR t$6635 sky130_fd_sc_hd__a22o_1
XU$$3631 t$6260 net1323 VGND VGND VPWR VPWR booth_b52_m31 sky130_fd_sc_hd__xor2_1
XU$$4376 t$6640 net1257 VGND VGND VPWR VPWR booth_b62_m61 sky130_fd_sc_hd__xor2_1
XFILLER_19_962 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3642 net967 net478 net958 net751 VGND VGND VPWR VPWR t$6266 sky130_fd_sc_hd__a22o_1
XU$$4387 net1812 notblock$6645\[1\] VGND VGND VPWR VPWR t$6646 sky130_fd_sc_hd__and2_1
XU$$4398 net939 sel_0$6647 net1678 net698 VGND VGND VPWR VPWR t$6653 sky130_fd_sc_hd__a22o_1
X_1083_ clknet_leaf_120_clk booth_b52_m50 VGND VGND VPWR VPWR pp_row102_8 sky130_fd_sc_hd__dfxtp_1
XU$$3653 t$6271 net1325 VGND VGND VPWR VPWR booth_b52_m42 sky130_fd_sc_hd__xor2_1
XU$$3664 net1701 net482 net1694 net755 VGND VGND VPWR VPWR t$6277 sky130_fd_sc_hd__a22o_1
XU$$2930 t$5902 net1372 VGND VGND VPWR VPWR booth_b42_m23 sky130_fd_sc_hd__xor2_1
XU$$3675 t$6282 net1326 VGND VGND VPWR VPWR booth_b52_m53 sky130_fd_sc_hd__xor2_1
XFILLER_34_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2941 net1051 net520 net1043 net793 VGND VGND VPWR VPWR t$5908 sky130_fd_sc_hd__a22o_1
XU$$3686 net1591 net483 net1583 net756 VGND VGND VPWR VPWR t$6288 sky130_fd_sc_hd__a22o_1
XU$$2952 t$5913 net1370 VGND VGND VPWR VPWR booth_b42_m34 sky130_fd_sc_hd__xor2_1
XU$$3697 t$6293 net1321 VGND VGND VPWR VPWR booth_b52_m64 sky130_fd_sc_hd__xor2_1
XTAP_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2963 net942 net521 net926 net794 VGND VGND VPWR VPWR t$5919 sky130_fd_sc_hd__a22o_1
XU$$2974 t$5924 net1369 VGND VGND VPWR VPWR booth_b42_m45 sky130_fd_sc_hd__xor2_1
XU$$2985 net1660 net524 net1652 net797 VGND VGND VPWR VPWR t$5930 sky130_fd_sc_hd__a22o_1
XU$$2996 t$5935 net1373 VGND VGND VPWR VPWR booth_b42_m56 sky130_fd_sc_hd__xor2_1
XFILLER_21_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_290 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1985_ clknet_leaf_79_clk booth_b8_m47 VGND VGND VPWR VPWR pp_row55_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_193_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0936_ clknet_leaf_104_clk booth_b58_m39 VGND VGND VPWR VPWR pp_row97_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0867_ clknet_leaf_111_clk booth_b42_m52 VGND VGND VPWR VPWR pp_row94_7 sky130_fd_sc_hd__dfxtp_1
X_0798_ clknet_leaf_123_clk booth_b38_m53 VGND VGND VPWR VPWR pp_row91_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_115_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2468_ clknet_leaf_102_clk booth_b46_m22 VGND VGND VPWR VPWR pp_row68_22 sky130_fd_sc_hd__dfxtp_1
Xdadda_ha_1_44_5 pp_row44_15 pp_row44_16 VGND VGND VPWR VPWR c$274 s$275 sky130_fd_sc_hd__ha_1
XFILLER_88_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$903 final_adder.$signal$1206 final_adder.g_new$975 final_adder.$signal$234
+ VGND VGND VPWR VPWR final_adder.g_new$1031 sky130_fd_sc_hd__a21o_1
X_1419_ clknet_leaf_56_clk booth_b8_m26 VGND VGND VPWR VPWR pp_row34_4 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$914 final_adder.$signal$1184 final_adder.g_new$997 final_adder.$signal$190
+ VGND VGND VPWR VPWR final_adder.g_new$1042 sky130_fd_sc_hd__a21o_1
X_2399_ clknet_leaf_74_clk booth_b52_m14 VGND VGND VPWR VPWR pp_row66_26 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$925 final_adder.$signal$1162 final_adder.g_new$1019 final_adder.$signal$146
+ VGND VGND VPWR VPWR final_adder.g_new$1053 sky130_fd_sc_hd__a21o_1
XFILLER_69_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$936 final_adder.$signal$103 final_adder.g_new$945 final_adder.$signal$102
+ VGND VGND VPWR VPWR final_adder.g_new$1064 sky130_fd_sc_hd__a21o_1
Xdadda_fa_1_50_4 pp_row50_12 pp_row50_13 pp_row50_14 VGND VGND VPWR VPWR c$356 s$357
+ sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$947 final_adder.$signal$1118 final_adder.g_new$855 final_adder.$signal$58
+ VGND VGND VPWR VPWR final_adder.g_new$1075 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$958 final_adder.$signal$1096 final_adder.g_new$633 final_adder.$signal$14
+ VGND VGND VPWR VPWR final_adder.g_new$1086 sky130_fd_sc_hd__a21o_1
XU$$808 t$4817 net1419 VGND VGND VPWR VPWR booth_b10_m58 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$969 final_adder.$signal$1098 final_adder.g_new$631 VGND VGND VPWR
+ VPWR net373 sky130_fd_sc_hd__xor2_2
XU$$819 net1527 net403 net1886 net669 VGND VGND VPWR VPWR t$4823 sky130_fd_sc_hd__a22o_1
XFILLER_83_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_43_3 pp_row43_9 pp_row43_10 pp_row43_11 VGND VGND VPWR VPWR c$260 s$261
+ sky130_fd_sc_hd__fa_1
XFILLER_28_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_20_2 s$2001 s$2003 s$2005 VGND VGND VPWR VPWR c$2814 s$2815 sky130_fd_sc_hd__fa_1
XFILLER_71_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_13_1 pp_row13_3 pp_row13_4 pp_row13_5 VGND VGND VPWR VPWR c$2770 s$2771
+ sky130_fd_sc_hd__fa_1
XFILLER_52_773 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1103 net1104 VGND VGND VPWR VPWR net1103 sky130_fd_sc_hd__buf_4
Xfanout1114 net1116 VGND VGND VPWR VPWR net1114 sky130_fd_sc_hd__buf_4
Xfanout1125 net76 VGND VGND VPWR VPWR net1125 sky130_fd_sc_hd__buf_4
Xfanout1136 net1137 VGND VGND VPWR VPWR net1136 sky130_fd_sc_hd__buf_6
XFILLER_66_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1147 net1154 VGND VGND VPWR VPWR net1147 sky130_fd_sc_hd__buf_4
Xfanout1158 net72 VGND VGND VPWR VPWR net1158 sky130_fd_sc_hd__buf_4
Xdadda_fa_3_58_3 s$1427 s$1429 s$1431 VGND VGND VPWR VPWR c$2308 s$2309 sky130_fd_sc_hd__fa_1
XFILLER_47_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1169 net71 VGND VGND VPWR VPWR net1169 sky130_fd_sc_hd__clkbuf_2
XFILLER_102_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2204 net1038 net572 net937 net845 VGND VGND VPWR VPWR t$5532 sky130_fd_sc_hd__a22o_1
XFILLER_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2215 t$5537 net1430 VGND VGND VPWR VPWR booth_b32_m8 sky130_fd_sc_hd__xor2_1
XFILLER_170_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2226 net1193 net569 net1174 net842 VGND VGND VPWR VPWR t$5543 sky130_fd_sc_hd__a22o_1
XU$$2237 t$5548 net1432 VGND VGND VPWR VPWR booth_b32_m19 sky130_fd_sc_hd__xor2_1
XU$$1503 t$5172 net1491 VGND VGND VPWR VPWR booth_b20_m63 sky130_fd_sc_hd__xor2_1
XFILLER_76_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2248 net1083 net570 net1074 net843 VGND VGND VPWR VPWR t$5554 sky130_fd_sc_hd__a22o_1
XFILLER_188_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2259 t$5559 net1431 VGND VGND VPWR VPWR booth_b32_m30 sky130_fd_sc_hd__xor2_1
XU$$1514 t$5179 net1478 VGND VGND VPWR VPWR booth_b22_m0 sky130_fd_sc_hd__xor2_1
XU$$1525 net1560 net610 net1519 net883 VGND VGND VPWR VPWR t$5185 sky130_fd_sc_hd__a22o_1
XFILLER_90_879 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1536 t$5190 net1479 VGND VGND VPWR VPWR booth_b22_m11 sky130_fd_sc_hd__xor2_1
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_21__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_5_21__leaf_clk sky130_fd_sc_hd__clkbuf_16
XU$$1547 net1157 net610 net1147 net883 VGND VGND VPWR VPWR t$5196 sky130_fd_sc_hd__a22o_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1558 t$5201 net1477 VGND VGND VPWR VPWR booth_b22_m22 sky130_fd_sc_hd__xor2_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1569 net1057 net613 net1049 net886 VGND VGND VPWR VPWR t$5207 sky130_fd_sc_hd__a22o_1
XFILLER_15_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1770_ clknet_leaf_238_clk booth_b12_m36 VGND VGND VPWR VPWR pp_row48_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_184_951 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0721_ clknet_leaf_132_clk booth_b56_m62 VGND VGND VPWR VPWR pp_row118_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_128_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0652_ clknet_leaf_169_clk booth_b38_m47 VGND VGND VPWR VPWR pp_row85_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_171_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0583_ clknet_leaf_173_clk booth_b60_m22 VGND VGND VPWR VPWR pp_row82_22 sky130_fd_sc_hd__dfxtp_1
XFILLER_170_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2322_ clknet_leaf_77_clk booth_b46_m18 VGND VGND VPWR VPWR pp_row64_23 sky130_fd_sc_hd__dfxtp_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_2_60_3 c$526 s$529 s$531 VGND VGND VPWR VPWR c$1452 s$1453 sky130_fd_sc_hd__fa_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2253_ clknet_leaf_150_clk booth_b56_m6 VGND VGND VPWR VPWR pp_row62_28 sky130_fd_sc_hd__dfxtp_1
XFILLER_85_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_53_2 c$394 c$396 c$398 VGND VGND VPWR VPWR c$1366 s$1367 sky130_fd_sc_hd__fa_1
Xfanout1670 net11 VGND VGND VPWR VPWR net1670 sky130_fd_sc_hd__buf_6
X_1204_ clknet_leaf_51_clk booth_b8_m14 VGND VGND VPWR VPWR pp_row22_4 sky130_fd_sc_hd__dfxtp_1
Xfanout1681 net108 VGND VGND VPWR VPWR net1681 sky130_fd_sc_hd__buf_6
XU$$4140 net1214 net434 net1205 net716 VGND VGND VPWR VPWR t$6521 sky130_fd_sc_hd__a22o_1
XFILLER_38_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2184_ clknet_leaf_216_clk booth_b60_m0 VGND VGND VPWR VPWR pp_row60_30 sky130_fd_sc_hd__dfxtp_1
Xfanout1692 net1694 VGND VGND VPWR VPWR net1692 sky130_fd_sc_hd__buf_6
Xdadda_fa_5_30_1 s$2871 s$2873 s$2875 VGND VGND VPWR VPWR c$3518 s$3519 sky130_fd_sc_hd__fa_1
XU$$4151 t$6526 net1267 VGND VGND VPWR VPWR booth_b60_m17 sky130_fd_sc_hd__xor2_1
XFILLER_66_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_46_1 pp_row46_23 pp_row46_24 pp_row46_25 VGND VGND VPWR VPWR c$1280 s$1281
+ sky130_fd_sc_hd__fa_1
XU$$4162 net1103 net436 net1095 net718 VGND VGND VPWR VPWR t$6532 sky130_fd_sc_hd__a22o_1
XFILLER_65_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1135_ clknet_leaf_16_clk booth_b0_m17 VGND VGND VPWR VPWR pp_row17_0 sky130_fd_sc_hd__dfxtp_1
XU$$4173 t$6537 net1265 VGND VGND VPWR VPWR booth_b60_m28 sky130_fd_sc_hd__xor2_1
XFILLER_25_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_23_0 c$2822 c$2824 c$2826 VGND VGND VPWR VPWR c$3488 s$3489 sky130_fd_sc_hd__fa_1
XU$$4184 net996 net441 net988 net723 VGND VGND VPWR VPWR t$6543 sky130_fd_sc_hd__a22o_1
XU$$4195 t$6548 net1271 VGND VGND VPWR VPWR booth_b60_m39 sky130_fd_sc_hd__xor2_1
XU$$3450 t$6168 net1329 VGND VGND VPWR VPWR booth_b50_m9 sky130_fd_sc_hd__xor2_1
XU$$3461 net1181 net488 net1172 net761 VGND VGND VPWR VPWR t$6174 sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_39_0 pp_row39_8 pp_row39_9 pp_row39_10 VGND VGND VPWR VPWR c$1194 s$1195
+ sky130_fd_sc_hd__fa_1
XU$$3472 t$6179 net1330 VGND VGND VPWR VPWR booth_b50_m20 sky130_fd_sc_hd__xor2_1
XFILLER_92_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1066_ clknet_leaf_248_clk net256 VGND VGND VPWR VPWR pp_row9_5 sky130_fd_sc_hd__dfxtp_2
XFILLER_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3483 net1076 net484 net1068 net757 VGND VGND VPWR VPWR t$6185 sky130_fd_sc_hd__a22o_1
XU$$3494 t$6190 net1331 VGND VGND VPWR VPWR booth_b50_m31 sky130_fd_sc_hd__xor2_1
XU$$2760 net1522 net535 net1514 net808 VGND VGND VPWR VPWR t$5816 sky130_fd_sc_hd__a22o_1
XU$$2771 t$5821 net1381 VGND VGND VPWR VPWR booth_b40_m12 sky130_fd_sc_hd__xor2_1
XFILLER_34_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2782 net1151 net536 net1141 net809 VGND VGND VPWR VPWR t$5827 sky130_fd_sc_hd__a22o_1
XFILLER_21_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2793 t$5832 net1380 VGND VGND VPWR VPWR booth_b40_m23 sky130_fd_sc_hd__xor2_1
XU$$4405_1823 VGND VGND VPWR VPWR U$$4405_1823/HI net1823 sky130_fd_sc_hd__conb_1
XFILLER_178_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1968_ clknet_leaf_62_clk booth_b38_m16 VGND VGND VPWR VPWR pp_row54_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_30_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0919_ clknet_leaf_111_clk booth_b64_m32 VGND VGND VPWR VPWR pp_row96_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1899_ clknet_leaf_63_clk booth_b28_m24 VGND VGND VPWR VPWR pp_row52_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_119_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_68_2 s$2385 s$2387 s$2389 VGND VGND VPWR VPWR c$3102 s$3103 sky130_fd_sc_hd__fa_1
XFILLER_88_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput206 c[54] VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkbuf_1
XFILLER_103_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput217 c[64] VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__clkbuf_1
Xinput228 c[74] VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput239 c[84] VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__clkbuf_1
XFILLER_57_810 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$700 final_adder.p_new$724 final_adder.p_new$708 VGND VGND VPWR VPWR
+ final_adder.p_new$828 sky130_fd_sc_hd__and2_1
XFILLER_124_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_38_0 s$3551 c$3970 s$3973 VGND VGND VPWR VPWR c$4228 s$4229 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$711 final_adder.p_new$718 final_adder.g_new$735 final_adder.g_new$719
+ VGND VGND VPWR VPWR final_adder.g_new$839 sky130_fd_sc_hd__a21o_1
XFILLER_25_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$733 final_adder.p_new$740 final_adder.g_new$633 final_adder.g_new$741
+ VGND VGND VPWR VPWR final_adder.g_new$861 sky130_fd_sc_hd__a21o_2
Xfinal_adder.U$$744 final_adder.p_new$792 final_adder.p_new$760 VGND VGND VPWR VPWR
+ final_adder.p_new$872 sky130_fd_sc_hd__and2_1
XFILLER_5_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$755 final_adder.p_new$770 final_adder.g_new$803 final_adder.g_new$771
+ VGND VGND VPWR VPWR final_adder.g_new$883 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$766 final_adder.p_new$814 final_adder.p_new$782 VGND VGND VPWR VPWR
+ final_adder.p_new$894 sky130_fd_sc_hd__and2_1
XU$$605 t$4714 net1239 VGND VGND VPWR VPWR booth_b8_m25 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$777 final_adder.p_new$792 final_adder.g_new$825 final_adder.g_new$793
+ VGND VGND VPWR VPWR final_adder.g_new$905 sky130_fd_sc_hd__a21o_1
XFILLER_72_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$616 net1025 net415 net1017 net681 VGND VGND VPWR VPWR t$4720 sky130_fd_sc_hd__a22o_1
Xdadda_fa_1_41_0 pp_row41_0 pp_row41_1 pp_row41_2 VGND VGND VPWR VPWR c$236 s$237
+ sky130_fd_sc_hd__fa_1
XU$$627 t$4725 net1236 VGND VGND VPWR VPWR booth_b8_m36 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$788 final_adder.p_new$836 final_adder.p_new$804 VGND VGND VPWR VPWR
+ final_adder.p_new$916 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$799 final_adder.p_new$814 final_adder.g_new$847 final_adder.g_new$815
+ VGND VGND VPWR VPWR final_adder.g_new$927 sky130_fd_sc_hd__a21o_1
XU$$638 net1745 net411 net1737 net677 VGND VGND VPWR VPWR t$4731 sky130_fd_sc_hd__a22o_1
XFILLER_71_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1028 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$649 t$4736 net1242 VGND VGND VPWR VPWR booth_b8_m47 sky130_fd_sc_hd__xor2_1
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_848 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_70_2 c$1564 s$1567 s$1569 VGND VGND VPWR VPWR c$2402 s$2403 sky130_fd_sc_hd__fa_1
XFILLER_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_63_1 c$1474 c$1476 c$1478 VGND VGND VPWR VPWR c$2344 s$2345 sky130_fd_sc_hd__fa_1
Xdadda_fa_6_40_0 c$3552 c$3554 s$3557 VGND VGND VPWR VPWR c$3976 s$3977 sky130_fd_sc_hd__fa_1
XFILLER_181_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_56_0 s$473 c$1386 c$1388 VGND VGND VPWR VPWR c$2286 s$2287 sky130_fd_sc_hd__fa_1
XFILLER_75_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2001 t$5427 net1452 VGND VGND VPWR VPWR booth_b28_m38 sky130_fd_sc_hd__xor2_1
XFILLER_47_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2012 net1730 net589 net1721 net862 VGND VGND VPWR VPWR t$5433 sky130_fd_sc_hd__a22o_1
XU$$2023 t$5438 net1455 VGND VGND VPWR VPWR booth_b28_m49 sky130_fd_sc_hd__xor2_1
XU$$2034 net1622 net589 net1613 net862 VGND VGND VPWR VPWR t$5444 sky130_fd_sc_hd__a22o_1
XU$$1300 t$5069 net1663 VGND VGND VPWR VPWR booth_b18_m30 sky130_fd_sc_hd__xor2_1
XU$$2045 t$5449 net1455 VGND VGND VPWR VPWR booth_b28_m60 sky130_fd_sc_hd__xor2_1
XU$$1311 net978 net638 net972 net911 VGND VGND VPWR VPWR t$5075 sky130_fd_sc_hd__a22o_1
XFILLER_16_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2056 net24 VGND VGND VPWR VPWR notblock$5455\[1\] sky130_fd_sc_hd__inv_1
XFILLER_63_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1322 t$5080 net1669 VGND VGND VPWR VPWR booth_b18_m41 sky130_fd_sc_hd__xor2_1
XU$$2067 net1036 net581 net936 net854 VGND VGND VPWR VPWR t$5462 sky130_fd_sc_hd__a22o_1
XU$$2078 t$5467 net1439 VGND VGND VPWR VPWR booth_b30_m8 sky130_fd_sc_hd__xor2_1
XFILLER_16_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1333 net1706 net642 net1698 net915 VGND VGND VPWR VPWR t$5086 sky130_fd_sc_hd__a22o_1
XFILLER_188_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2089 net1195 net577 net1175 net850 VGND VGND VPWR VPWR t$5473 sky130_fd_sc_hd__a22o_1
XU$$1344 t$5091 net1670 VGND VGND VPWR VPWR booth_b18_m52 sky130_fd_sc_hd__xor2_1
XU$$1355 net1595 net640 net1586 net913 VGND VGND VPWR VPWR t$5097 sky130_fd_sc_hd__a22o_1
XU$$1366 t$5102 net1669 VGND VGND VPWR VPWR booth_b18_m63 sky130_fd_sc_hd__xor2_1
XU$$1377 t$5109 net1487 VGND VGND VPWR VPWR booth_b20_m0 sky130_fd_sc_hd__xor2_1
XU$$1388 net1560 net627 net1519 net900 VGND VGND VPWR VPWR t$5115 sky130_fd_sc_hd__a22o_1
XFILLER_128_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1399 t$5120 net1485 VGND VGND VPWR VPWR booth_b20_m11 sky130_fd_sc_hd__xor2_1
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1822_ clknet_leaf_232_clk booth_b0_m50 VGND VGND VPWR VPWR pp_row50_0 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_7_113_0 s$3851 c$4120 s$4123 VGND VGND VPWR VPWR c$4378 s$4379 sky130_fd_sc_hd__fa_1
XFILLER_157_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1753_ clknet_leaf_223_clk booth_b30_m17 VGND VGND VPWR VPWR pp_row47_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_144_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0704_ clknet_leaf_170_clk booth_b40_m47 VGND VGND VPWR VPWR pp_row87_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_116_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1684_ clknet_leaf_19_clk booth_b6_m39 VGND VGND VPWR VPWR pp_row45_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_132_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_78_1 s$3159 s$3161 s$3163 VGND VGND VPWR VPWR c$3710 s$3711 sky130_fd_sc_hd__fa_1
XFILLER_89_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0635_ clknet_leaf_174_clk booth_b54_m30 VGND VGND VPWR VPWR pp_row84_18 sky130_fd_sc_hd__dfxtp_1
XU$$4435_1838 VGND VGND VPWR VPWR U$$4435_1838/HI net1838 sky130_fd_sc_hd__conb_1
XFILLER_143_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout907 sel_1$5108 VGND VGND VPWR VPWR net907 sky130_fd_sc_hd__buf_6
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout918 net919 VGND VGND VPWR VPWR net918 sky130_fd_sc_hd__clkbuf_8
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0566_ clknet_leaf_126_clk booth_b58_m58 VGND VGND VPWR VPWR pp_row116_4 sky130_fd_sc_hd__dfxtp_1
Xfanout929 net930 VGND VGND VPWR VPWR net929 sky130_fd_sc_hd__clkbuf_8
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_607 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2305_ clknet_leaf_133_clk booth_b64_m46 VGND VGND VPWR VPWR pp_row110_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_135_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0497_ clknet_leaf_158_clk booth_b60_m19 VGND VGND VPWR VPWR pp_row79_23 sky130_fd_sc_hd__dfxtp_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2236_ clknet_leaf_228_clk booth_b26_m36 VGND VGND VPWR VPWR pp_row62_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_39_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2167_ clknet_leaf_27_clk booth_b32_m28 VGND VGND VPWR VPWR pp_row60_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_94_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1118_ clknet_leaf_14_clk booth_b8_m7 VGND VGND VPWR VPWR pp_row15_4 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$40 c$4230 s$4233 VGND VGND VPWR VPWR final_adder.$signal$82 final_adder.$signal$1130
+ sky130_fd_sc_hd__ha_2
X_2098_ clknet_leaf_86_clk booth_b32_m26 VGND VGND VPWR VPWR pp_row58_16 sky130_fd_sc_hd__dfxtp_1
XU$$3280 t$6080 net1356 VGND VGND VPWR VPWR booth_b46_m61 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$51 c$4252 s$4255 VGND VGND VPWR VPWR final_adder.$signal$104 final_adder.$signal$105
+ sky130_fd_sc_hd__ha_1
XU$$3291 net1340 notblock$6085\[1\] VGND VGND VPWR VPWR t$6086 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$62 c$4274 s$4277 VGND VGND VPWR VPWR final_adder.$signal$126 final_adder.$signal$1152
+ sky130_fd_sc_hd__ha_2
XFILLER_0_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$73 c$4296 s$4299 VGND VGND VPWR VPWR final_adder.$signal$148 final_adder.$signal$1163
+ sky130_fd_sc_hd__ha_1
XFILLER_13_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$84 c$4318 s$4321 VGND VGND VPWR VPWR final_adder.$signal$170 final_adder.$signal$1174
+ sky130_fd_sc_hd__ha_1
X_1049_ clknet_leaf_120_clk booth_b46_m56 VGND VGND VPWR VPWR pp_row102_5 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$95 c$4340 s$4343 VGND VGND VPWR VPWR final_adder.$signal$192 final_adder.$signal$1185
+ sky130_fd_sc_hd__ha_1
XFILLER_94_1072 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2590 net1593 net557 net1585 net830 VGND VGND VPWR VPWR t$5728 sky130_fd_sc_hd__a22o_1
XFILLER_34_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_80_1 c$2474 c$2476 s$2479 VGND VGND VPWR VPWR c$3172 s$3173 sky130_fd_sc_hd__fa_1
XFILLER_150_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_73_0 s$1613 c$2414 c$2416 VGND VGND VPWR VPWR c$3128 s$3129 sky130_fd_sc_hd__fa_1
Xdadda_fa_1_89_0 pp_row89_0 pp_row89_1 pp_row89_2 VGND VGND VPWR VPWR c$1010 s$1011
+ sky130_fd_sc_hd__fa_2
XFILLER_135_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$530 final_adder.p_new$542 final_adder.p_new$534 VGND VGND VPWR VPWR
+ final_adder.p_new$658 sky130_fd_sc_hd__and2_1
XTAP_3812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$541 final_adder.p_new$544 final_adder.g_new$553 final_adder.g_new$545
+ VGND VGND VPWR VPWR final_adder.g_new$669 sky130_fd_sc_hd__a21o_1
XTAP_3823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$552 final_adder.p_new$564 final_adder.p_new$556 VGND VGND VPWR VPWR
+ final_adder.p_new$680 sky130_fd_sc_hd__and2_1
XTAP_3834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$402 net1555 net533 net1547 net806 VGND VGND VPWR VPWR t$4610 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$563 final_adder.p_new$566 final_adder.g_new$575 final_adder.g_new$567
+ VGND VGND VPWR VPWR final_adder.g_new$691 sky130_fd_sc_hd__a21o_1
XTAP_3845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$413 net1246 VGND VGND VPWR VPWR notblock$4615\[2\] sky130_fd_sc_hd__inv_1
XFILLER_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$574 final_adder.p_new$586 final_adder.p_new$578 VGND VGND VPWR VPWR
+ final_adder.p_new$702 sky130_fd_sc_hd__and2_1
XTAP_3856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$585 final_adder.p_new$588 final_adder.g_new$597 final_adder.g_new$589
+ VGND VGND VPWR VPWR final_adder.g_new$713 sky130_fd_sc_hd__a21o_1
XU$$424 t$4622 net1248 VGND VGND VPWR VPWR booth_b6_m3 sky130_fd_sc_hd__xor2_1
XTAP_3867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$435 net1505 net431 net1496 net713 VGND VGND VPWR VPWR t$4628 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$596 final_adder.p_new$608 final_adder.p_new$600 VGND VGND VPWR VPWR
+ final_adder.p_new$724 sky130_fd_sc_hd__and2_1
XTAP_3878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$446 t$4633 net1249 VGND VGND VPWR VPWR booth_b6_m14 sky130_fd_sc_hd__xor2_1
XFILLER_189_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$457 net1130 net426 net1114 net708 VGND VGND VPWR VPWR t$4639 sky130_fd_sc_hd__a22o_1
XU$$468 t$4644 net1245 VGND VGND VPWR VPWR booth_b6_m25 sky130_fd_sc_hd__xor2_1
XU$$479 net1025 net431 net1017 net713 VGND VGND VPWR VPWR t$4650 sky130_fd_sc_hd__a22o_1
XFILLER_44_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_160_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_160_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_154_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_88_0 c$3744 c$3746 s$3749 VGND VGND VPWR VPWR c$4072 s$4073 sky130_fd_sc_hd__fa_2
XFILLER_5_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_0_78_0 net1915 pp_row78_1 VGND VGND VPWR VPWR c$202 s$203 sky130_fd_sc_hd__ha_1
XFILLER_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0420_ clknet_leaf_145_clk booth_b28_m49 VGND VGND VPWR VPWR pp_row77_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_69_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0351_ clknet_leaf_200_clk booth_b16_m59 VGND VGND VPWR VPWR pp_row75_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_121_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0282_ clknet_leaf_198_clk net226 VGND VGND VPWR VPWR pp_row72_30 sky130_fd_sc_hd__dfxtp_1
XFILLER_36_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2021_ clknet_leaf_33_clk booth_b16_m40 VGND VGND VPWR VPWR pp_row56_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_35_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$980 t$4906 net1187 VGND VGND VPWR VPWR booth_b14_m7 sky130_fd_sc_hd__xor2_1
XFILLER_35_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$991 net1201 net385 net1192 net651 VGND VGND VPWR VPWR t$4912 sky130_fd_sc_hd__a22o_1
XU$$1130 net1192 net643 net1173 net916 VGND VGND VPWR VPWR t$4983 sky130_fd_sc_hd__a22o_1
XFILLER_165_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1141 t$4988 net1010 VGND VGND VPWR VPWR booth_b16_m19 sky130_fd_sc_hd__xor2_1
XU$$1152 net1080 net644 net1071 net917 VGND VGND VPWR VPWR t$4994 sky130_fd_sc_hd__a22o_1
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1163 t$4999 net1007 VGND VGND VPWR VPWR booth_b16_m30 sky130_fd_sc_hd__xor2_1
XU$$1174 net977 net645 net969 net918 VGND VGND VPWR VPWR t$5005 sky130_fd_sc_hd__a22o_1
XFILLER_189_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1185 t$5010 net1011 VGND VGND VPWR VPWR booth_b16_m41 sky130_fd_sc_hd__xor2_1
XFILLER_149_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1196 net1703 net648 net1695 net921 VGND VGND VPWR VPWR t$5016 sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_151_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_151_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_176_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1805_ clknet_leaf_141_clk booth_b44_m63 VGND VGND VPWR VPWR pp_row107_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_129_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_90_0 c$3224 c$3226 c$3228 VGND VGND VPWR VPWR c$3756 s$3757 sky130_fd_sc_hd__fa_2
XFILLER_191_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1736_ clknet_leaf_236_clk booth_b0_m47 VGND VGND VPWR VPWR pp_row47_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_172_773 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1667_ clknet_leaf_21_clk booth_b26_m18 VGND VGND VPWR VPWR pp_row44_13 sky130_fd_sc_hd__dfxtp_1
X_0618_ clknet_leaf_187_clk booth_b24_m60 VGND VGND VPWR VPWR pp_row84_3 sky130_fd_sc_hd__dfxtp_1
Xfanout704 net707 VGND VGND VPWR VPWR net704 sky130_fd_sc_hd__buf_4
Xfanout715 sel_1$4618 VGND VGND VPWR VPWR net715 sky130_fd_sc_hd__buf_6
X_1598_ clknet_leaf_5_clk booth_b40_m1 VGND VGND VPWR VPWR pp_row41_20 sky130_fd_sc_hd__dfxtp_1
Xfanout726 net727 VGND VGND VPWR VPWR net726 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_75_6 pp_row75_24 pp_row75_25 pp_row75_26 VGND VGND VPWR VPWR c$810 s$811
+ sky130_fd_sc_hd__fa_1
XFILLER_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout737 net740 VGND VGND VPWR VPWR net737 sky130_fd_sc_hd__clkbuf_8
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0549_ clknet_leaf_171_clk booth_b48_m33 VGND VGND VPWR VPWR pp_row81_16 sky130_fd_sc_hd__dfxtp_1
Xfanout748 sel_1$6298 VGND VGND VPWR VPWR net748 sky130_fd_sc_hd__buf_6
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout759 net760 VGND VGND VPWR VPWR net759 sky130_fd_sc_hd__clkbuf_4
XFILLER_105_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_68_5 pp_row68_32 c$120 c$122 VGND VGND VPWR VPWR c$682 s$683 sky130_fd_sc_hd__fa_1
XFILLER_140_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2219_ clknet_leaf_216_clk booth_b58_m3 VGND VGND VPWR VPWR pp_row61_29 sky130_fd_sc_hd__dfxtp_1
XFILLER_2_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_108 net602 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_119 net644 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_142_clk clknet_5_25__leaf_clk VGND VGND VPWR VPWR clknet_leaf_142_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_10_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_120_0 c$3872 c$3874 s$3877 VGND VGND VPWR VPWR c$4136 s$4137 sky130_fd_sc_hd__fa_1
XTAP_4310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_63_4 pp_row63_12 pp_row63_13 pp_row63_14 VGND VGND VPWR VPWR c$80 s$81
+ sky130_fd_sc_hd__fa_1
XTAP_4332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_40_3 s$1211 s$1213 s$1215 VGND VGND VPWR VPWR c$2164 s$2165 sky130_fd_sc_hd__fa_1
XTAP_4365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$360 final_adder.p_new$362 final_adder.p_new$360 VGND VGND VPWR VPWR
+ final_adder.p_new$488 sky130_fd_sc_hd__and2_1
XTAP_3642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$371 final_adder.p_new$370 final_adder.g_new$373 final_adder.g_new$371
+ VGND VGND VPWR VPWR final_adder.g_new$499 sky130_fd_sc_hd__a21o_1
XU$$210 t$4512 net1389 VGND VGND VPWR VPWR booth_b2_m33 sky130_fd_sc_hd__xor2_1
XTAP_4387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$221 net948 net619 net940 net892 VGND VGND VPWR VPWR t$4518 sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_33_2 c$1120 s$1123 s$1125 VGND VGND VPWR VPWR c$2106 s$2107 sky130_fd_sc_hd__fa_1
XTAP_4398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$393 final_adder.p_new$394 final_adder.g_new$399 final_adder.g_new$395
+ VGND VGND VPWR VPWR final_adder.g_new$521 sky130_fd_sc_hd__a21o_1
XU$$232 t$4523 net1386 VGND VGND VPWR VPWR booth_b2_m44 sky130_fd_sc_hd__xor2_1
XTAP_3675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$243 net1683 net626 net1658 net899 VGND VGND VPWR VPWR t$4529 sky130_fd_sc_hd__a22o_1
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$254 t$4534 net1392 VGND VGND VPWR VPWR booth_b2_m55 sky130_fd_sc_hd__xor2_1
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$265 net1551 net621 net1543 net894 VGND VGND VPWR VPWR t$4540 sky130_fd_sc_hd__a22o_1
XFILLER_44_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_26_1 pp_row26_11 pp_row26_12 pp_row26_13 VGND VGND VPWR VPWR c$2048 s$2049
+ sky130_fd_sc_hd__fa_1
XFILLER_73_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$276 net1275 VGND VGND VPWR VPWR notblock$4545\[2\] sky130_fd_sc_hd__inv_1
XFILLER_72_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$287 t$4552 net1277 VGND VGND VPWR VPWR booth_b4_m3 sky130_fd_sc_hd__xor2_1
XTAP_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$298 net1509 net531 net1500 net804 VGND VGND VPWR VPWR t$4558 sky130_fd_sc_hd__a22o_1
XTAP_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_19_0 pp_row19_0 pp_row19_1 pp_row19_2 VGND VGND VPWR VPWR c$1992 s$1993
+ sky130_fd_sc_hd__fa_1
XTAP_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_133_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_133_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_139_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4 notblock\[2\] net1 net1802 t notblock\[0\] VGND VGND VPWR VPWR sel_0 sky130_fd_sc_hd__a32o_1
Xoutput307 net307 VGND VGND VPWR VPWR o[2] sky130_fd_sc_hd__buf_2
Xoutput318 net318 VGND VGND VPWR VPWR o[3] sky130_fd_sc_hd__buf_2
X_1521_ clknet_leaf_246_clk booth_b32_m6 VGND VGND VPWR VPWR pp_row38_16 sky130_fd_sc_hd__dfxtp_1
Xoutput329 net329 VGND VGND VPWR VPWR o[4] sky130_fd_sc_hd__buf_2
XFILLER_113_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_85_5 s$971 s$973 s$975 VGND VGND VPWR VPWR c$1756 s$1757 sky130_fd_sc_hd__fa_2
XFILLER_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1452_ clknet_leaf_64_clk booth_b28_m7 VGND VGND VPWR VPWR pp_row35_14 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_78_4 s$857 s$859 s$861 VGND VGND VPWR VPWR c$1670 s$1671 sky130_fd_sc_hd__fa_1
X_0403_ clknet_leaf_208_clk booth_b52_m24 VGND VGND VPWR VPWR pp_row76_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_171_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1383_ clknet_leaf_44_clk booth_b20_m12 VGND VGND VPWR VPWR pp_row32_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_68_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0334_ clknet_leaf_225_clk booth_b42_m32 VGND VGND VPWR VPWR pp_row74_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_110_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0265_ clknet_leaf_150_clk booth_b38_m34 VGND VGND VPWR VPWR pp_row72_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_82_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2004_ clknet_leaf_74_clk booth_b44_m11 VGND VGND VPWR VPWR pp_row55_22 sky130_fd_sc_hd__dfxtp_1
X_0196_ clknet_leaf_154_clk booth_b34_m36 VGND VGND VPWR VPWR pp_row70_15 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_101_3 pp_row101_9 pp_row101_10 pp_row101_11 VGND VGND VPWR VPWR c$1940
+ s$1941 sky130_fd_sc_hd__fa_1
XFILLER_63_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_124_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_124_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_17_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_578 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_115_1 s$3381 s$3383 s$3385 VGND VGND VPWR VPWR c$3858 s$3859 sky130_fd_sc_hd__fa_1
Xdadda_fa_5_108_0 c$3332 c$3334 c$3336 VGND VGND VPWR VPWR c$3828 s$3829 sky130_fd_sc_hd__fa_1
X_1719_ clknet_leaf_21_clk booth_b22_m24 VGND VGND VPWR VPWR pp_row46_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_105_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_80_4 pp_row80_12 pp_row80_13 pp_row80_14 VGND VGND VPWR VPWR c$896 s$897
+ sky130_fd_sc_hd__fa_1
XFILLER_132_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout501 net502 VGND VGND VPWR VPWR net501 sky130_fd_sc_hd__buf_4
XFILLER_99_860 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout512 net518 VGND VGND VPWR VPWR net512 sky130_fd_sc_hd__buf_4
Xfanout523 net526 VGND VGND VPWR VPWR net523 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_73_3 pp_row73_18 pp_row73_19 pp_row73_20 VGND VGND VPWR VPWR c$768 s$769
+ sky130_fd_sc_hd__fa_1
Xfanout534 sel_0$4547 VGND VGND VPWR VPWR net534 sky130_fd_sc_hd__buf_4
XFILLER_150_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout545 net546 VGND VGND VPWR VPWR net545 sky130_fd_sc_hd__buf_6
Xfanout556 net558 VGND VGND VPWR VPWR net556 sky130_fd_sc_hd__buf_6
Xdadda_fa_4_50_2 s$2241 s$2243 s$2245 VGND VGND VPWR VPWR c$2994 s$2995 sky130_fd_sc_hd__fa_1
Xdadda_fa_1_66_2 pp_row66_24 pp_row66_25 pp_row66_26 VGND VGND VPWR VPWR c$640 s$641
+ sky130_fd_sc_hd__fa_1
Xfanout567 net568 VGND VGND VPWR VPWR net567 sky130_fd_sc_hd__clkbuf_8
Xfanout578 net579 VGND VGND VPWR VPWR net578 sky130_fd_sc_hd__buf_4
XFILLER_150_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout589 net592 VGND VGND VPWR VPWR net589 sky130_fd_sc_hd__clkbuf_8
Xdadda_fa_4_43_1 c$2178 c$2180 s$2183 VGND VGND VPWR VPWR c$2950 s$2951 sky130_fd_sc_hd__fa_1
XFILLER_101_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_59_1 pp_row59_14 pp_row59_15 pp_row59_16 VGND VGND VPWR VPWR c$512 s$513
+ sky130_fd_sc_hd__fa_1
XU$$4487_1864 VGND VGND VPWR VPWR U$$4487_1864/HI net1864 sky130_fd_sc_hd__conb_1
Xdadda_fa_7_20_0 s$3479 c$3934 s$3937 VGND VGND VPWR VPWR c$4192 s$4193 sky130_fd_sc_hd__fa_1
XFILLER_6_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_36_0 s$1169 c$2118 c$2120 VGND VGND VPWR VPWR c$2906 s$2907 sky130_fd_sc_hd__fa_1
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_5_2__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_5_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_115_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_115_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_167_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_88_3 s$1787 s$1789 s$1791 VGND VGND VPWR VPWR c$2548 s$2549 sky130_fd_sc_hd__fa_1
XFILLER_68_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_786 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4503 t$6705 net1872 VGND VGND VPWR VPWR booth_b64_m56 sky130_fd_sc_hd__xor2_1
XU$$4514 net1544 sel_0$6647 net1536 net693 VGND VGND VPWR VPWR t$6711 sky130_fd_sc_hd__a22o_1
Xdadda_fa_0_61_1 pp_row61_3 pp_row61_4 pp_row61_5 VGND VGND VPWR VPWR c$52 s$53 sky130_fd_sc_hd__fa_1
XTAP_4140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$17 t$4415 net1573 VGND VGND VPWR VPWR booth_b0_m5 sky130_fd_sc_hd__xor2_1
XU$$3802 t$6347 net1307 VGND VGND VPWR VPWR booth_b54_m48 sky130_fd_sc_hd__xor2_1
XU$$3813 net1634 net473 net1624 net746 VGND VGND VPWR VPWR t$6353 sky130_fd_sc_hd__a22o_1
XU$$28 net1224 net446 net1216 net688 VGND VGND VPWR VPWR t$4421 sky130_fd_sc_hd__a22o_1
XTAP_4162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_54_0 pp_row54_0 pp_row54_1 pp_row54_2 VGND VGND VPWR VPWR c$4 s$5 sky130_fd_sc_hd__fa_1
XFILLER_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3824 t$6358 net1306 VGND VGND VPWR VPWR booth_b54_m59 sky130_fd_sc_hd__xor2_1
XTAP_4173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$39 t$4426 net1568 VGND VGND VPWR VPWR booth_b0_m16 sky130_fd_sc_hd__xor2_1
XU$$3835 net1302 VGND VGND VPWR VPWR notsign$6364 sky130_fd_sc_hd__inv_1
XTAP_4184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3846 net1129 net464 net1037 net737 VGND VGND VPWR VPWR t$6371 sky130_fd_sc_hd__a22o_1
XTAP_4195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3857 t$6376 net1291 VGND VGND VPWR VPWR booth_b56_m7 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$190 final_adder.$signal$1154 final_adder.$signal$1155 VGND VGND VPWR
+ VPWR final_adder.p_new$318 sky130_fd_sc_hd__and2_1
XU$$3868 net1208 net464 net1200 net737 VGND VGND VPWR VPWR t$6382 sky130_fd_sc_hd__a22o_1
XTAP_3472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3879 t$6387 net1291 VGND VGND VPWR VPWR booth_b56_m18 sky130_fd_sc_hd__xor2_1
XTAP_3483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_450 net1506 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_461 net1683 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_106_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_106_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_19 sel_0$5247 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0952_ clknet_leaf_114_clk booth_b52_m46 VGND VGND VPWR VPWR pp_row98_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_14_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0883_ clknet_leaf_110_clk booth_b34_m61 VGND VGND VPWR VPWR pp_row95_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_158_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_90_3 pp_row90_20 pp_row90_21 c$1010 VGND VGND VPWR VPWR c$1812 s$1813
+ sky130_fd_sc_hd__fa_1
XFILLER_127_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_83_2 c$926 c$928 c$930 VGND VGND VPWR VPWR c$1726 s$1727 sky130_fd_sc_hd__fa_1
X_1504_ clknet_leaf_20_clk booth_b4_m34 VGND VGND VPWR VPWR pp_row38_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_141_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2484_ clknet_leaf_146_clk booth_b10_m59 VGND VGND VPWR VPWR pp_row69_3 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_60_1 s$3051 s$3053 s$3055 VGND VGND VPWR VPWR c$3638 s$3639 sky130_fd_sc_hd__fa_2
XFILLER_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_76_1 c$802 c$804 c$806 VGND VGND VPWR VPWR c$1640 s$1641 sky130_fd_sc_hd__fa_1
X_1435_ clknet_leaf_244_clk net184 VGND VGND VPWR VPWR pp_row34_19 sky130_fd_sc_hd__dfxtp_2
XFILLER_114_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_53_0 c$3002 c$3004 c$3006 VGND VGND VPWR VPWR c$3608 s$3609 sky130_fd_sc_hd__fa_1
Xdadda_fa_2_69_0 s$153 c$672 c$674 VGND VGND VPWR VPWR c$1554 s$1555 sky130_fd_sc_hd__fa_1
X_1366_ clknet_leaf_3_clk booth_b24_m7 VGND VGND VPWR VPWR pp_row31_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_56_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0317_ clknet_leaf_196_clk booth_b12_m62 VGND VGND VPWR VPWR pp_row74_2 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_52_8 pp_row52_26 pp_row52_27 pp_row52_28 VGND VGND VPWR VPWR c$400 s$401
+ sky130_fd_sc_hd__fa_2
X_1297_ clknet_leaf_251_clk booth_b0_m28 VGND VGND VPWR VPWR pp_row28_0 sky130_fd_sc_hd__dfxtp_1
X_0248_ clknet_leaf_197_clk net225 VGND VGND VPWR VPWR pp_row71_30 sky130_fd_sc_hd__dfxtp_2
XFILLER_110_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0179_ clknet_leaf_141_clk booth_b64_m5 VGND VGND VPWR VPWR pp_row69_30 sky130_fd_sc_hd__dfxtp_1
XFILLER_169_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_98_2 s$2625 s$2627 s$2629 VGND VGND VPWR VPWR c$3282 s$3283 sky130_fd_sc_hd__fa_1
XFILLER_152_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_68_0 s$3671 c$4030 s$4033 VGND VGND VPWR VPWR c$4288 s$4289 sky130_fd_sc_hd__fa_1
XFILLER_79_808 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1307 net1308 VGND VGND VPWR VPWR net1307 sky130_fd_sc_hd__buf_6
XFILLER_121_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1318 net5 VGND VGND VPWR VPWR net1318 sky130_fd_sc_hd__buf_8
Xdadda_fa_1_71_0 pp_row71_12 pp_row71_13 pp_row71_14 VGND VGND VPWR VPWR c$726 s$727
+ sky130_fd_sc_hd__fa_1
XFILLER_132_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1329 net1332 VGND VGND VPWR VPWR net1329 sky130_fd_sc_hd__buf_6
XFILLER_87_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout386 net392 VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__buf_4
XFILLER_86_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout397 net398 VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__buf_4
XU$$3109 t$5993 net1360 VGND VGND VPWR VPWR booth_b44_m44 sky130_fd_sc_hd__xor2_1
XFILLER_98_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2408 t$5635 net1425 VGND VGND VPWR VPWR booth_b34_m36 sky130_fd_sc_hd__xor2_1
XFILLER_28_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2419 net1747 net565 net1739 net838 VGND VGND VPWR VPWR t$5641 sky130_fd_sc_hd__a22o_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1707 t$5277 net1469 VGND VGND VPWR VPWR booth_b24_m28 sky130_fd_sc_hd__xor2_1
XFILLER_36_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1718 net996 net609 net988 net882 VGND VGND VPWR VPWR t$5283 sky130_fd_sc_hd__a22o_1
XFILLER_42_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1729 t$5288 net1473 VGND VGND VPWR VPWR booth_b24_m39 sky130_fd_sc_hd__xor2_1
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput17 a[24] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_2
XFILLER_168_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput28 a[34] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput39 a[44] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_93_1 c$1834 c$1836 c$1838 VGND VGND VPWR VPWR c$2584 s$2585 sky130_fd_sc_hd__fa_1
XFILLER_7_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_70_0 c$3672 c$3674 s$3677 VGND VGND VPWR VPWR c$4036 s$4037 sky130_fd_sc_hd__fa_1
XFILLER_182_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_86_0 s$989 c$1746 c$1748 VGND VGND VPWR VPWR c$2526 s$2527 sky130_fd_sc_hd__fa_1
XFILLER_170_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1220_ clknet_leaf_48_clk booth_b8_m15 VGND VGND VPWR VPWR pp_row23_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_81_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4300 t$6602 net1255 VGND VGND VPWR VPWR booth_b62_m23 sky130_fd_sc_hd__xor2_1
XFILLER_120_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4311 net1053 net422 net1045 net704 VGND VGND VPWR VPWR t$6608 sky130_fd_sc_hd__a22o_1
XU$$4322 t$6613 net1262 VGND VGND VPWR VPWR booth_b62_m34 sky130_fd_sc_hd__xor2_1
XU$$4333 net945 net424 net929 net706 VGND VGND VPWR VPWR t$6619 sky130_fd_sc_hd__a22o_1
XFILLER_38_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1151_ clknet_leaf_15_clk booth_b8_m10 VGND VGND VPWR VPWR pp_row18_4 sky130_fd_sc_hd__dfxtp_1
XU$$4344 t$6624 net1260 VGND VGND VPWR VPWR booth_b62_m45 sky130_fd_sc_hd__xor2_1
XU$$3610 net1120 net476 net1111 net749 VGND VGND VPWR VPWR t$6250 sky130_fd_sc_hd__a22o_1
XU$$4355 net1659 net423 net1651 net705 VGND VGND VPWR VPWR t$6630 sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_48_5 s$325 s$327 s$329 VGND VGND VPWR VPWR c$1312 s$1313 sky130_fd_sc_hd__fa_1
XU$$3621 t$6255 net1319 VGND VGND VPWR VPWR booth_b52_m26 sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_115_0 pp_row115_3 pp_row115_4 pp_row115_5 VGND VGND VPWR VPWR c$3380 s$3381
+ sky130_fd_sc_hd__fa_2
XFILLER_65_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4366 t$6635 net1260 VGND VGND VPWR VPWR booth_b62_m56 sky130_fd_sc_hd__xor2_1
XU$$3632 net1020 net477 net1003 net750 VGND VGND VPWR VPWR t$6261 sky130_fd_sc_hd__a22o_1
XU$$4377 net1545 net420 net1537 net702 VGND VGND VPWR VPWR t$6641 sky130_fd_sc_hd__a22o_1
X_1082_ clknet_leaf_248_clk net151 VGND VGND VPWR VPWR pp_row11_6 sky130_fd_sc_hd__dfxtp_2
XU$$3643 t$6266 net1322 VGND VGND VPWR VPWR booth_b52_m37 sky130_fd_sc_hd__xor2_1
XU$$4388 notblock$6645\[2\] net1813 net1260 t$6646 notblock$6645\[0\] VGND VGND VPWR
+ VPWR sel_0$6647 sky130_fd_sc_hd__a32o_1
XU$$4399 t$6653 net1820 VGND VGND VPWR VPWR booth_b64_m4 sky130_fd_sc_hd__xor2_1
XU$$3654 net1741 net480 net1733 net753 VGND VGND VPWR VPWR t$6272 sky130_fd_sc_hd__a22o_1
XFILLER_19_974 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3665 t$6277 net1326 VGND VGND VPWR VPWR booth_b52_m48 sky130_fd_sc_hd__xor2_1
XU$$2920 t$5897 net1367 VGND VGND VPWR VPWR booth_b42_m18 sky130_fd_sc_hd__xor2_1
XU$$2931 net1096 net526 net1087 net799 VGND VGND VPWR VPWR t$5903 sky130_fd_sc_hd__a22o_1
XFILLER_34_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3676 net1634 net483 net1624 net756 VGND VGND VPWR VPWR t$6283 sky130_fd_sc_hd__a22o_1
XTAP_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2942 t$5908 net1368 VGND VGND VPWR VPWR booth_b42_m29 sky130_fd_sc_hd__xor2_1
XU$$3687 t$6288 net1327 VGND VGND VPWR VPWR booth_b52_m59 sky130_fd_sc_hd__xor2_1
XTAP_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2953 net985 net520 net976 net793 VGND VGND VPWR VPWR t$5914 sky130_fd_sc_hd__a22o_1
XU$$3698 net1322 VGND VGND VPWR VPWR notsign$6294 sky130_fd_sc_hd__inv_1
XU$$2964 t$5919 net1370 VGND VGND VPWR VPWR booth_b42_m40 sky130_fd_sc_hd__xor2_1
XU$$2975 net1719 net522 net1710 net795 VGND VGND VPWR VPWR t$5925 sky130_fd_sc_hd__a22o_1
XU$$2986 t$5930 net1373 VGND VGND VPWR VPWR booth_b42_m51 sky130_fd_sc_hd__xor2_1
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2997 net1609 net525 net1602 net798 VGND VGND VPWR VPWR t$5936 sky130_fd_sc_hd__a22o_1
XANTENNA_280 c$580 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_291 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1984_ clknet_leaf_79_clk booth_b6_m49 VGND VGND VPWR VPWR pp_row55_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0935_ clknet_leaf_104_clk booth_b56_m41 VGND VGND VPWR VPWR pp_row97_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0866_ clknet_leaf_134_clk booth_b56_m64 VGND VGND VPWR VPWR pp_row120_1 sky130_fd_sc_hd__dfxtp_1
X_0797_ clknet_leaf_139_clk booth_b36_m55 VGND VGND VPWR VPWR pp_row91_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2467_ clknet_leaf_95_clk booth_b44_m24 VGND VGND VPWR VPWR pp_row68_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_69_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1418_ clknet_leaf_56_clk booth_b6_m28 VGND VGND VPWR VPWR pp_row34_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_69_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2398_ clknet_leaf_74_clk booth_b50_m16 VGND VGND VPWR VPWR pp_row66_25 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$904 final_adder.$signal$1204 final_adder.g_new$977 final_adder.$signal$230
+ VGND VGND VPWR VPWR final_adder.g_new$1032 sky130_fd_sc_hd__a21o_1
XFILLER_84_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$915 final_adder.$signal$1182 final_adder.g_new$999 final_adder.$signal$186
+ VGND VGND VPWR VPWR final_adder.g_new$1043 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$926 final_adder.$signal$1160 final_adder.g_new$1021 final_adder.$signal$142
+ VGND VGND VPWR VPWR final_adder.g_new$1054 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$937 final_adder.$signal$1138 final_adder.g_new$947 final_adder.$signal$98
+ VGND VGND VPWR VPWR final_adder.g_new$1065 sky130_fd_sc_hd__a21o_1
XFILLER_96_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1349_ clknet_leaf_123_clk booth_b42_m62 VGND VGND VPWR VPWR pp_row104_2 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_50_5 pp_row50_15 pp_row50_16 pp_row50_17 VGND VGND VPWR VPWR c$358 s$359
+ sky130_fd_sc_hd__fa_1
XFILLER_113_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$948 final_adder.$signal$1116 final_adder.g_new$857 final_adder.$signal$54
+ VGND VGND VPWR VPWR final_adder.g_new$1076 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$959 final_adder.$signal$1094 final_adder.g_new$509 final_adder.$signal$10
+ VGND VGND VPWR VPWR final_adder.g_new$1087 sky130_fd_sc_hd__a21o_1
XU$$809 net1590 net407 net1582 net673 VGND VGND VPWR VPWR t$4818 sky130_fd_sc_hd__a22o_1
XFILLER_84_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_1008 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1104 net79 VGND VGND VPWR VPWR net1104 sky130_fd_sc_hd__buf_4
XFILLER_191_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1115 net1116 VGND VGND VPWR VPWR net1115 sky130_fd_sc_hd__buf_2
XFILLER_105_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_746 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1126 net1128 VGND VGND VPWR VPWR net1126 sky130_fd_sc_hd__buf_4
XFILLER_120_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1137 net75 VGND VGND VPWR VPWR net1137 sky130_fd_sc_hd__clkbuf_8
Xfanout1148 net1154 VGND VGND VPWR VPWR net1148 sky130_fd_sc_hd__clkbuf_4
Xfanout1159 net72 VGND VGND VPWR VPWR net1159 sky130_fd_sc_hd__buf_6
XFILLER_47_524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2205 t$5532 net1432 VGND VGND VPWR VPWR booth_b32_m3 sky130_fd_sc_hd__xor2_1
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2216 net1503 net569 net1495 net842 VGND VGND VPWR VPWR t$5538 sky130_fd_sc_hd__a22o_1
XFILLER_170_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2227 t$5543 net1430 VGND VGND VPWR VPWR booth_b32_m14 sky130_fd_sc_hd__xor2_1
XU$$2238 net1133 net571 net1117 net844 VGND VGND VPWR VPWR t$5549 sky130_fd_sc_hd__a22o_1
XU$$1504 net1528 net633 net1762 net906 VGND VGND VPWR VPWR t$5173 sky130_fd_sc_hd__a22o_1
XU$$2249 t$5554 net1432 VGND VGND VPWR VPWR booth_b32_m25 sky130_fd_sc_hd__xor2_1
XU$$1515 net1230 net613 net1126 net886 VGND VGND VPWR VPWR t$5180 sky130_fd_sc_hd__a22o_1
XU$$1526 t$5185 net1475 VGND VGND VPWR VPWR booth_b22_m6 sky130_fd_sc_hd__xor2_1
XFILLER_43_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1537 net1216 net613 net1206 net886 VGND VGND VPWR VPWR t$5191 sky130_fd_sc_hd__a22o_1
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1548 t$5196 net1476 VGND VGND VPWR VPWR booth_b22_m17 sky130_fd_sc_hd__xor2_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1559 net1099 net611 net1089 net884 VGND VGND VPWR VPWR t$5202 sky130_fd_sc_hd__a22o_1
XFILLER_187_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0720_ clknet_leaf_161_clk booth_b26_m62 VGND VGND VPWR VPWR pp_row88_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_7_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0651_ clknet_leaf_168_clk booth_b36_m49 VGND VGND VPWR VPWR pp_row85_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_171_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0582_ clknet_leaf_173_clk booth_b58_m24 VGND VGND VPWR VPWR pp_row82_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_98_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2321_ clknet_leaf_77_clk booth_b44_m20 VGND VGND VPWR VPWR pp_row64_22 sky130_fd_sc_hd__dfxtp_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_2_60_4 s$533 s$535 s$537 VGND VGND VPWR VPWR c$1454 s$1455 sky130_fd_sc_hd__fa_2
X_2252_ clknet_leaf_149_clk booth_b54_m8 VGND VGND VPWR VPWR pp_row62_27 sky130_fd_sc_hd__dfxtp_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1660 net1661 VGND VGND VPWR VPWR net1660 sky130_fd_sc_hd__buf_4
XFILLER_84_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1203_ clknet_leaf_51_clk booth_b6_m16 VGND VGND VPWR VPWR pp_row22_3 sky130_fd_sc_hd__dfxtp_1
Xfanout1671 net1673 VGND VGND VPWR VPWR net1671 sky130_fd_sc_hd__buf_4
XFILLER_66_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_53_3 c$400 s$403 s$405 VGND VGND VPWR VPWR c$1368 s$1369 sky130_fd_sc_hd__fa_1
X_2183_ clknet_leaf_136_clk booth_b64_m45 VGND VGND VPWR VPWR pp_row109_10 sky130_fd_sc_hd__dfxtp_1
XU$$4130 net1525 net438 net1517 net720 VGND VGND VPWR VPWR t$6516 sky130_fd_sc_hd__a22o_1
Xfanout1682 net1683 VGND VGND VPWR VPWR net1682 sky130_fd_sc_hd__buf_4
Xfanout1693 net1694 VGND VGND VPWR VPWR net1693 sky130_fd_sc_hd__buf_4
XU$$4141 t$6521 net1263 VGND VGND VPWR VPWR booth_b60_m12 sky130_fd_sc_hd__xor2_1
XU$$4152 net1152 net434 net1142 net716 VGND VGND VPWR VPWR t$6527 sky130_fd_sc_hd__a22o_1
X_1134_ clknet_leaf_247_clk net164 VGND VGND VPWR VPWR pp_row16_10 sky130_fd_sc_hd__dfxtp_1
XU$$4163 t$6532 net1268 VGND VGND VPWR VPWR booth_b60_m23 sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_46_2 c$276 c$278 c$280 VGND VGND VPWR VPWR c$1282 s$1283 sky130_fd_sc_hd__fa_1
XFILLER_53_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_888 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4174 net1053 net437 net1045 net719 VGND VGND VPWR VPWR t$6538 sky130_fd_sc_hd__a22o_1
XU$$3440 t$6163 net1333 VGND VGND VPWR VPWR booth_b50_m4 sky130_fd_sc_hd__xor2_1
XFILLER_168_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_23_1 s$2829 s$2831 s$2833 VGND VGND VPWR VPWR c$3490 s$3491 sky130_fd_sc_hd__fa_1
XU$$4185 t$6543 net1272 VGND VGND VPWR VPWR booth_b60_m34 sky130_fd_sc_hd__xor2_1
XU$$4196 net945 net440 net929 net722 VGND VGND VPWR VPWR t$6549 sky130_fd_sc_hd__a22o_1
XU$$3451 net1498 net484 net1222 net757 VGND VGND VPWR VPWR t$6169 sky130_fd_sc_hd__a22o_1
XFILLER_25_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_39_1 pp_row39_11 pp_row39_12 pp_row39_13 VGND VGND VPWR VPWR c$1196 s$1197
+ sky130_fd_sc_hd__fa_1
XU$$3462 t$6174 net1333 VGND VGND VPWR VPWR booth_b50_m15 sky130_fd_sc_hd__xor2_1
XU$$3473 net1120 net487 net1111 net760 VGND VGND VPWR VPWR t$6180 sky130_fd_sc_hd__a22o_1
X_1065_ clknet_leaf_59_clk booth_b8_m1 VGND VGND VPWR VPWR pp_row9_4 sky130_fd_sc_hd__dfxtp_1
XU$$3484 t$6185 net1329 VGND VGND VPWR VPWR booth_b50_m26 sky130_fd_sc_hd__xor2_1
XFILLER_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2750 net1122 net535 net1031 net808 VGND VGND VPWR VPWR t$5811 sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_16_0 c$2780 c$2782 c$2784 VGND VGND VPWR VPWR c$3460 s$3461 sky130_fd_sc_hd__fa_1
XU$$3495 net1019 net485 net1002 net758 VGND VGND VPWR VPWR t$6191 sky130_fd_sc_hd__a22o_1
XU$$2761 t$5816 net1376 VGND VGND VPWR VPWR booth_b40_m7 sky130_fd_sc_hd__xor2_1
XU$$2772 net1207 net539 net1199 net812 VGND VGND VPWR VPWR t$5822 sky130_fd_sc_hd__a22o_1
XU$$2783 t$5827 net1377 VGND VGND VPWR VPWR booth_b40_m18 sky130_fd_sc_hd__xor2_1
XU$$2794 net1092 net539 net1084 net812 VGND VGND VPWR VPWR t$5833 sky130_fd_sc_hd__a22o_1
XFILLER_22_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1967_ clknet_leaf_63_clk booth_b36_m18 VGND VGND VPWR VPWR pp_row54_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0918_ clknet_leaf_104_clk booth_b62_m34 VGND VGND VPWR VPWR pp_row96_16 sky130_fd_sc_hd__dfxtp_1
X_1898_ clknet_leaf_64_clk booth_b26_m26 VGND VGND VPWR VPWR pp_row52_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_147_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0849_ clknet_leaf_109_clk booth_b48_m45 VGND VGND VPWR VPWR pp_row93_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_146_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput207 c[55] VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__clkbuf_1
Xinput218 c[65] VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__clkbuf_1
Xinput229 c[75] VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$701 final_adder.p_new$708 final_adder.g_new$725 final_adder.g_new$709
+ VGND VGND VPWR VPWR final_adder.g_new$829 sky130_fd_sc_hd__a21o_1
XFILLER_57_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$712 final_adder.p_new$736 final_adder.p_new$720 VGND VGND VPWR VPWR
+ final_adder.p_new$840 sky130_fd_sc_hd__and2_1
XFILLER_99_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$723 final_adder.p_new$730 final_adder.g_new$747 final_adder.g_new$731
+ VGND VGND VPWR VPWR final_adder.g_new$851 sky130_fd_sc_hd__a21o_2
Xclkbuf_leaf_95_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_95_clk sky130_fd_sc_hd__clkbuf_16
Xfinal_adder.U$$745 final_adder.p_new$760 final_adder.g_new$793 final_adder.g_new$761
+ VGND VGND VPWR VPWR final_adder.g_new$873 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$756 final_adder.p_new$804 final_adder.p_new$772 VGND VGND VPWR VPWR
+ final_adder.p_new$884 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$767 final_adder.p_new$782 final_adder.g_new$815 final_adder.g_new$783
+ VGND VGND VPWR VPWR final_adder.g_new$895 sky130_fd_sc_hd__a21o_1
XU$$606 net1075 net413 net1067 net679 VGND VGND VPWR VPWR t$4715 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$778 final_adder.p_new$826 final_adder.p_new$794 VGND VGND VPWR VPWR
+ final_adder.p_new$906 sky130_fd_sc_hd__and2_1
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$617 t$4720 net1241 VGND VGND VPWR VPWR booth_b8_m31 sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_41_1 pp_row41_3 pp_row41_4 pp_row41_5 VGND VGND VPWR VPWR c$238 s$239
+ sky130_fd_sc_hd__fa_1
XU$$628 net968 net415 net960 net681 VGND VGND VPWR VPWR t$4726 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$789 final_adder.p_new$804 final_adder.g_new$837 final_adder.g_new$805
+ VGND VGND VPWR VPWR final_adder.g_new$917 sky130_fd_sc_hd__a21o_1
XU$$639 t$4731 net1237 VGND VGND VPWR VPWR booth_b8_m42 sky130_fd_sc_hd__xor2_1
XFILLER_44_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_941 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_70_3 s$1571 s$1573 s$1575 VGND VGND VPWR VPWR c$2404 s$2405 sky130_fd_sc_hd__fa_1
XFILLER_140_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_63_2 c$1480 s$1483 s$1485 VGND VGND VPWR VPWR c$2346 s$2347 sky130_fd_sc_hd__fa_1
XFILLER_94_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_56_1 c$1390 c$1392 c$1394 VGND VGND VPWR VPWR c$2288 s$2289 sky130_fd_sc_hd__fa_1
XFILLER_48_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_33_0 c$3524 c$3526 s$3529 VGND VGND VPWR VPWR c$3962 s$3963 sky130_fd_sc_hd__fa_2
XFILLER_59_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_86_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_86_clk sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_3_49_0 s$347 c$1302 c$1304 VGND VGND VPWR VPWR c$2230 s$2231 sky130_fd_sc_hd__fa_2
XU$$2002 net954 net591 net946 net864 VGND VGND VPWR VPWR t$5428 sky130_fd_sc_hd__a22o_1
XU$$2013 t$5433 net1454 VGND VGND VPWR VPWR booth_b28_m44 sky130_fd_sc_hd__xor2_1
XFILLER_74_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2024 net1680 net590 net1655 net863 VGND VGND VPWR VPWR t$5439 sky130_fd_sc_hd__a22o_1
XFILLER_74_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2035 t$5444 net1454 VGND VGND VPWR VPWR booth_b28_m55 sky130_fd_sc_hd__xor2_1
XU$$1301 net1024 net636 net1015 net909 VGND VGND VPWR VPWR t$5070 sky130_fd_sc_hd__a22o_1
XU$$2046 net1556 net591 net1548 net864 VGND VGND VPWR VPWR t$5450 sky130_fd_sc_hd__a22o_1
XU$$1312 t$5075 net1666 VGND VGND VPWR VPWR booth_b18_m36 sky130_fd_sc_hd__xor2_1
XU$$2057 net1444 VGND VGND VPWR VPWR notblock$5455\[2\] sky130_fd_sc_hd__inv_1
XU$$1323 net1746 net640 net1738 net913 VGND VGND VPWR VPWR t$5081 sky130_fd_sc_hd__a22o_1
XU$$2068 t$5462 net1441 VGND VGND VPWR VPWR booth_b30_m3 sky130_fd_sc_hd__xor2_1
XU$$2079 net1505 net577 net1496 net850 VGND VGND VPWR VPWR t$5468 sky130_fd_sc_hd__a22o_1
XU$$1334 t$5086 net1670 VGND VGND VPWR VPWR booth_b18_m47 sky130_fd_sc_hd__xor2_1
XU$$1345 net1638 net640 net1629 net913 VGND VGND VPWR VPWR t$5092 sky130_fd_sc_hd__a22o_1
XU$$1356 t$5097 net1669 VGND VGND VPWR VPWR booth_b18_m58 sky130_fd_sc_hd__xor2_1
XU$$1367 net1528 net641 net1759 net914 VGND VGND VPWR VPWR t$5103 sky130_fd_sc_hd__a22o_1
Xdadda_ha_3_114_1 pp_row114_3 pp_row114_4 VGND VGND VPWR VPWR c$2744 s$2745 sky130_fd_sc_hd__ha_1
XU$$1378 net1230 net630 net1126 net903 VGND VGND VPWR VPWR t$5110 sky130_fd_sc_hd__a22o_1
XFILLER_30_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1389 t$5115 net1485 VGND VGND VPWR VPWR booth_b20_m6 sky130_fd_sc_hd__xor2_1
XFILLER_188_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1821_ clknet_leaf_235_clk net200 VGND VGND VPWR VPWR pp_row49_25 sky130_fd_sc_hd__dfxtp_1
XFILLER_175_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_106_0 s$3823 c$4106 s$4109 VGND VGND VPWR VPWR c$4364 s$4365 sky130_fd_sc_hd__fa_1
X_1752_ clknet_leaf_234_clk booth_b28_m19 VGND VGND VPWR VPWR pp_row47_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_10_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_156_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0703_ clknet_leaf_174_clk booth_b38_m49 VGND VGND VPWR VPWR pp_row87_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_183_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1683_ clknet_leaf_123_clk booth_b48_m58 VGND VGND VPWR VPWR pp_row106_4 sky130_fd_sc_hd__dfxtp_1
X_0634_ clknet_leaf_178_clk booth_b52_m32 VGND VGND VPWR VPWR pp_row84_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_171_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout908 net909 VGND VGND VPWR VPWR net908 sky130_fd_sc_hd__buf_4
X_0565_ clknet_leaf_188_clk booth_b28_m54 VGND VGND VPWR VPWR pp_row82_6 sky130_fd_sc_hd__dfxtp_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout919 net920 VGND VGND VPWR VPWR net919 sky130_fd_sc_hd__buf_6
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2304_ clknet_leaf_91_clk booth_b14_m50 VGND VGND VPWR VPWR pp_row64_7 sky130_fd_sc_hd__dfxtp_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0496_ clknet_leaf_158_clk booth_b58_m21 VGND VGND VPWR VPWR pp_row79_22 sky130_fd_sc_hd__dfxtp_1
XFILLER_98_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2235_ clknet_leaf_228_clk booth_b24_m38 VGND VGND VPWR VPWR pp_row62_12 sky130_fd_sc_hd__dfxtp_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_77_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_77_clk sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_2_51_0 pp_row51_26 c$348 c$350 VGND VGND VPWR VPWR c$1338 s$1339 sky130_fd_sc_hd__fa_2
XFILLER_38_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1490 net14 VGND VGND VPWR VPWR net1490 sky130_fd_sc_hd__buf_4
X_2166_ clknet_leaf_28_clk booth_b30_m30 VGND VGND VPWR VPWR pp_row60_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1117_ clknet_leaf_47_clk booth_b6_m9 VGND VGND VPWR VPWR pp_row15_3 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$30 c$4210 s$4213 VGND VGND VPWR VPWR final_adder.$signal$62 final_adder.$signal$1120
+ sky130_fd_sc_hd__ha_1
XFILLER_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2097_ clknet_leaf_86_clk booth_b30_m28 VGND VGND VPWR VPWR pp_row58_15 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$41 c$4232 s$4235 VGND VGND VPWR VPWR final_adder.$signal$84 final_adder.$signal$1131
+ sky130_fd_sc_hd__ha_2
XU$$3270 t$6075 net1356 VGND VGND VPWR VPWR booth_b46_m56 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$52 c$4254 s$4257 VGND VGND VPWR VPWR final_adder.$signal$106 final_adder.$signal$107
+ sky130_fd_sc_hd__ha_1
XFILLER_0_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3281 net1548 net508 net1540 net781 VGND VGND VPWR VPWR t$6081 sky130_fd_sc_hd__a22o_1
XU$$3292 notblock$6085\[2\] net43 net1352 t$6086 notblock$6085\[0\] VGND VGND VPWR
+ VPWR sel_0$6087 sky130_fd_sc_hd__a32o_2
Xfinal_adder.U$$63 c$4276 s$4279 VGND VGND VPWR VPWR final_adder.$signal$128 final_adder.$signal$1153
+ sky130_fd_sc_hd__ha_1
X_1048_ clknet_leaf_57_clk booth_b4_m3 VGND VGND VPWR VPWR pp_row7_2 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$74 c$4298 s$4301 VGND VGND VPWR VPWR final_adder.$signal$150 final_adder.$signal$1164
+ sky130_fd_sc_hd__ha_1
XFILLER_179_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$85 c$4320 s$4323 VGND VGND VPWR VPWR final_adder.$signal$172 final_adder.$signal$1175
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$96 c$4342 s$4345 VGND VGND VPWR VPWR final_adder.$signal$194 final_adder.$signal$1186
+ sky130_fd_sc_hd__ha_1
XFILLER_179_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2580 net1634 net557 net1624 net830 VGND VGND VPWR VPWR t$5723 sky130_fd_sc_hd__a22o_1
XU$$2591 t$5728 net1410 VGND VGND VPWR VPWR booth_b36_m59 sky130_fd_sc_hd__xor2_1
XFILLER_94_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1890 t$5370 net1465 VGND VGND VPWR VPWR booth_b26_m51 sky130_fd_sc_hd__xor2_1
XFILLER_10_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_80_2 s$2481 s$2483 s$2485 VGND VGND VPWR VPWR c$3174 s$3175 sky130_fd_sc_hd__fa_1
XFILLER_150_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_73_1 c$2418 c$2420 s$2423 VGND VGND VPWR VPWR c$3130 s$3131 sky130_fd_sc_hd__fa_1
XFILLER_162_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_89_1 pp_row89_3 pp_row89_4 pp_row89_5 VGND VGND VPWR VPWR c$1012 s$1013
+ sky130_fd_sc_hd__fa_1
XFILLER_122_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_50_0 s$3599 c$3994 s$3997 VGND VGND VPWR VPWR c$4252 s$4253 sky130_fd_sc_hd__fa_2
XU$$554_1882 VGND VGND VPWR VPWR U$$554_1882/HI net1882 sky130_fd_sc_hd__conb_1
Xdadda_fa_4_66_0 s$1529 c$2358 c$2360 VGND VGND VPWR VPWR c$3086 s$3087 sky130_fd_sc_hd__fa_1
XFILLER_48_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$520 final_adder.p_new$532 final_adder.p_new$524 VGND VGND VPWR VPWR
+ final_adder.p_new$648 sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_68_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_68_clk sky130_fd_sc_hd__clkbuf_16
XTAP_3802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$531 final_adder.p_new$534 final_adder.g_new$543 final_adder.g_new$535
+ VGND VGND VPWR VPWR final_adder.g_new$659 sky130_fd_sc_hd__a21o_1
XTAP_3813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$542 final_adder.p_new$554 final_adder.p_new$546 VGND VGND VPWR VPWR
+ final_adder.p_new$670 sky130_fd_sc_hd__and2_1
XTAP_3824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$553 final_adder.p_new$556 final_adder.g_new$565 final_adder.g_new$557
+ VGND VGND VPWR VPWR final_adder.g_new$681 sky130_fd_sc_hd__a21o_1
XFILLER_57_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$403 t$4610 net1280 VGND VGND VPWR VPWR booth_b4_m61 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$564 final_adder.p_new$576 final_adder.p_new$568 VGND VGND VPWR VPWR
+ final_adder.p_new$692 sky130_fd_sc_hd__and2_1
XTAP_3846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$414 net1246 notblock$4615\[1\] VGND VGND VPWR VPWR t$4616 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$575 final_adder.p_new$578 final_adder.g_new$587 final_adder.g_new$579
+ VGND VGND VPWR VPWR final_adder.g_new$703 sky130_fd_sc_hd__a21o_1
XFILLER_178_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$425 net936 net430 net1676 net712 VGND VGND VPWR VPWR t$4623 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$586 final_adder.p_new$598 final_adder.p_new$590 VGND VGND VPWR VPWR
+ final_adder.p_new$714 sky130_fd_sc_hd__and2_1
XTAP_3868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$436 t$4628 net1250 VGND VGND VPWR VPWR booth_b6_m9 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$597 final_adder.p_new$600 final_adder.g_new$609 final_adder.g_new$601
+ VGND VGND VPWR VPWR final_adder.g_new$725 sky130_fd_sc_hd__a21o_1
XTAP_3879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$447 net1180 net429 net1171 net711 VGND VGND VPWR VPWR t$4634 sky130_fd_sc_hd__a22o_1
XFILLER_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$458 t$4639 net1244 VGND VGND VPWR VPWR booth_b6_m20 sky130_fd_sc_hd__xor2_1
XU$$469 net1072 net427 net1064 net709 VGND VGND VPWR VPWR t$4645 sky130_fd_sc_hd__a22o_1
XFILLER_60_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1001 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0350_ clknet_leaf_200_clk booth_b14_m61 VGND VGND VPWR VPWR pp_row75_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_67_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0281_ clknet_leaf_196_clk booth_b64_m8 VGND VGND VPWR VPWR pp_row72_29 sky130_fd_sc_hd__dfxtp_1
XFILLER_48_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_59_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_59_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_76_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2020_ clknet_leaf_38_clk booth_b14_m42 VGND VGND VPWR VPWR pp_row56_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_47_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$970 t$4901 net1183 VGND VGND VPWR VPWR booth_b14_m2 sky130_fd_sc_hd__xor2_1
XU$$1120 net1505 net644 net1496 net917 VGND VGND VPWR VPWR t$4978 sky130_fd_sc_hd__a22o_1
XU$$981 net1513 net387 net1505 net653 VGND VGND VPWR VPWR t$4907 sky130_fd_sc_hd__a22o_1
XFILLER_189_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$992 t$4912 net1183 VGND VGND VPWR VPWR booth_b14_m13 sky130_fd_sc_hd__xor2_1
XU$$1131 t$4983 net1006 VGND VGND VPWR VPWR booth_b16_m14 sky130_fd_sc_hd__xor2_1
XU$$1142 net1133 net645 net1117 net918 VGND VGND VPWR VPWR t$4989 sky130_fd_sc_hd__a22o_1
XU$$1153 t$4994 net1007 VGND VGND VPWR VPWR booth_b16_m25 sky130_fd_sc_hd__xor2_1
XU$$1164 net1023 net644 net1015 net917 VGND VGND VPWR VPWR t$5000 sky130_fd_sc_hd__a22o_1
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1175 t$5005 net1010 VGND VGND VPWR VPWR booth_b16_m36 sky130_fd_sc_hd__xor2_1
XFILLER_149_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1186 net1749 net645 net1741 net918 VGND VGND VPWR VPWR t$5011 sky130_fd_sc_hd__a22o_1
XU$$1197 t$5016 net1008 VGND VGND VPWR VPWR booth_b16_m47 sky130_fd_sc_hd__xor2_1
XFILLER_191_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1804_ clknet_leaf_220_clk booth_b20_m29 VGND VGND VPWR VPWR pp_row49_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_163_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_90_1 s$3231 s$3233 s$3235 VGND VGND VPWR VPWR c$3758 s$3759 sky130_fd_sc_hd__fa_1
XFILLER_163_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1735_ clknet_leaf_235_clk net197 VGND VGND VPWR VPWR pp_row46_25 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_83_0 c$3182 c$3184 c$3186 VGND VGND VPWR VPWR c$3728 s$3729 sky130_fd_sc_hd__fa_1
XFILLER_116_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_99_0 pp_row99_0 pp_row99_1 pp_row99_2 VGND VGND VPWR VPWR c$1914 s$1915
+ sky130_fd_sc_hd__fa_1
XFILLER_176_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_1107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1666_ clknet_leaf_21_clk booth_b24_m20 VGND VGND VPWR VPWR pp_row44_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_104_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0617_ clknet_leaf_187_clk booth_b22_m62 VGND VGND VPWR VPWR pp_row84_2 sky130_fd_sc_hd__dfxtp_1
Xfanout705 net707 VGND VGND VPWR VPWR net705 sky130_fd_sc_hd__buf_4
X_1597_ clknet_leaf_5_clk booth_b38_m3 VGND VGND VPWR VPWR pp_row41_19 sky130_fd_sc_hd__dfxtp_1
Xfanout716 net719 VGND VGND VPWR VPWR net716 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_75_7 pp_row75_27 pp_row75_28 c$186 VGND VGND VPWR VPWR c$812 s$813 sky130_fd_sc_hd__fa_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout727 net732 VGND VGND VPWR VPWR net727 sky130_fd_sc_hd__buf_4
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout738 net740 VGND VGND VPWR VPWR net738 sky130_fd_sc_hd__clkbuf_8
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0548_ clknet_leaf_171_clk booth_b46_m35 VGND VGND VPWR VPWR pp_row81_15 sky130_fd_sc_hd__dfxtp_1
Xfanout749 net752 VGND VGND VPWR VPWR net749 sky130_fd_sc_hd__buf_6
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_68_6 c$124 c$126 c$128 VGND VGND VPWR VPWR c$684 s$685 sky130_fd_sc_hd__fa_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0479_ clknet_leaf_205_clk booth_b26_m53 VGND VGND VPWR VPWR pp_row79_6 sky130_fd_sc_hd__dfxtp_1
XTAP_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_972 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2218_ clknet_leaf_29_clk booth_b56_m5 VGND VGND VPWR VPWR pp_row61_28 sky130_fd_sc_hd__dfxtp_1
XFILLER_27_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_109 net615 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2149_ clknet_leaf_144_clk booth_b58_m51 VGND VGND VPWR VPWR pp_row109_7 sky130_fd_sc_hd__dfxtp_1
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_7_98_0 s$3791 c$4090 s$4093 VGND VGND VPWR VPWR c$4348 s$4349 sky130_fd_sc_hd__fa_1
XFILLER_155_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_885 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_113_0 c$3844 c$3846 s$3849 VGND VGND VPWR VPWR c$4122 s$4123 sky130_fd_sc_hd__fa_1
XTAP_4344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$350 final_adder.p_new$352 final_adder.p_new$350 VGND VGND VPWR VPWR
+ final_adder.p_new$478 sky130_fd_sc_hd__and2_1
XTAP_4377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$200 t$4507 net1385 VGND VGND VPWR VPWR booth_b2_m28 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$361 final_adder.p_new$360 final_adder.g_new$363 final_adder.g_new$361
+ VGND VGND VPWR VPWR final_adder.g_new$489 sky130_fd_sc_hd__a21o_1
XTAP_4388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$372 final_adder.p_new$374 final_adder.p_new$372 VGND VGND VPWR VPWR
+ final_adder.p_new$500 sky130_fd_sc_hd__and2_1
XU$$211 net992 net625 net987 net898 VGND VGND VPWR VPWR t$4513 sky130_fd_sc_hd__a22o_1
XTAP_4399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$222 t$4518 net1385 VGND VGND VPWR VPWR booth_b2_m39 sky130_fd_sc_hd__xor2_1
XFILLER_57_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_33_3 s$1127 s$1129 s$1131 VGND VGND VPWR VPWR c$2108 s$2109 sky130_fd_sc_hd__fa_1
XTAP_3665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$233 net1720 net621 net1711 net894 VGND VGND VPWR VPWR t$4524 sky130_fd_sc_hd__a22o_1
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$394 final_adder.p_new$400 final_adder.p_new$396 VGND VGND VPWR VPWR
+ final_adder.p_new$522 sky130_fd_sc_hd__and2_1
XFILLER_18_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$244 t$4529 net1392 VGND VGND VPWR VPWR booth_b2_m50 sky130_fd_sc_hd__xor2_1
XTAP_3687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$255 net1615 net626 net1607 net899 VGND VGND VPWR VPWR t$4535 sky130_fd_sc_hd__a22o_1
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$266 t$4540 net1387 VGND VGND VPWR VPWR booth_b2_m61 sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_26_2 pp_row26_14 pp_row26_15 c$1058 VGND VGND VPWR VPWR c$2050 s$2051
+ sky130_fd_sc_hd__fa_1
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$277 net1275 notblock$4545\[1\] VGND VGND VPWR VPWR t$4546 sky130_fd_sc_hd__and2_1
XTAP_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$288 net937 net531 net1675 net804 VGND VGND VPWR VPWR t$4553 sky130_fd_sc_hd__a22o_1
XTAP_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$299 t$4558 net1278 VGND VGND VPWR VPWR booth_b4_m9 sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_19_1 pp_row19_3 pp_row19_4 pp_row19_5 VGND VGND VPWR VPWR c$1994 s$1995
+ sky130_fd_sc_hd__fa_1
XTAP_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4505_1873 VGND VGND VPWR VPWR U$$4505_1873/HI net1873 sky130_fd_sc_hd__conb_1
XFILLER_40_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$5 net1 net1880 VGND VGND VPWR VPWR sel_1 sky130_fd_sc_hd__xor2_1
XFILLER_173_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput308 net308 VGND VGND VPWR VPWR o[30] sky130_fd_sc_hd__buf_2
XFILLER_154_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_903 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput319 net319 VGND VGND VPWR VPWR o[40] sky130_fd_sc_hd__buf_2
X_1520_ clknet_leaf_246_clk booth_b30_m8 VGND VGND VPWR VPWR pp_row38_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1451_ clknet_leaf_65_clk booth_b26_m9 VGND VGND VPWR VPWR pp_row35_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_45_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_78_5 s$863 s$865 s$867 VGND VGND VPWR VPWR c$1672 s$1673 sky130_fd_sc_hd__fa_1
X_0402_ clknet_leaf_208_clk booth_b50_m26 VGND VGND VPWR VPWR pp_row76_20 sky130_fd_sc_hd__dfxtp_1
X_1382_ clknet_leaf_110_clk booth_b48_m56 VGND VGND VPWR VPWR pp_row104_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_45_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_990 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0333_ clknet_leaf_128_clk booth_b50_m64 VGND VGND VPWR VPWR pp_row114_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_121_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0264_ clknet_leaf_150_clk booth_b36_m36 VGND VGND VPWR VPWR pp_row72_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_95_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2003_ clknet_leaf_73_clk booth_b42_m13 VGND VGND VPWR VPWR pp_row55_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_64_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0195_ clknet_leaf_155_clk booth_b32_m38 VGND VGND VPWR VPWR pp_row70_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_23_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_108_1 s$3339 s$3341 s$3343 VGND VGND VPWR VPWR c$3830 s$3831 sky130_fd_sc_hd__fa_1
X_1718_ clknet_leaf_21_clk booth_b20_m26 VGND VGND VPWR VPWR pp_row46_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_172_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1649_ clknet_leaf_239_clk booth_b40_m3 VGND VGND VPWR VPWR pp_row43_20 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_80_5 pp_row80_15 pp_row80_16 pp_row80_17 VGND VGND VPWR VPWR c$898 s$899
+ sky130_fd_sc_hd__fa_1
XFILLER_104_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout502 net509 VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__clkbuf_4
Xfanout513 net518 VGND VGND VPWR VPWR net513 sky130_fd_sc_hd__buf_4
XFILLER_116_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout524 net525 VGND VGND VPWR VPWR net524 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_73_4 pp_row73_21 pp_row73_22 pp_row73_23 VGND VGND VPWR VPWR c$770 s$771
+ sky130_fd_sc_hd__fa_1
XFILLER_113_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout535 net536 VGND VGND VPWR VPWR net535 sky130_fd_sc_hd__clkbuf_8
XFILLER_98_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout546 net550 VGND VGND VPWR VPWR net546 sky130_fd_sc_hd__buf_6
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout557 net558 VGND VGND VPWR VPWR net557 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_66_3 pp_row66_27 pp_row66_28 pp_row66_29 VGND VGND VPWR VPWR c$642 s$643
+ sky130_fd_sc_hd__fa_1
XFILLER_150_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout568 sel_0$5597 VGND VGND VPWR VPWR net568 sky130_fd_sc_hd__buf_8
XFILLER_58_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout579 net583 VGND VGND VPWR VPWR net579 sky130_fd_sc_hd__buf_6
XFILLER_112_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_43_2 s$2185 s$2187 s$2189 VGND VGND VPWR VPWR c$2952 s$2953 sky130_fd_sc_hd__fa_1
XFILLER_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_59_2 pp_row59_17 pp_row59_18 pp_row59_19 VGND VGND VPWR VPWR c$514 s$515
+ sky130_fd_sc_hd__fa_1
Xdadda_fa_4_36_1 c$2122 c$2124 s$2127 VGND VGND VPWR VPWR c$2908 s$2909 sky130_fd_sc_hd__fa_1
XFILLER_55_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_13_0 s$3451 c$3920 s$3923 VGND VGND VPWR VPWR c$4178 s$4179 sky130_fd_sc_hd__fa_1
Xdadda_fa_4_29_0 s$1089 c$2062 c$2064 VGND VGND VPWR VPWR c$2864 s$2865 sky130_fd_sc_hd__fa_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_798 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4504 net1605 sel_0$6647 net1597 net693 VGND VGND VPWR VPWR t$6706 sky130_fd_sc_hd__a22o_1
XFILLER_77_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4515 t$6711 net1878 VGND VGND VPWR VPWR booth_b64_m62 sky130_fd_sc_hd__xor2_1
Xdadda_fa_0_61_2 pp_row61_6 pp_row61_7 pp_row61_8 VGND VGND VPWR VPWR c$54 s$55 sky130_fd_sc_hd__fa_1
XTAP_4130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3803 net1693 net474 net1684 net747 VGND VGND VPWR VPWR t$6348 sky130_fd_sc_hd__a22o_1
XTAP_4152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$18 net1565 net447 net1524 net689 VGND VGND VPWR VPWR t$4416 sky130_fd_sc_hd__a22o_1
XU$$3814 t$6353 net1306 VGND VGND VPWR VPWR booth_b54_m54 sky130_fd_sc_hd__xor2_1
XTAP_4163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$29 t$4421 net1573 VGND VGND VPWR VPWR booth_b0_m11 sky130_fd_sc_hd__xor2_1
XTAP_4174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3825 net1583 net473 net1556 net746 VGND VGND VPWR VPWR t$6359 sky130_fd_sc_hd__a22o_1
XTAP_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3836 net1302 VGND VGND VPWR VPWR notblock$6365\[0\] sky130_fd_sc_hd__inv_1
XTAP_4185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_31_0 pp_row31_14 pp_row31_15 pp_row31_16 VGND VGND VPWR VPWR c$2086 s$2087
+ sky130_fd_sc_hd__fa_1
XU$$3847 t$6371 net1296 VGND VGND VPWR VPWR booth_b56_m2 sky130_fd_sc_hd__xor2_1
XFILLER_131_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3858 net1517 net467 net1510 net740 VGND VGND VPWR VPWR t$6377 sky130_fd_sc_hd__a22o_1
XTAP_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$180 final_adder.$signal$1164 final_adder.$signal$1165 VGND VGND VPWR
+ VPWR final_adder.p_new$308 sky130_fd_sc_hd__and2_1
XU$$3869 t$6382 net1299 VGND VGND VPWR VPWR booth_b56_m13 sky130_fd_sc_hd__xor2_1
XTAP_3462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$191 final_adder.$signal$1155 final_adder.$signal$130 final_adder.$signal$132
+ VGND VGND VPWR VPWR final_adder.g_new$319 sky130_fd_sc_hd__a21o_1
XTAP_3473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_440 net967 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_451 net1518 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_462 net1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0951_ clknet_leaf_114_clk booth_b50_m48 VGND VGND VPWR VPWR pp_row98_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0882_ clknet_leaf_110_clk booth_b32_m63 VGND VGND VPWR VPWR pp_row95_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_174_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_90_4 c$1012 c$1014 c$1016 VGND VGND VPWR VPWR c$1814 s$1815 sky130_fd_sc_hd__fa_2
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_83_3 c$932 c$934 c$936 VGND VGND VPWR VPWR c$1728 s$1729 sky130_fd_sc_hd__fa_1
X_1503_ clknet_leaf_17_clk booth_b2_m36 VGND VGND VPWR VPWR pp_row38_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_173_1137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2483_ clknet_leaf_147_clk booth_b8_m61 VGND VGND VPWR VPWR pp_row69_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_142_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_76_2 c$808 c$810 c$812 VGND VGND VPWR VPWR c$1642 s$1643 sky130_fd_sc_hd__fa_1
X_1434_ clknet_leaf_40_clk net1423 VGND VGND VPWR VPWR pp_row34_18 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_53_1 s$3009 s$3011 s$3013 VGND VGND VPWR VPWR c$3610 s$3611 sky130_fd_sc_hd__fa_1
XFILLER_68_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_69_1 c$676 c$678 c$680 VGND VGND VPWR VPWR c$1556 s$1557 sky130_fd_sc_hd__fa_2
XFILLER_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1365_ clknet_leaf_9_clk booth_b22_m9 VGND VGND VPWR VPWR pp_row31_11 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_46_0 c$2960 c$2962 c$2964 VGND VGND VPWR VPWR c$3580 s$3581 sky130_fd_sc_hd__fa_1
XFILLER_28_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0316_ clknet_leaf_196_clk booth_b10_m64 VGND VGND VPWR VPWR pp_row74_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1296_ clknet_leaf_248_clk net176 VGND VGND VPWR VPWR pp_row27_14 sky130_fd_sc_hd__dfxtp_1
X_0247_ clknet_leaf_146_clk booth_b64_m7 VGND VGND VPWR VPWR pp_row71_29 sky130_fd_sc_hd__dfxtp_1
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0178_ clknet_leaf_125_clk booth_b60_m52 VGND VGND VPWR VPWR pp_row112_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_120_0 pp_row120_5 pp_row120_6 c$3404 VGND VGND VPWR VPWR c$3876 s$3877
+ sky130_fd_sc_hd__fa_1
XFILLER_137_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1308 net1309 VGND VGND VPWR VPWR net1308 sky130_fd_sc_hd__buf_4
Xfanout1319 net1328 VGND VGND VPWR VPWR net1319 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_71_1 pp_row71_15 pp_row71_16 pp_row71_17 VGND VGND VPWR VPWR c$728 s$729
+ sky130_fd_sc_hd__fa_1
XFILLER_99_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_64_0 pp_row64_18 pp_row64_19 pp_row64_20 VGND VGND VPWR VPWR c$600 s$601
+ sky130_fd_sc_hd__fa_2
XFILLER_8_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout387 net389 VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__buf_4
XFILLER_115_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout398 net399 VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__clkbuf_4
XFILLER_189_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2409 net967 net565 net958 net838 VGND VGND VPWR VPWR t$5636 sky130_fd_sc_hd__a22o_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1708 net1049 net605 net1041 net878 VGND VGND VPWR VPWR t$5278 sky130_fd_sc_hd__a22o_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1719 t$5283 net1474 VGND VGND VPWR VPWR booth_b24_m34 sky130_fd_sc_hd__xor2_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$408_1803 VGND VGND VPWR VPWR U$$408_1803/HI net1803 sky130_fd_sc_hd__conb_1
XFILLER_188_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput18 a[25] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_6
XFILLER_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput29 a[35] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_128_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_93_2 c$1840 s$1843 s$1845 VGND VGND VPWR VPWR c$2586 s$2587 sky130_fd_sc_hd__fa_1
XFILLER_182_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_86_1 c$1750 c$1752 c$1754 VGND VGND VPWR VPWR c$2528 s$2529 sky130_fd_sc_hd__fa_1
XFILLER_124_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_63_0 c$3644 c$3646 s$3649 VGND VGND VPWR VPWR c$4022 s$4023 sky130_fd_sc_hd__fa_1
XFILLER_184_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_79_0 s$887 c$1662 c$1664 VGND VGND VPWR VPWR c$2470 s$2471 sky130_fd_sc_hd__fa_1
XFILLER_69_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_777 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_0_53_0 pp_row53_0 pp_row53_1 VGND VGND VPWR VPWR c$2 s$3 sky130_fd_sc_hd__ha_1
XFILLER_123_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4301 net1095 net420 net1085 net702 VGND VGND VPWR VPWR t$6603 sky130_fd_sc_hd__a22o_1
XFILLER_42_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4312 t$6608 net1259 VGND VGND VPWR VPWR booth_b62_m29 sky130_fd_sc_hd__xor2_1
XU$$4323 net989 net423 net980 net705 VGND VGND VPWR VPWR t$6614 sky130_fd_sc_hd__a22o_1
XFILLER_78_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1150_ clknet_leaf_14_clk booth_b6_m12 VGND VGND VPWR VPWR pp_row18_3 sky130_fd_sc_hd__dfxtp_1
XU$$4334 t$6619 net1261 VGND VGND VPWR VPWR booth_b62_m40 sky130_fd_sc_hd__xor2_1
XU$$3600 net1172 net481 net1163 net754 VGND VGND VPWR VPWR t$6245 sky130_fd_sc_hd__a22o_1
XU$$4345 net1719 net420 net1710 net702 VGND VGND VPWR VPWR t$6625 sky130_fd_sc_hd__a22o_1
XU$$3611 t$6250 net1319 VGND VGND VPWR VPWR booth_b52_m21 sky130_fd_sc_hd__xor2_1
XFILLER_93_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4356 t$6630 net1260 VGND VGND VPWR VPWR booth_b62_m51 sky130_fd_sc_hd__xor2_1
XU$$3622 net1068 net478 net1060 net751 VGND VGND VPWR VPWR t$6256 sky130_fd_sc_hd__a22o_1
XU$$4367 net1610 net423 net1601 net705 VGND VGND VPWR VPWR t$6636 sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_115_1 pp_row115_6 pp_row115_7 pp_row115_8 VGND VGND VPWR VPWR c$3382 s$3383
+ sky130_fd_sc_hd__fa_1
XU$$3633 t$6261 net1323 VGND VGND VPWR VPWR booth_b52_m32 sky130_fd_sc_hd__xor2_1
XFILLER_19_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1081_ clknet_leaf_53_clk booth_b10_m1 VGND VGND VPWR VPWR pp_row11_5 sky130_fd_sc_hd__dfxtp_1
XU$$4378 t$6641 net1257 VGND VGND VPWR VPWR booth_b62_m62 sky130_fd_sc_hd__xor2_1
XFILLER_34_901 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4389 net1814 net1256 VGND VGND VPWR VPWR sel_1$6648 sky130_fd_sc_hd__xor2_2
XU$$3644 net962 net483 net954 net756 VGND VGND VPWR VPWR t$6267 sky130_fd_sc_hd__a22o_1
XU$$2910 t$5892 net1372 VGND VGND VPWR VPWR booth_b42_m13 sky130_fd_sc_hd__xor2_1
XU$$3655 t$6272 net1325 VGND VGND VPWR VPWR booth_b52_m43 sky130_fd_sc_hd__xor2_1
XFILLER_19_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3666 net1694 net482 net1686 net755 VGND VGND VPWR VPWR t$6278 sky130_fd_sc_hd__a22o_1
XU$$2921 net1141 net520 net1136 net793 VGND VGND VPWR VPWR t$5898 sky130_fd_sc_hd__a22o_1
XFILLER_92_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_108_0 s$1973 c$2694 c$2696 VGND VGND VPWR VPWR c$3338 s$3339 sky130_fd_sc_hd__fa_1
XU$$2932 t$5903 net1372 VGND VGND VPWR VPWR booth_b42_m24 sky130_fd_sc_hd__xor2_1
XU$$3677 t$6283 net1327 VGND VGND VPWR VPWR booth_b52_m54 sky130_fd_sc_hd__xor2_1
XTAP_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2943 net1040 net519 net1024 net792 VGND VGND VPWR VPWR t$5909 sky130_fd_sc_hd__a22o_1
XU$$3688 net1583 net483 net1556 net756 VGND VGND VPWR VPWR t$6289 sky130_fd_sc_hd__a22o_1
XTAP_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2954 t$5914 net1368 VGND VGND VPWR VPWR booth_b42_m35 sky130_fd_sc_hd__xor2_1
XTAP_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3699 net1321 VGND VGND VPWR VPWR notblock$6295\[0\] sky130_fd_sc_hd__inv_1
XU$$2965 net926 net522 net1747 net795 VGND VGND VPWR VPWR t$5920 sky130_fd_sc_hd__a22o_1
XU$$2976 t$5925 net1371 VGND VGND VPWR VPWR booth_b42_m46 sky130_fd_sc_hd__xor2_1
XFILLER_179_939 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2987 net1652 net524 net1644 net797 VGND VGND VPWR VPWR t$5931 sky130_fd_sc_hd__a22o_1
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_270 net1741 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2998 t$5936 net1373 VGND VGND VPWR VPWR booth_b42_m57 sky130_fd_sc_hd__xor2_1
XANTENNA_281 final_adder.p_new$604 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_292 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1983_ clknet_leaf_136_clk booth_b52_m56 VGND VGND VPWR VPWR pp_row108_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_193_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0934_ clknet_leaf_112_clk booth_b54_m43 VGND VGND VPWR VPWR pp_row97_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0865_ clknet_leaf_111_clk booth_b40_m54 VGND VGND VPWR VPWR pp_row94_6 sky130_fd_sc_hd__dfxtp_1
X_0796_ clknet_leaf_140_clk booth_b34_m57 VGND VGND VPWR VPWR pp_row91_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_114_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_81_0 pp_row81_24 pp_row81_25 c$888 VGND VGND VPWR VPWR c$1698 s$1699 sky130_fd_sc_hd__fa_1
XFILLER_138_1043 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_1_51_8 pp_row51_24 pp_row51_25 VGND VGND VPWR VPWR c$382 s$383 sky130_fd_sc_hd__ha_1
X_2466_ clknet_leaf_95_clk booth_b42_m26 VGND VGND VPWR VPWR pp_row68_20 sky130_fd_sc_hd__dfxtp_1
XFILLER_142_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1417_ clknet_leaf_121_clk booth_b54_m50 VGND VGND VPWR VPWR pp_row104_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_60_1115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2397_ clknet_leaf_74_clk booth_b48_m18 VGND VGND VPWR VPWR pp_row66_24 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$905 final_adder.$signal$1202 final_adder.g_new$979 final_adder.$signal$226
+ VGND VGND VPWR VPWR final_adder.g_new$1033 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$916 final_adder.$signal$1180 final_adder.g_new$1001 final_adder.$signal$182
+ VGND VGND VPWR VPWR final_adder.g_new$1044 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$927 final_adder.$signal$1158 final_adder.g_new$1023 final_adder.$signal$138
+ VGND VGND VPWR VPWR final_adder.g_new$1055 sky130_fd_sc_hd__a21o_1
XFILLER_29_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1348_ clknet_leaf_241_clk booth_b28_m2 VGND VGND VPWR VPWR pp_row30_14 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$938 final_adder.$signal$1136 final_adder.g_new$949 final_adder.$signal$94
+ VGND VGND VPWR VPWR final_adder.g_new$1066 sky130_fd_sc_hd__a21o_1
Xdadda_fa_1_50_6 pp_row50_18 pp_row50_19 pp_row50_20 VGND VGND VPWR VPWR c$360 s$361
+ sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$949 final_adder.$signal$1114 final_adder.g_new$859 final_adder.$signal$50
+ VGND VGND VPWR VPWR final_adder.g_new$1077 sky130_fd_sc_hd__a21o_1
XFILLER_44_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1279_ clknet_leaf_251_clk booth_b0_m27 VGND VGND VPWR VPWR pp_row27_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_58_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_2_0 pp_row2_2 pp_row2_3 s$3901 VGND VGND VPWR VPWR c$4156 s$4157 sky130_fd_sc_hd__fa_1
XFILLER_58_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1025 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_80_0 s$3719 c$4054 s$4057 VGND VGND VPWR VPWR c$4312 s$4313 sky130_fd_sc_hd__fa_2
XFILLER_193_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_96_0 s$1889 c$2598 c$2600 VGND VGND VPWR VPWR c$3266 s$3267 sky130_fd_sc_hd__fa_1
XFILLER_4_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1105 net1110 VGND VGND VPWR VPWR net1105 sky130_fd_sc_hd__buf_4
Xfanout1116 net77 VGND VGND VPWR VPWR net1116 sky130_fd_sc_hd__buf_6
XFILLER_121_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1127 net1128 VGND VGND VPWR VPWR net1127 sky130_fd_sc_hd__clkbuf_4
Xfanout1138 net1140 VGND VGND VPWR VPWR net1138 sky130_fd_sc_hd__buf_4
XFILLER_121_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1149 net1154 VGND VGND VPWR VPWR net1149 sky130_fd_sc_hd__clkbuf_8
XFILLER_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_878 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_1081 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2206 net936 net571 net1676 net844 VGND VGND VPWR VPWR t$5533 sky130_fd_sc_hd__a22o_1
XU$$2217 t$5538 net1430 VGND VGND VPWR VPWR booth_b32_m9 sky130_fd_sc_hd__xor2_1
XU$$2228 net1174 net570 net1165 net843 VGND VGND VPWR VPWR t$5544 sky130_fd_sc_hd__a22o_1
XFILLER_76_1111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2239 t$5549 net1432 VGND VGND VPWR VPWR booth_b32_m20 sky130_fd_sc_hd__xor2_1
XFILLER_28_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1505 t$5173 net1491 VGND VGND VPWR VPWR booth_b20_m64 sky130_fd_sc_hd__xor2_1
XU$$1516 t$5180 net1478 VGND VGND VPWR VPWR booth_b22_m1 sky130_fd_sc_hd__xor2_1
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1527 net1519 net610 net1511 net883 VGND VGND VPWR VPWR t$5186 sky130_fd_sc_hd__a22o_1
XU$$1538 t$5191 net1479 VGND VGND VPWR VPWR booth_b22_m12 sky130_fd_sc_hd__xor2_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1549 net1146 net611 net1139 net884 VGND VGND VPWR VPWR t$5197 sky130_fd_sc_hd__a22o_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0650_ clknet_leaf_165_clk booth_b34_m51 VGND VGND VPWR VPWR pp_row85_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_155_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0581_ clknet_leaf_205_clk booth_b56_m26 VGND VGND VPWR VPWR pp_row82_20 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_245_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_245_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2320_ clknet_leaf_77_clk booth_b42_m22 VGND VGND VPWR VPWR pp_row64_21 sky130_fd_sc_hd__dfxtp_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2251_ clknet_leaf_212_clk booth_b52_m10 VGND VGND VPWR VPWR pp_row62_26 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_60_5 s$539 s$541 s$543 VGND VGND VPWR VPWR c$1456 s$1457 sky130_fd_sc_hd__fa_2
XFILLER_66_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1650 net111 VGND VGND VPWR VPWR net1650 sky130_fd_sc_hd__clkbuf_4
XFILLER_78_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1202_ clknet_leaf_51_clk booth_b4_m18 VGND VGND VPWR VPWR pp_row22_2 sky130_fd_sc_hd__dfxtp_1
Xfanout1661 net110 VGND VGND VPWR VPWR net1661 sky130_fd_sc_hd__clkbuf_4
XFILLER_38_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_53_4 s$407 s$409 s$411 VGND VGND VPWR VPWR c$1370 s$1371 sky130_fd_sc_hd__fa_1
X_2182_ clknet_leaf_216_clk booth_b58_m2 VGND VGND VPWR VPWR pp_row60_29 sky130_fd_sc_hd__dfxtp_1
Xfanout1672 net1673 VGND VGND VPWR VPWR net1672 sky130_fd_sc_hd__buf_4
XU$$4120 net1125 net437 net1034 net719 VGND VGND VPWR VPWR t$6511 sky130_fd_sc_hd__a22o_1
Xfanout1683 net108 VGND VGND VPWR VPWR net1683 sky130_fd_sc_hd__buf_4
XU$$4131 t$6516 net1269 VGND VGND VPWR VPWR booth_b60_m7 sky130_fd_sc_hd__xor2_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1694 net107 VGND VGND VPWR VPWR net1694 sky130_fd_sc_hd__clkbuf_4
XU$$4142 net1205 net434 net1196 net716 VGND VGND VPWR VPWR t$6522 sky130_fd_sc_hd__a22o_1
XFILLER_66_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4153 t$6527 net1263 VGND VGND VPWR VPWR booth_b60_m18 sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_46_3 c$282 c$284 c$286 VGND VGND VPWR VPWR c$1284 s$1285 sky130_fd_sc_hd__fa_1
X_1133_ clknet_leaf_13_clk net1008 VGND VGND VPWR VPWR pp_row16_9 sky130_fd_sc_hd__dfxtp_1
XU$$4164 net1095 net436 net1085 net718 VGND VGND VPWR VPWR t$6533 sky130_fd_sc_hd__a22o_1
XFILLER_92_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4175 t$6538 net1264 VGND VGND VPWR VPWR booth_b60_m29 sky130_fd_sc_hd__xor2_1
XU$$3430 net46 net1342 VGND VGND VPWR VPWR sel_1$6158 sky130_fd_sc_hd__xor2_4
XU$$3441 net1677 net488 net1566 net761 VGND VGND VPWR VPWR t$6164 sky130_fd_sc_hd__a22o_1
XU$$4186 net988 net438 net979 net720 VGND VGND VPWR VPWR t$6544 sky130_fd_sc_hd__a22o_1
XFILLER_53_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_826 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4197 t$6549 net1271 VGND VGND VPWR VPWR booth_b60_m40 sky130_fd_sc_hd__xor2_1
XU$$3452 t$6169 net1329 VGND VGND VPWR VPWR booth_b50_m10 sky130_fd_sc_hd__xor2_1
XU$$3463 net1172 net488 net1163 net761 VGND VGND VPWR VPWR t$6175 sky130_fd_sc_hd__a22o_1
XFILLER_19_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_39_2 pp_row39_14 pp_row39_15 pp_row39_16 VGND VGND VPWR VPWR c$1198 s$1199
+ sky130_fd_sc_hd__fa_1
X_1064_ clknet_leaf_59_clk booth_b6_m3 VGND VGND VPWR VPWR pp_row9_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_65_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3474 t$6180 net1332 VGND VGND VPWR VPWR booth_b50_m21 sky130_fd_sc_hd__xor2_1
XU$$2740 net1398 VGND VGND VPWR VPWR notblock$5805\[0\] sky130_fd_sc_hd__inv_1
Xdadda_fa_5_16_1 s$2787 s$2789 s$2791 VGND VGND VPWR VPWR c$3462 s$3463 sky130_fd_sc_hd__fa_1
XU$$3485 net1068 net486 net1060 net759 VGND VGND VPWR VPWR t$6186 sky130_fd_sc_hd__a22o_1
XU$$2751 t$5811 net1376 VGND VGND VPWR VPWR booth_b40_m2 sky130_fd_sc_hd__xor2_1
XU$$3496 t$6191 net1331 VGND VGND VPWR VPWR booth_b50_m32 sky130_fd_sc_hd__xor2_1
XU$$2762 net1512 net535 net1504 net808 VGND VGND VPWR VPWR t$5817 sky130_fd_sc_hd__a22o_1
XU$$2773 t$5822 net1381 VGND VGND VPWR VPWR booth_b40_m13 sky130_fd_sc_hd__xor2_1
XFILLER_61_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2784 net1140 net536 net1132 net809 VGND VGND VPWR VPWR t$5828 sky130_fd_sc_hd__a22o_1
XU$$2795 t$5833 net1381 VGND VGND VPWR VPWR booth_b40_m24 sky130_fd_sc_hd__xor2_1
XFILLER_21_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1966_ clknet_leaf_63_clk booth_b34_m20 VGND VGND VPWR VPWR pp_row54_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_147_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0917_ clknet_leaf_103_clk booth_b60_m36 VGND VGND VPWR VPWR pp_row96_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_975 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1897_ clknet_leaf_64_clk booth_b24_m28 VGND VGND VPWR VPWR pp_row52_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0848_ clknet_leaf_109_clk booth_b46_m47 VGND VGND VPWR VPWR pp_row93_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_108_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0779_ clknet_leaf_153_clk booth_b44_m46 VGND VGND VPWR VPWR pp_row90_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_115_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_236_clk clknet_5_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_236_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_102_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_1_42_4 pp_row42_12 pp_row42_13 VGND VGND VPWR VPWR c$252 s$253 sky130_fd_sc_hd__ha_1
Xinput208 c[56] VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_1
Xinput219 c[66] VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2449_ clknet_leaf_91_clk booth_b10_m58 VGND VGND VPWR VPWR pp_row68_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_124_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$702 final_adder.p_new$726 final_adder.p_new$710 VGND VGND VPWR VPWR
+ final_adder.p_new$830 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$713 final_adder.p_new$720 final_adder.g_new$737 final_adder.g_new$721
+ VGND VGND VPWR VPWR final_adder.g_new$841 sky130_fd_sc_hd__a21o_1
XFILLER_151_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_4_12_2 pp_row12_6 pp_row12_7 VGND VGND VPWR VPWR c$2766 s$2767 sky130_fd_sc_hd__ha_1
XFILLER_84_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$735 final_adder.p_new$742 final_adder.g_new$509 final_adder.g_new$743
+ VGND VGND VPWR VPWR final_adder.g_new$863 sky130_fd_sc_hd__a21o_2
Xfinal_adder.U$$746 final_adder.p_new$794 final_adder.p_new$762 VGND VGND VPWR VPWR
+ final_adder.p_new$874 sky130_fd_sc_hd__and2_1
XFILLER_110_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$757 final_adder.p_new$772 final_adder.g_new$805 final_adder.g_new$773
+ VGND VGND VPWR VPWR final_adder.g_new$885 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$768 final_adder.p_new$816 final_adder.p_new$784 VGND VGND VPWR VPWR
+ final_adder.p_new$896 sky130_fd_sc_hd__and2_1
XFILLER_17_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$607 t$4715 net1240 VGND VGND VPWR VPWR booth_b8_m26 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$779 final_adder.p_new$794 final_adder.g_new$827 final_adder.g_new$795
+ VGND VGND VPWR VPWR final_adder.g_new$907 sky130_fd_sc_hd__a21o_1
XU$$618 net1016 net410 net998 net676 VGND VGND VPWR VPWR t$4721 sky130_fd_sc_hd__a22o_1
Xdadda_fa_1_41_2 pp_row41_6 pp_row41_7 pp_row41_8 VGND VGND VPWR VPWR c$240 s$241
+ sky130_fd_sc_hd__fa_1
XFILLER_84_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$629 t$4726 net1241 VGND VGND VPWR VPWR booth_b8_m37 sky130_fd_sc_hd__xor2_1
XFILLER_186_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_11_0 pp_row11_0 pp_row11_1 pp_row11_2 VGND VGND VPWR VPWR c$2758 s$2759
+ sky130_fd_sc_hd__fa_1
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_115_0 pp_row115_0 pp_row115_1 pp_row115_2 VGND VGND VPWR VPWR c$2746 s$2747
+ sky130_fd_sc_hd__fa_1
XFILLER_193_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_227_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_227_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_133_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_63_3 s$1487 s$1489 s$1491 VGND VGND VPWR VPWR c$2348 s$2349 sky130_fd_sc_hd__fa_1
XFILLER_43_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_56_2 c$1396 s$1399 s$1401 VGND VGND VPWR VPWR c$2290 s$2291 sky130_fd_sc_hd__fa_1
XFILLER_94_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_49_1 c$1306 c$1308 c$1310 VGND VGND VPWR VPWR c$2232 s$2233 sky130_fd_sc_hd__fa_2
XFILLER_48_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_26_0 c$3496 c$3498 s$3501 VGND VGND VPWR VPWR c$3948 s$3949 sky130_fd_sc_hd__fa_1
XU$$2003 t$5428 net1455 VGND VGND VPWR VPWR booth_b28_m39 sky130_fd_sc_hd__xor2_1
XU$$2014 net1720 net589 net1711 net862 VGND VGND VPWR VPWR t$5434 sky130_fd_sc_hd__a22o_1
XFILLER_16_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2025 t$5439 net1453 VGND VGND VPWR VPWR booth_b28_m50 sky130_fd_sc_hd__xor2_1
XFILLER_74_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2036 net1613 net589 net1605 net862 VGND VGND VPWR VPWR t$5445 sky130_fd_sc_hd__a22o_1
XFILLER_62_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1302 t$5070 net1663 VGND VGND VPWR VPWR booth_b18_m31 sky130_fd_sc_hd__xor2_1
XU$$2047 t$5450 net1455 VGND VGND VPWR VPWR booth_b28_m61 sky130_fd_sc_hd__xor2_1
XU$$1313 net969 net638 net961 net911 VGND VGND VPWR VPWR t$5076 sky130_fd_sc_hd__a22o_1
XU$$2058 net1444 notblock$5455\[1\] VGND VGND VPWR VPWR t$5456 sky130_fd_sc_hd__and2_1
XU$$2069 net937 net580 net1675 net853 VGND VGND VPWR VPWR t$5463 sky130_fd_sc_hd__a22o_1
XU$$1324 t$5081 net1667 VGND VGND VPWR VPWR booth_b18_m42 sky130_fd_sc_hd__xor2_1
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1335 net1698 net642 net1690 net915 VGND VGND VPWR VPWR t$5087 sky130_fd_sc_hd__a22o_1
XFILLER_188_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1346 t$5092 net1669 VGND VGND VPWR VPWR booth_b18_m53 sky130_fd_sc_hd__xor2_1
XU$$1357 net1587 net640 net1581 net913 VGND VGND VPWR VPWR t$5098 sky130_fd_sc_hd__a22o_1
XU$$1368 t$5103 net1668 VGND VGND VPWR VPWR booth_b18_m64 sky130_fd_sc_hd__xor2_1
XFILLER_43_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1379 t$5110 net1487 VGND VGND VPWR VPWR booth_b20_m1 sky130_fd_sc_hd__xor2_1
XFILLER_176_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1820_ clknet_leaf_220_clk booth_b48_m1 VGND VGND VPWR VPWR pp_row49_24 sky130_fd_sc_hd__dfxtp_1
XFILLER_129_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1751_ clknet_leaf_233_clk booth_b26_m21 VGND VGND VPWR VPWR pp_row47_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_117_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0702_ clknet_leaf_174_clk booth_b36_m51 VGND VGND VPWR VPWR pp_row87_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_172_945 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1682_ clknet_leaf_24_clk booth_b4_m41 VGND VGND VPWR VPWR pp_row45_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_183_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0633_ clknet_leaf_164_clk booth_b54_m63 VGND VGND VPWR VPWR pp_row117_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_125_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_218_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_218_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_98_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0564_ clknet_leaf_186_clk booth_b26_m56 VGND VGND VPWR VPWR pp_row82_5 sky130_fd_sc_hd__dfxtp_1
Xfanout909 net912 VGND VGND VPWR VPWR net909 sky130_fd_sc_hd__buf_6
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2303_ clknet_leaf_91_clk booth_b12_m52 VGND VGND VPWR VPWR pp_row64_6 sky130_fd_sc_hd__dfxtp_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0495_ clknet_leaf_158_clk booth_b56_m23 VGND VGND VPWR VPWR pp_row79_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_140_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2234_ clknet_leaf_232_clk booth_b22_m40 VGND VGND VPWR VPWR pp_row62_11 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_51_1 c$352 c$354 c$356 VGND VGND VPWR VPWR c$1340 s$1341 sky130_fd_sc_hd__fa_1
XFILLER_38_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1480 net16 VGND VGND VPWR VPWR net1480 sky130_fd_sc_hd__buf_6
Xfanout1491 net1492 VGND VGND VPWR VPWR net1491 sky130_fd_sc_hd__clkbuf_8
X_2165_ clknet_leaf_28_clk booth_b28_m32 VGND VGND VPWR VPWR pp_row60_14 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_44_0 pp_row44_17 pp_row44_18 pp_row44_19 VGND VGND VPWR VPWR c$1254 s$1255
+ sky130_fd_sc_hd__fa_1
XFILLER_81_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1116_ clknet_leaf_121_clk booth_b58_m44 VGND VGND VPWR VPWR pp_row102_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_93_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$20 c$4190 s$4193 VGND VGND VPWR VPWR final_adder.$signal$42 final_adder.$signal$1110
+ sky130_fd_sc_hd__ha_1
XU$$3260 t$6070 net1355 VGND VGND VPWR VPWR booth_b46_m51 sky130_fd_sc_hd__xor2_1
X_2096_ clknet_leaf_86_clk booth_b28_m30 VGND VGND VPWR VPWR pp_row58_14 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$31 c$4212 s$4215 VGND VGND VPWR VPWR final_adder.$signal$64 final_adder.$signal$1121
+ sky130_fd_sc_hd__ha_1
XFILLER_19_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3271 net1608 net504 net1600 net777 VGND VGND VPWR VPWR t$6076 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$42 c$4234 s$4237 VGND VGND VPWR VPWR final_adder.$signal$86 final_adder.$signal$1132
+ sky130_fd_sc_hd__ha_2
XFILLER_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3282 t$6081 net1356 VGND VGND VPWR VPWR booth_b46_m62 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$53 c$4256 s$4259 VGND VGND VPWR VPWR final_adder.$signal$108 final_adder.$signal$109
+ sky130_fd_sc_hd__ha_1
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$64 c$4278 s$4281 VGND VGND VPWR VPWR final_adder.$signal$130 final_adder.$signal$1154
+ sky130_fd_sc_hd__ha_2
X_1047_ clknet_leaf_61_clk booth_b2_m5 VGND VGND VPWR VPWR pp_row7_1 sky130_fd_sc_hd__dfxtp_1
XU$$3293 net43 net1352 VGND VGND VPWR VPWR sel_1$6088 sky130_fd_sc_hd__xor2_4
Xfinal_adder.U$$75 c$4300 s$4303 VGND VGND VPWR VPWR final_adder.$signal$152 final_adder.$signal$1165
+ sky130_fd_sc_hd__ha_2
XU$$2570 net1689 net556 net1681 net829 VGND VGND VPWR VPWR t$5718 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$86 c$4322 s$4325 VGND VGND VPWR VPWR final_adder.$signal$174 final_adder.$signal$1176
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$97 c$4344 s$4347 VGND VGND VPWR VPWR final_adder.$signal$196 final_adder.$signal$1187
+ sky130_fd_sc_hd__ha_1
XFILLER_0_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2581 t$5723 net1410 VGND VGND VPWR VPWR booth_b36_m54 sky130_fd_sc_hd__xor2_1
XU$$2592 net1585 net557 net1555 net830 VGND VGND VPWR VPWR t$5729 sky130_fd_sc_hd__a22o_1
XFILLER_139_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1880 t$5365 net1464 VGND VGND VPWR VPWR booth_b26_m46 sky130_fd_sc_hd__xor2_1
XFILLER_107_1137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1891 net1647 net598 net1638 net871 VGND VGND VPWR VPWR t$5371 sky130_fd_sc_hd__a22o_1
XFILLER_148_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1949_ clknet_leaf_137_clk booth_b46_m62 VGND VGND VPWR VPWR pp_row108_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_175_761 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_934 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_209_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_209_clk
+ sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_4_73_2 s$2425 s$2427 s$2429 VGND VGND VPWR VPWR c$3132 s$3133 sky130_fd_sc_hd__fa_1
Xdadda_fa_1_89_2 pp_row89_6 pp_row89_7 pp_row89_8 VGND VGND VPWR VPWR c$1014 s$1015
+ sky130_fd_sc_hd__fa_1
XFILLER_1_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_66_1 c$2362 c$2364 s$2367 VGND VGND VPWR VPWR c$3088 s$3089 sky130_fd_sc_hd__fa_1
XFILLER_153_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_7_43_0 s$3571 c$3980 s$3983 VGND VGND VPWR VPWR c$4238 s$4239 sky130_fd_sc_hd__fa_2
XFILLER_77_929 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_59_0 s$1445 c$2302 c$2304 VGND VGND VPWR VPWR c$3044 s$3045 sky130_fd_sc_hd__fa_1
XFILLER_130_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$510 final_adder.p_new$522 final_adder.p_new$514 VGND VGND VPWR VPWR
+ final_adder.p_new$638 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$521 final_adder.p_new$524 final_adder.g_new$533 final_adder.g_new$525
+ VGND VGND VPWR VPWR final_adder.g_new$649 sky130_fd_sc_hd__a21o_1
XTAP_3803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$532 final_adder.p_new$544 final_adder.p_new$536 VGND VGND VPWR VPWR
+ final_adder.p_new$660 sky130_fd_sc_hd__and2_1
XTAP_3814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$543 final_adder.p_new$546 final_adder.g_new$555 final_adder.g_new$547
+ VGND VGND VPWR VPWR final_adder.g_new$671 sky130_fd_sc_hd__a21o_1
XTAP_3825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$554 final_adder.p_new$566 final_adder.p_new$558 VGND VGND VPWR VPWR
+ final_adder.p_new$682 sky130_fd_sc_hd__and2_1
XTAP_3836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$404 net1547 net533 net1539 net806 VGND VGND VPWR VPWR t$4611 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$565 final_adder.p_new$568 final_adder.g_new$577 final_adder.g_new$569
+ VGND VGND VPWR VPWR final_adder.g_new$693 sky130_fd_sc_hd__a21o_1
XTAP_3847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$576 final_adder.p_new$588 final_adder.p_new$580 VGND VGND VPWR VPWR
+ final_adder.p_new$704 sky130_fd_sc_hd__and2_1
XU$$415 notblock$4615\[2\] net61 net1275 t$4616 notblock$4615\[0\] VGND VGND VPWR
+ VPWR sel_0$4617 sky130_fd_sc_hd__a32o_1
XTAP_3858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$426 t$4623 net1248 VGND VGND VPWR VPWR booth_b6_m4 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$587 final_adder.p_new$590 final_adder.g_new$599 final_adder.g_new$591
+ VGND VGND VPWR VPWR final_adder.g_new$715 sky130_fd_sc_hd__a21o_1
XTAP_3869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$437 net1496 net427 net1221 net709 VGND VGND VPWR VPWR t$4629 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$598 final_adder.p_new$610 final_adder.p_new$602 VGND VGND VPWR VPWR
+ final_adder.p_new$726 sky130_fd_sc_hd__and2_1
XFILLER_84_494 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$448 t$4634 net1248 VGND VGND VPWR VPWR booth_b6_m15 sky130_fd_sc_hd__xor2_1
XU$$459 net1114 net426 net1105 net708 VGND VGND VPWR VPWR t$4640 sky130_fd_sc_hd__a22o_1
XFILLER_71_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_717 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_61_0 s$563 c$1446 c$1448 VGND VGND VPWR VPWR c$2326 s$2327 sky130_fd_sc_hd__fa_1
XFILLER_192_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_0_77_0 pp_row77_0 pp_row77_1 pp_row77_2 VGND VGND VPWR VPWR c$200 s$201
+ sky130_fd_sc_hd__fa_1
XFILLER_79_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0280_ clknet_leaf_201_clk booth_b62_m10 VGND VGND VPWR VPWR pp_row72_28 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$960 net6 VGND VGND VPWR VPWR notblock$4895\[1\] sky130_fd_sc_hd__inv_1
Xdadda_ha_4_8_0 pp_row8_0 pp_row8_1 VGND VGND VPWR VPWR c$2750 s$2751 sky130_fd_sc_hd__ha_1
XFILLER_35_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$971 net1032 net385 net933 net651 VGND VGND VPWR VPWR t$4902 sky130_fd_sc_hd__a22o_1
XU$$1110 net936 net646 net1676 net919 VGND VGND VPWR VPWR t$4973 sky130_fd_sc_hd__a22o_1
XU$$1121 t$4978 net1008 VGND VGND VPWR VPWR booth_b16_m9 sky130_fd_sc_hd__xor2_1
XU$$982 t$4907 net1185 VGND VGND VPWR VPWR booth_b14_m8 sky130_fd_sc_hd__xor2_1
XU$$1132 net1173 net643 net1164 net916 VGND VGND VPWR VPWR t$4984 sky130_fd_sc_hd__a22o_1
XFILLER_189_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$993 net1192 net385 net1173 net651 VGND VGND VPWR VPWR t$4913 sky130_fd_sc_hd__a22o_1
XFILLER_90_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1143 t$4989 net1009 VGND VGND VPWR VPWR booth_b16_m20 sky130_fd_sc_hd__xor2_1
XU$$1154 net1071 net644 net1063 net917 VGND VGND VPWR VPWR t$4995 sky130_fd_sc_hd__a22o_1
XU$$1165 t$5000 net1007 VGND VGND VPWR VPWR booth_b16_m31 sky130_fd_sc_hd__xor2_1
XU$$1176 net969 net647 net961 net920 VGND VGND VPWR VPWR t$5006 sky130_fd_sc_hd__a22o_1
XFILLER_189_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1187 t$5011 net1011 VGND VGND VPWR VPWR booth_b16_m42 sky130_fd_sc_hd__xor2_1
XU$$1198 net1698 net650 net1690 net923 VGND VGND VPWR VPWR t$5017 sky130_fd_sc_hd__a22o_1
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1803_ clknet_leaf_220_clk booth_b18_m31 VGND VGND VPWR VPWR pp_row49_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1734_ clknet_leaf_23_clk net1348 VGND VGND VPWR VPWR pp_row46_24 sky130_fd_sc_hd__dfxtp_1
XFILLER_145_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_83_1 s$3189 s$3191 s$3193 VGND VGND VPWR VPWR c$3730 s$3731 sky130_fd_sc_hd__fa_2
XFILLER_85_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_99_1 pp_row99_3 pp_row99_4 pp_row99_5 VGND VGND VPWR VPWR c$1916 s$1917
+ sky130_fd_sc_hd__fa_1
XFILLER_105_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1665_ clknet_leaf_24_clk booth_b22_m22 VGND VGND VPWR VPWR pp_row44_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_144_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_76_0 c$3140 c$3142 c$3144 VGND VGND VPWR VPWR c$3700 s$3701 sky130_fd_sc_hd__fa_1
XFILLER_137_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0616_ clknet_leaf_187_clk booth_b20_m64 VGND VGND VPWR VPWR pp_row84_1 sky130_fd_sc_hd__dfxtp_1
X_1596_ clknet_leaf_5_clk booth_b36_m5 VGND VGND VPWR VPWR pp_row41_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_98_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout706 net707 VGND VGND VPWR VPWR net706 sky130_fd_sc_hd__clkbuf_4
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout717 net718 VGND VGND VPWR VPWR net717 sky130_fd_sc_hd__clkbuf_4
Xfanout728 net731 VGND VGND VPWR VPWR net728 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_75_8 c$188 c$190 s$193 VGND VGND VPWR VPWR c$814 s$815 sky130_fd_sc_hd__fa_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0547_ clknet_leaf_171_clk booth_b44_m37 VGND VGND VPWR VPWR pp_row81_14 sky130_fd_sc_hd__dfxtp_1
Xfanout739 net740 VGND VGND VPWR VPWR net739 sky130_fd_sc_hd__clkbuf_4
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_68_7 c$130 s$133 s$135 VGND VGND VPWR VPWR c$686 s$687 sky130_fd_sc_hd__fa_1
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0478_ clknet_leaf_193_clk booth_b24_m55 VGND VGND VPWR VPWR pp_row79_5 sky130_fd_sc_hd__dfxtp_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2217_ clknet_leaf_29_clk booth_b54_m7 VGND VGND VPWR VPWR pp_row61_27 sky130_fd_sc_hd__dfxtp_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_984 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2148_ clknet_leaf_231_clk net211 VGND VGND VPWR VPWR pp_row59_30 sky130_fd_sc_hd__dfxtp_2
XFILLER_26_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2079_ clknet_leaf_231_clk net209 VGND VGND VPWR VPWR pp_row57_29 sky130_fd_sc_hd__dfxtp_2
XU$$3090 net985 net513 net976 net786 VGND VGND VPWR VPWR t$5984 sky130_fd_sc_hd__a22o_1
XFILLER_179_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_94_0 net1903 pp_row94_1 pp_row94_2 VGND VGND VPWR VPWR c$1042 s$1043 sky130_fd_sc_hd__fa_1
XFILLER_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$340 final_adder.p_new$342 final_adder.p_new$340 VGND VGND VPWR VPWR
+ final_adder.p_new$468 sky130_fd_sc_hd__and2_1
XTAP_4367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$351 final_adder.p_new$350 final_adder.g_new$353 final_adder.g_new$351
+ VGND VGND VPWR VPWR final_adder.g_new$479 sky130_fd_sc_hd__a21o_1
XTAP_3633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_106_0 c$3816 c$3818 s$3821 VGND VGND VPWR VPWR c$4108 s$4109 sky130_fd_sc_hd__fa_1
XFILLER_29_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$201 net1047 net619 net1039 net892 VGND VGND VPWR VPWR t$4508 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$362 final_adder.p_new$364 final_adder.p_new$362 VGND VGND VPWR VPWR
+ final_adder.p_new$490 sky130_fd_sc_hd__and2_1
XTAP_4378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$373 final_adder.p_new$372 final_adder.g_new$375 final_adder.g_new$373
+ VGND VGND VPWR VPWR final_adder.g_new$501 sky130_fd_sc_hd__a21o_1
XU$$212 t$4513 net1391 VGND VGND VPWR VPWR booth_b2_m34 sky130_fd_sc_hd__xor2_1
XTAP_3655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$223 net940 net619 net924 net892 VGND VGND VPWR VPWR t$4519 sky130_fd_sc_hd__a22o_1
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$384 final_adder.p_new$390 final_adder.p_new$386 VGND VGND VPWR VPWR
+ final_adder.p_new$512 sky130_fd_sc_hd__and2_1
XTAP_3666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$234 t$4524 net1387 VGND VGND VPWR VPWR booth_b2_m45 sky130_fd_sc_hd__xor2_1
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$395 final_adder.p_new$396 final_adder.g_new$401 final_adder.g_new$397
+ VGND VGND VPWR VPWR final_adder.g_new$523 sky130_fd_sc_hd__a21o_1
XU$$245 net1658 net626 net1650 net899 VGND VGND VPWR VPWR t$4530 sky130_fd_sc_hd__a22o_1
XTAP_3677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$256 t$4535 net1392 VGND VGND VPWR VPWR booth_b2_m56 sky130_fd_sc_hd__xor2_1
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_26_3 c$1060 s$1063 s$1065 VGND VGND VPWR VPWR c$2052 s$2053 sky130_fd_sc_hd__fa_1
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$267 net1543 net621 net1535 net894 VGND VGND VPWR VPWR t$4541 sky130_fd_sc_hd__a22o_1
XU$$278 notblock$4545\[2\] net45 net1388 t$4546 notblock$4545\[0\] VGND VGND VPWR
+ VPWR sel_0$4547 sky130_fd_sc_hd__a32o_4
XTAP_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$289 t$4553 net1277 VGND VGND VPWR VPWR booth_b4_m4 sky130_fd_sc_hd__xor2_1
XFILLER_189_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_93_0 c$3764 c$3766 s$3769 VGND VGND VPWR VPWR c$4082 s$4083 sky130_fd_sc_hd__fa_1
XU$$6 net1883 net446 net1232 net688 VGND VGND VPWR VPWR t$4410 sky130_fd_sc_hd__a22o_1
XFILLER_138_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput309 net309 VGND VGND VPWR VPWR o[31] sky130_fd_sc_hd__buf_2
XFILLER_181_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1450_ clknet_leaf_110_clk booth_b60_m44 VGND VGND VPWR VPWR pp_row104_11 sky130_fd_sc_hd__dfxtp_1
X_0401_ clknet_leaf_190_clk booth_b48_m28 VGND VGND VPWR VPWR pp_row76_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_84_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1381_ clknet_leaf_43_clk booth_b18_m14 VGND VGND VPWR VPWR pp_row32_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_95_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_5_27__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_5_27__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_68_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_523 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0332_ clknet_leaf_224_clk booth_b40_m34 VGND VGND VPWR VPWR pp_row74_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_834 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0263_ clknet_leaf_150_clk booth_b34_m38 VGND VGND VPWR VPWR pp_row72_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_83_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2002_ clknet_leaf_73_clk booth_b40_m15 VGND VGND VPWR VPWR pp_row55_20 sky130_fd_sc_hd__dfxtp_1
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0194_ clknet_leaf_146_clk booth_b30_m40 VGND VGND VPWR VPWR pp_row70_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_35_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$790 t$4808 net1418 VGND VGND VPWR VPWR booth_b10_m49 sky130_fd_sc_hd__xor2_1
XFILLER_56_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_912 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1717_ clknet_leaf_21_clk booth_b18_m28 VGND VGND VPWR VPWR pp_row46_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_118_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1648_ clknet_leaf_5_clk booth_b38_m5 VGND VGND VPWR VPWR pp_row43_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_116_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_80_6 pp_row80_18 pp_row80_19 pp_row80_20 VGND VGND VPWR VPWR c$900 s$901
+ sky130_fd_sc_hd__fa_1
Xfanout503 net509 VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__buf_4
XFILLER_132_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout514 net517 VGND VGND VPWR VPWR net514 sky130_fd_sc_hd__buf_4
Xfanout525 net526 VGND VGND VPWR VPWR net525 sky130_fd_sc_hd__buf_4
X_1579_ clknet_leaf_243_clk booth_b6_m35 VGND VGND VPWR VPWR pp_row41_3 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_73_5 pp_row73_24 pp_row73_25 pp_row73_26 VGND VGND VPWR VPWR c$772 s$773
+ sky130_fd_sc_hd__fa_1
XFILLER_116_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout536 net542 VGND VGND VPWR VPWR net536 sky130_fd_sc_hd__buf_4
Xfanout547 net548 VGND VGND VPWR VPWR net547 sky130_fd_sc_hd__buf_4
XFILLER_101_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout558 net559 VGND VGND VPWR VPWR net558 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_66_4 pp_row66_30 pp_row66_31 pp_row66_32 VGND VGND VPWR VPWR c$644 s$645
+ sky130_fd_sc_hd__fa_1
Xfanout569 net570 VGND VGND VPWR VPWR net569 sky130_fd_sc_hd__buf_6
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_59_3 pp_row59_20 pp_row59_21 pp_row59_22 VGND VGND VPWR VPWR c$516 s$517
+ sky130_fd_sc_hd__fa_1
Xdadda_fa_4_36_2 s$2129 s$2131 s$2133 VGND VGND VPWR VPWR c$2910 s$2911 sky130_fd_sc_hd__fa_1
XFILLER_73_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_29_1 c$2066 c$2068 s$2071 VGND VGND VPWR VPWR c$2866 s$2867 sky130_fd_sc_hd__fa_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_0_62_5 pp_row62_15 pp_row62_16 VGND VGND VPWR VPWR c$70 s$71 sky130_fd_sc_hd__ha_2
XFILLER_135_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4505 t$6706 net1873 VGND VGND VPWR VPWR booth_b64_m57 sky130_fd_sc_hd__xor2_1
XU$$4516 net1536 sel_0$6647 net1528 net693 VGND VGND VPWR VPWR t$6712 sky130_fd_sc_hd__a22o_1
XTAP_4120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_61_3 pp_row61_9 pp_row61_10 pp_row61_11 VGND VGND VPWR VPWR c$56 s$57
+ sky130_fd_sc_hd__fa_1
XTAP_4131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3804 t$6348 net1307 VGND VGND VPWR VPWR booth_b54_m49 sky130_fd_sc_hd__xor2_1
XU$$19 t$4416 net1574 VGND VGND VPWR VPWR booth_b0_m6 sky130_fd_sc_hd__xor2_1
XTAP_4153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3815 net1624 net473 net1616 net746 VGND VGND VPWR VPWR t$6354 sky130_fd_sc_hd__a22o_1
XTAP_4164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_932 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3826 t$6359 net1306 VGND VGND VPWR VPWR booth_b54_m60 sky130_fd_sc_hd__xor2_1
XFILLER_131_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3837 net52 VGND VGND VPWR VPWR notblock$6365\[1\] sky130_fd_sc_hd__inv_1
XTAP_4186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$170 final_adder.$signal$1174 final_adder.$signal$1175 VGND VGND VPWR
+ VPWR final_adder.p_new$298 sky130_fd_sc_hd__and2_1
XTAP_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_31_1 c$1090 c$1092 c$1094 VGND VGND VPWR VPWR c$2088 s$2089 sky130_fd_sc_hd__fa_1
XU$$3848 net1037 net461 net935 net734 VGND VGND VPWR VPWR t$6372 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$181 final_adder.$signal$1165 final_adder.$signal$150 final_adder.$signal$152
+ VGND VGND VPWR VPWR final_adder.g_new$309 sky130_fd_sc_hd__a21o_1
XTAP_4197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3859 t$6377 net1296 VGND VGND VPWR VPWR booth_b56_m8 sky130_fd_sc_hd__xor2_1
XFILLER_17_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$192 final_adder.$signal$1152 final_adder.$signal$1153 VGND VGND VPWR
+ VPWR final_adder.p_new$320 sky130_fd_sc_hd__and2_1
XTAP_3474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_430 net710 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1028 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_24_0 pp_row24_5 pp_row24_6 pp_row24_7 VGND VGND VPWR VPWR c$2030 s$2031
+ sky130_fd_sc_hd__fa_1
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_441 net986 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_452 net1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_463 net1751 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0950_ clknet_leaf_114_clk booth_b48_m50 VGND VGND VPWR VPWR pp_row98_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_158_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0881_ clknet_leaf_111_clk notsign$5524 VGND VGND VPWR VPWR pp_row95_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_146_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_90_5 s$1019 s$1021 s$1023 VGND VGND VPWR VPWR c$1816 s$1817 sky130_fd_sc_hd__fa_1
XFILLER_142_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1502_ clknet_leaf_20_clk booth_b0_m38 VGND VGND VPWR VPWR pp_row38_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_99_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_83_4 s$939 s$941 s$943 VGND VGND VPWR VPWR c$1730 s$1731 sky130_fd_sc_hd__fa_1
X_2482_ clknet_leaf_142_clk booth_b6_m63 VGND VGND VPWR VPWR pp_row69_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_181_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1433_ clknet_leaf_40_clk booth_b34_m0 VGND VGND VPWR VPWR pp_row34_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_142_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_76_3 c$814 s$817 s$819 VGND VGND VPWR VPWR c$1644 s$1645 sky130_fd_sc_hd__fa_1
XFILLER_68_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_ha_1_96_0_1916 VGND VGND VPWR VPWR net1916 dadda_ha_1_96_0_1916/LO sky130_fd_sc_hd__conb_1
Xdadda_fa_2_69_2 c$682 c$684 c$686 VGND VGND VPWR VPWR c$1558 s$1559 sky130_fd_sc_hd__fa_1
X_1364_ clknet_leaf_9_clk booth_b20_m11 VGND VGND VPWR VPWR pp_row31_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_110_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_46_1 s$2967 s$2969 s$2971 VGND VGND VPWR VPWR c$3582 s$3583 sky130_fd_sc_hd__fa_1
X_0315_ clknet_leaf_197_clk net227 VGND VGND VPWR VPWR pp_row73_29 sky130_fd_sc_hd__dfxtp_1
XFILLER_68_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1295_ clknet_leaf_3_clk booth_b26_m1 VGND VGND VPWR VPWR pp_row27_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_39_0 c$2918 c$2920 c$2922 VGND VGND VPWR VPWR c$3552 s$3553 sky130_fd_sc_hd__fa_1
X_0246_ clknet_leaf_145_clk booth_b62_m9 VGND VGND VPWR VPWR pp_row71_28 sky130_fd_sc_hd__dfxtp_1
XFILLER_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_976 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0177_ clknet_leaf_100_clk booth_b62_m7 VGND VGND VPWR VPWR pp_row69_29 sky130_fd_sc_hd__dfxtp_1
XFILLER_24_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_120_1 c$3406 s$3409 s$3411 VGND VGND VPWR VPWR c$3878 s$3879 sky130_fd_sc_hd__fa_1
XFILLER_20_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_113_0 c$3362 c$3364 c$3366 VGND VGND VPWR VPWR c$3848 s$3849 sky130_fd_sc_hd__fa_1
XFILLER_192_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1309 net51 VGND VGND VPWR VPWR net1309 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_71_2 pp_row71_18 pp_row71_19 pp_row71_20 VGND VGND VPWR VPWR c$730 s$731
+ sky130_fd_sc_hd__fa_1
XFILLER_120_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_64_1 pp_row64_21 pp_row64_22 pp_row64_23 VGND VGND VPWR VPWR c$602 s$603
+ sky130_fd_sc_hd__fa_2
Xclkbuf_5_10__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_5_10__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xfanout388 net389 VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__clkbuf_4
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_41_0 s$1229 c$2158 c$2160 VGND VGND VPWR VPWR c$2936 s$2937 sky130_fd_sc_hd__fa_1
Xfanout399 net400 VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__clkbuf_8
XFILLER_46_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_57_0 pp_row57_8 pp_row57_9 pp_row57_10 VGND VGND VPWR VPWR c$474 s$475
+ sky130_fd_sc_hd__fa_1
XFILLER_189_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1709 t$5278 net1470 VGND VGND VPWR VPWR booth_b24_m29 sky130_fd_sc_hd__xor2_1
XFILLER_15_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput19 a[26] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_93_3 s$1847 s$1849 s$1851 VGND VGND VPWR VPWR c$2588 s$2589 sky130_fd_sc_hd__fa_2
XFILLER_182_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_86_2 c$1756 s$1759 s$1761 VGND VGND VPWR VPWR c$2530 s$2531 sky130_fd_sc_hd__fa_1
XFILLER_163_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_79_1 c$1666 c$1668 c$1670 VGND VGND VPWR VPWR c$2472 s$2473 sky130_fd_sc_hd__fa_1
XFILLER_112_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_789 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_56_0 c$3616 c$3618 s$3621 VGND VGND VPWR VPWR c$4008 s$4009 sky130_fd_sc_hd__fa_1
XFILLER_105_992 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4302 t$6603 net1256 VGND VGND VPWR VPWR booth_b62_m24 sky130_fd_sc_hd__xor2_1
XU$$4313 net1045 net425 net1029 net707 VGND VGND VPWR VPWR t$6609 sky130_fd_sc_hd__a22o_1
XFILLER_42_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4324 t$6614 net1261 VGND VGND VPWR VPWR booth_b62_m35 sky130_fd_sc_hd__xor2_1
XU$$4335 net929 net423 net1750 net705 VGND VGND VPWR VPWR t$6620 sky130_fd_sc_hd__a22o_1
XFILLER_120_995 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3601 t$6245 net1324 VGND VGND VPWR VPWR booth_b52_m16 sky130_fd_sc_hd__xor2_1
XU$$4346 t$6625 net1256 VGND VGND VPWR VPWR booth_b62_m46 sky130_fd_sc_hd__xor2_1
XU$$3612 net1111 net476 net1102 net749 VGND VGND VPWR VPWR t$6251 sky130_fd_sc_hd__a22o_1
XU$$4357 net1653 net423 net1645 net705 VGND VGND VPWR VPWR t$6631 sky130_fd_sc_hd__a22o_1
XU$$3623 t$6256 net1322 VGND VGND VPWR VPWR booth_b52_m27 sky130_fd_sc_hd__xor2_1
XU$$4368 t$6636 net1261 VGND VGND VPWR VPWR booth_b62_m57 sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_115_2 c$2742 c$2744 s$2747 VGND VGND VPWR VPWR c$3384 s$3385 sky130_fd_sc_hd__fa_1
X_1080_ clknet_leaf_52_clk booth_b8_m3 VGND VGND VPWR VPWR pp_row11_4 sky130_fd_sc_hd__dfxtp_1
XU$$3634 net1003 net477 net995 net750 VGND VGND VPWR VPWR t$6262 sky130_fd_sc_hd__a22o_1
XU$$4379 net1536 net419 net1528 net701 VGND VGND VPWR VPWR t$6642 sky130_fd_sc_hd__a22o_1
XU$$2900 t$5887 net1372 VGND VGND VPWR VPWR booth_b42_m8 sky130_fd_sc_hd__xor2_1
XU$$3645 t$6267 net1327 VGND VGND VPWR VPWR booth_b52_m38 sky130_fd_sc_hd__xor2_1
XU$$2911 net1200 net523 net1181 net796 VGND VGND VPWR VPWR t$5893 sky130_fd_sc_hd__a22o_1
XU$$3656 net1734 net482 net1726 net755 VGND VGND VPWR VPWR t$6273 sky130_fd_sc_hd__a22o_1
XFILLER_34_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2922 t$5898 net1368 VGND VGND VPWR VPWR booth_b42_m19 sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_108_1 c$2698 c$2700 s$2703 VGND VGND VPWR VPWR c$3340 s$3341 sky130_fd_sc_hd__fa_1
XTAP_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3667 t$6278 net1326 VGND VGND VPWR VPWR booth_b52_m49 sky130_fd_sc_hd__xor2_1
XTAP_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2933 net1087 net526 net1078 net799 VGND VGND VPWR VPWR t$5904 sky130_fd_sc_hd__a22o_1
XU$$3678 net1624 net478 net1616 net751 VGND VGND VPWR VPWR t$6284 sky130_fd_sc_hd__a22o_1
XU$$2944 t$5909 net1367 VGND VGND VPWR VPWR booth_b42_m30 sky130_fd_sc_hd__xor2_1
XU$$3689 t$6289 net1327 VGND VGND VPWR VPWR booth_b52_m60 sky130_fd_sc_hd__xor2_1
XTAP_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2955 net975 net521 net966 net794 VGND VGND VPWR VPWR t$5915 sky130_fd_sc_hd__a22o_1
XTAP_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2966 t$5920 net1369 VGND VGND VPWR VPWR booth_b42_m41 sky130_fd_sc_hd__xor2_1
XFILLER_60_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2977 net1705 net522 net1697 net795 VGND VGND VPWR VPWR t$5926 sky130_fd_sc_hd__a22o_1
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_260 net1667 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_271 net1744 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2988 t$5931 net1373 VGND VGND VPWR VPWR booth_b42_m52 sky130_fd_sc_hd__xor2_1
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2999 net1602 net524 net1592 net797 VGND VGND VPWR VPWR t$5937 sky130_fd_sc_hd__a22o_1
XANTENNA_282 final_adder.p_new$840 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_293 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1982_ clknet_leaf_78_clk booth_b4_m51 VGND VGND VPWR VPWR pp_row55_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_14_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0933_ clknet_leaf_112_clk booth_b52_m45 VGND VGND VPWR VPWR pp_row97_10 sky130_fd_sc_hd__dfxtp_1
XU$$4397_1819 VGND VGND VPWR VPWR U$$4397_1819/HI net1819 sky130_fd_sc_hd__conb_1
XFILLER_14_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0864_ clknet_leaf_111_clk booth_b38_m56 VGND VGND VPWR VPWR pp_row94_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_146_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0795_ clknet_leaf_139_clk booth_b32_m59 VGND VGND VPWR VPWR pp_row91_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_170_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$691_1885 VGND VGND VPWR VPWR U$$691_1885/HI net1885 sky130_fd_sc_hd__conb_1
Xdadda_fa_2_81_1 c$890 c$892 c$894 VGND VGND VPWR VPWR c$1700 s$1701 sky130_fd_sc_hd__fa_1
XFILLER_114_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1055 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2465_ clknet_leaf_95_clk booth_b40_m28 VGND VGND VPWR VPWR pp_row68_19 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_74_0 s$191 c$762 c$764 VGND VGND VPWR VPWR c$1614 s$1615 sky130_fd_sc_hd__fa_1
XFILLER_87_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1416_ clknet_leaf_56_clk booth_b4_m30 VGND VGND VPWR VPWR pp_row34_2 sky130_fd_sc_hd__dfxtp_1
X_2396_ clknet_leaf_96_clk booth_b46_m20 VGND VGND VPWR VPWR pp_row66_23 sky130_fd_sc_hd__dfxtp_1
XFILLER_60_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$906 final_adder.$signal$1200 final_adder.g_new$981 final_adder.$signal$222
+ VGND VGND VPWR VPWR final_adder.g_new$1034 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$917 final_adder.$signal$1178 final_adder.g_new$1003 final_adder.$signal$178
+ VGND VGND VPWR VPWR final_adder.g_new$1045 sky130_fd_sc_hd__a21o_1
XFILLER_69_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$928 final_adder.$signal$1156 final_adder.g_new$1025 final_adder.$signal$134
+ VGND VGND VPWR VPWR final_adder.g_new$1056 sky130_fd_sc_hd__a21o_1
X_1347_ clknet_leaf_3_clk booth_b26_m4 VGND VGND VPWR VPWR pp_row30_13 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$939 final_adder.$signal$1134 final_adder.g_new$951 final_adder.$signal$90
+ VGND VGND VPWR VPWR final_adder.g_new$1067 sky130_fd_sc_hd__a21o_1
Xdadda_fa_1_50_7 pp_row50_21 pp_row50_22 pp_row50_23 VGND VGND VPWR VPWR c$362 s$363
+ sky130_fd_sc_hd__fa_1
XFILLER_3_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1278_ clknet_leaf_244_clk net175 VGND VGND VPWR VPWR pp_row26_15 sky130_fd_sc_hd__dfxtp_2
X_0229_ clknet_leaf_153_clk booth_b32_m39 VGND VGND VPWR VPWR pp_row71_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_1075 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4421_1831 VGND VGND VPWR VPWR U$$4421_1831/HI net1831 sky130_fd_sc_hd__conb_1
XFILLER_165_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_96_1 c$2602 c$2604 s$2607 VGND VGND VPWR VPWR c$3268 s$3269 sky130_fd_sc_hd__fa_1
XFILLER_137_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_73_0 s$3691 c$4040 s$4043 VGND VGND VPWR VPWR c$4298 s$4299 sky130_fd_sc_hd__fa_1
XFILLER_121_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_89_0 s$1805 c$2542 c$2544 VGND VGND VPWR VPWR c$3224 s$3225 sky130_fd_sc_hd__fa_1
XFILLER_118_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1106 net1110 VGND VGND VPWR VPWR net1106 sky130_fd_sc_hd__clkbuf_4
Xfanout1117 net1118 VGND VGND VPWR VPWR net1117 sky130_fd_sc_hd__buf_4
Xfanout1128 net76 VGND VGND VPWR VPWR net1128 sky130_fd_sc_hd__clkbuf_4
Xfanout1139 net1140 VGND VGND VPWR VPWR net1139 sky130_fd_sc_hd__buf_4
XFILLER_102_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2207 t$5533 net1432 VGND VGND VPWR VPWR booth_b32_m4 sky130_fd_sc_hd__xor2_1
XFILLER_34_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2218 net1494 net569 net1219 net842 VGND VGND VPWR VPWR t$5539 sky130_fd_sc_hd__a22o_1
XFILLER_27_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2229 t$5544 net1431 VGND VGND VPWR VPWR booth_b32_m15 sky130_fd_sc_hd__xor2_1
XFILLER_55_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1506 net1491 VGND VGND VPWR VPWR notsign$5174 sky130_fd_sc_hd__inv_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1517 net1123 net610 net1032 net883 VGND VGND VPWR VPWR t$5181 sky130_fd_sc_hd__a22o_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1528 t$5186 net1475 VGND VGND VPWR VPWR booth_b22_m7 sky130_fd_sc_hd__xor2_1
XFILLER_15_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1539 net1206 net614 net1198 net887 VGND VGND VPWR VPWR t$5192 sky130_fd_sc_hd__a22o_1
XFILLER_188_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_190_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_190_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_91_0 s$1031 c$1806 c$1808 VGND VGND VPWR VPWR c$2566 s$2567 sky130_fd_sc_hd__fa_1
XFILLER_6_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0580_ clknet_leaf_189_clk booth_b54_m28 VGND VGND VPWR VPWR pp_row82_19 sky130_fd_sc_hd__dfxtp_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2250_ clknet_leaf_149_clk booth_b50_m12 VGND VGND VPWR VPWR pp_row62_25 sky130_fd_sc_hd__dfxtp_1
XFILLER_111_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_759 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1640 net112 VGND VGND VPWR VPWR net1640 sky130_fd_sc_hd__buf_6
X_1201_ clknet_leaf_49_clk booth_b2_m20 VGND VGND VPWR VPWR pp_row22_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_66_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1651 net1653 VGND VGND VPWR VPWR net1651 sky130_fd_sc_hd__buf_4
Xfanout1662 net1667 VGND VGND VPWR VPWR net1662 sky130_fd_sc_hd__buf_6
X_2181_ clknet_leaf_218_clk booth_b56_m4 VGND VGND VPWR VPWR pp_row60_28 sky130_fd_sc_hd__dfxtp_1
XU$$4110 net1284 VGND VGND VPWR VPWR notblock$6505\[0\] sky130_fd_sc_hd__inv_1
Xdadda_fa_2_53_5 s$413 s$415 s$417 VGND VGND VPWR VPWR c$1372 s$1373 sky130_fd_sc_hd__fa_1
XFILLER_38_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_120_0 net1913 pp_row120_1 pp_row120_2 VGND VGND VPWR VPWR c$3408 s$3409
+ sky130_fd_sc_hd__fa_1
Xfanout1673 net1674 VGND VGND VPWR VPWR net1673 sky130_fd_sc_hd__clkbuf_4
XU$$4121 t$6511 net1264 VGND VGND VPWR VPWR booth_b60_m2 sky130_fd_sc_hd__xor2_1
XU$$4132 net1517 net438 net127 net720 VGND VGND VPWR VPWR t$6517 sky130_fd_sc_hd__a22o_1
Xfanout1684 net1686 VGND VGND VPWR VPWR net1684 sky130_fd_sc_hd__buf_4
XFILLER_77_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4143 t$6522 net1263 VGND VGND VPWR VPWR booth_b60_m13 sky130_fd_sc_hd__xor2_1
Xfanout1695 net1697 VGND VGND VPWR VPWR net1695 sky130_fd_sc_hd__buf_6
X_1132_ clknet_leaf_13_clk booth_b16_m0 VGND VGND VPWR VPWR pp_row16_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_65_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4154 net1142 net436 net1135 net718 VGND VGND VPWR VPWR t$6528 sky130_fd_sc_hd__a22o_1
XFILLER_168_1015 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4165 t$6533 net1268 VGND VGND VPWR VPWR booth_b60_m24 sky130_fd_sc_hd__xor2_1
XFILLER_19_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_46_4 s$289 s$291 s$293 VGND VGND VPWR VPWR c$1286 s$1287 sky130_fd_sc_hd__fa_2
XU$$3420 net1541 net499 net1532 net772 VGND VGND VPWR VPWR t$6152 sky130_fd_sc_hd__a22o_1
XU$$3431 net1793 net484 net1228 net757 VGND VGND VPWR VPWR t$6159 sky130_fd_sc_hd__a22o_1
XU$$4176 net1045 net439 net1029 net721 VGND VGND VPWR VPWR t$6539 sky130_fd_sc_hd__a22o_1
XU$$4187 t$6544 net1269 VGND VGND VPWR VPWR booth_b60_m35 sky130_fd_sc_hd__xor2_1
XU$$3442 t$6164 net1333 VGND VGND VPWR VPWR booth_b50_m5 sky130_fd_sc_hd__xor2_1
XU$$4198 net929 net440 net1750 net722 VGND VGND VPWR VPWR t$6550 sky130_fd_sc_hd__a22o_1
X_1063_ clknet_leaf_60_clk booth_b4_m5 VGND VGND VPWR VPWR pp_row9_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_53_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3453 net1222 net484 net1214 net757 VGND VGND VPWR VPWR t$6170 sky130_fd_sc_hd__a22o_1
XFILLER_65_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3464 t$6175 net1333 VGND VGND VPWR VPWR booth_b50_m16 sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_39_3 pp_row39_17 pp_row39_18 pp_row39_19 VGND VGND VPWR VPWR c$1200 s$1201
+ sky130_fd_sc_hd__fa_1
XU$$2730 t$5799 net1400 VGND VGND VPWR VPWR booth_b38_m60 sky130_fd_sc_hd__xor2_1
XU$$3475 net1107 net484 net1098 net757 VGND VGND VPWR VPWR t$6181 sky130_fd_sc_hd__a22o_1
XU$$2741 net35 VGND VGND VPWR VPWR notblock$5805\[1\] sky130_fd_sc_hd__inv_1
XFILLER_92_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3486 t$6186 net1330 VGND VGND VPWR VPWR booth_b50_m27 sky130_fd_sc_hd__xor2_1
XTAP_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2752 net1031 net535 net934 net808 VGND VGND VPWR VPWR t$5812 sky130_fd_sc_hd__a22o_1
XU$$3497 net1003 net485 net995 net758 VGND VGND VPWR VPWR t$6192 sky130_fd_sc_hd__a22o_1
XFILLER_34_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2763 t$5817 net1376 VGND VGND VPWR VPWR booth_b40_m8 sky130_fd_sc_hd__xor2_1
XFILLER_179_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2774 net1199 net539 net1181 net812 VGND VGND VPWR VPWR t$5823 sky130_fd_sc_hd__a22o_1
XU$$2785 t$5828 net1377 VGND VGND VPWR VPWR booth_b40_m19 sky130_fd_sc_hd__xor2_1
XU$$2796 net1084 net539 net1075 net812 VGND VGND VPWR VPWR t$5834 sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_181_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_181_clk
+ sky130_fd_sc_hd__clkbuf_16
X_1965_ clknet_leaf_62_clk booth_b32_m22 VGND VGND VPWR VPWR pp_row54_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0916_ clknet_leaf_103_clk booth_b58_m38 VGND VGND VPWR VPWR pp_row96_14 sky130_fd_sc_hd__dfxtp_1
X_1896_ clknet_leaf_64_clk booth_b22_m30 VGND VGND VPWR VPWR pp_row52_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0847_ clknet_leaf_105_clk booth_b44_m49 VGND VGND VPWR VPWR pp_row93_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_161_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0778_ clknet_leaf_153_clk booth_b42_m48 VGND VGND VPWR VPWR pp_row90_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_1_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4451_1846 VGND VGND VPWR VPWR U$$4451_1846/HI net1846 sky130_fd_sc_hd__conb_1
XFILLER_130_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput209 c[57] VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_1
X_2448_ clknet_leaf_91_clk booth_b8_m60 VGND VGND VPWR VPWR pp_row68_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_75_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$703 final_adder.p_new$710 final_adder.g_new$727 final_adder.g_new$711
+ VGND VGND VPWR VPWR final_adder.g_new$831 sky130_fd_sc_hd__a21o_1
XFILLER_69_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$714 final_adder.p_new$738 final_adder.p_new$722 VGND VGND VPWR VPWR
+ final_adder.p_new$842 sky130_fd_sc_hd__and2_1
X_2379_ clknet_leaf_83_clk booth_b18_m48 VGND VGND VPWR VPWR pp_row66_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_111_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$725 final_adder.p_new$732 final_adder.g_new$749 final_adder.g_new$733
+ VGND VGND VPWR VPWR final_adder.g_new$853 sky130_fd_sc_hd__a21o_2
Xfinal_adder.U$$747 final_adder.p_new$762 final_adder.g_new$795 final_adder.g_new$763
+ VGND VGND VPWR VPWR final_adder.g_new$875 sky130_fd_sc_hd__a21o_1
XFILLER_84_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$758 final_adder.p_new$806 final_adder.p_new$774 VGND VGND VPWR VPWR
+ final_adder.p_new$886 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$769 final_adder.p_new$784 final_adder.g_new$817 final_adder.g_new$785
+ VGND VGND VPWR VPWR final_adder.g_new$897 sky130_fd_sc_hd__a21o_1
XU$$608 net1066 net413 net1058 net679 VGND VGND VPWR VPWR t$4716 sky130_fd_sc_hd__a22o_1
XU$$619 t$4721 net1236 VGND VGND VPWR VPWR booth_b8_m32 sky130_fd_sc_hd__xor2_1
XFILLER_16_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_172_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_172_clk
+ sky130_fd_sc_hd__clkbuf_16
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_913 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_108_0 pp_row108_2 pp_row108_3 pp_row108_4 VGND VGND VPWR VPWR c$2702 s$2703
+ sky130_fd_sc_hd__fa_1
XFILLER_165_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_5_8__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_5_8__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_106_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_895 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_56_3 s$1403 s$1405 s$1407 VGND VGND VPWR VPWR c$2292 s$2293 sky130_fd_sc_hd__fa_1
XFILLER_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_49_2 c$1312 s$1315 s$1317 VGND VGND VPWR VPWR c$2234 s$2235 sky130_fd_sc_hd__fa_1
XFILLER_63_805 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2004 net942 net591 net926 net864 VGND VGND VPWR VPWR t$5429 sky130_fd_sc_hd__a22o_1
XU$$2015 t$5434 net1450 VGND VGND VPWR VPWR booth_b28_m45 sky130_fd_sc_hd__xor2_1
XFILLER_74_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2026 net1655 net589 net1647 net862 VGND VGND VPWR VPWR t$5440 sky130_fd_sc_hd__a22o_1
Xdadda_fa_6_19_0 c$3468 c$3470 s$3473 VGND VGND VPWR VPWR c$3934 s$3935 sky130_fd_sc_hd__fa_1
XU$$2037 t$5445 net1453 VGND VGND VPWR VPWR booth_b28_m56 sky130_fd_sc_hd__xor2_1
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1303 net1015 net639 net998 net912 VGND VGND VPWR VPWR t$5071 sky130_fd_sc_hd__a22o_1
XU$$2048 net1548 net592 net1540 net865 VGND VGND VPWR VPWR t$5451 sky130_fd_sc_hd__a22o_1
XFILLER_188_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2059 notblock$5455\[2\] net24 net1454 t$5456 notblock$5455\[0\] VGND VGND VPWR
+ VPWR sel_0$5457 sky130_fd_sc_hd__a32o_1
XU$$1314 t$5076 net1666 VGND VGND VPWR VPWR booth_b18_m37 sky130_fd_sc_hd__xor2_1
XU$$1325 net1737 net636 net1729 net909 VGND VGND VPWR VPWR t$5082 sky130_fd_sc_hd__a22o_1
XFILLER_71_860 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1336 t$5087 net1667 VGND VGND VPWR VPWR booth_b18_m48 sky130_fd_sc_hd__xor2_1
XFILLER_167_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1347 net1629 net640 net1620 net913 VGND VGND VPWR VPWR t$5093 sky130_fd_sc_hd__a22o_1
XFILLER_71_882 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1358 t$5098 net1668 VGND VGND VPWR VPWR booth_b18_m59 sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_163_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_163_clk
+ sky130_fd_sc_hd__clkbuf_16
XU$$1369 net1668 VGND VGND VPWR VPWR notsign$5104 sky130_fd_sc_hd__inv_1
XFILLER_43_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1750_ clknet_leaf_123_clk booth_b60_m46 VGND VGND VPWR VPWR pp_row106_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_12_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0701_ clknet_leaf_174_clk booth_b34_m53 VGND VGND VPWR VPWR pp_row87_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_128_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1681_ clknet_leaf_24_clk booth_b2_m43 VGND VGND VPWR VPWR pp_row45_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_7_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_957 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0632_ clknet_leaf_178_clk booth_b50_m34 VGND VGND VPWR VPWR pp_row84_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0563_ clknet_leaf_186_clk booth_b24_m58 VGND VGND VPWR VPWR pp_row82_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2302_ clknet_leaf_198_clk booth_b10_m54 VGND VGND VPWR VPWR pp_row64_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_97_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0494_ clknet_leaf_159_clk booth_b54_m25 VGND VGND VPWR VPWR pp_row79_20 sky130_fd_sc_hd__dfxtp_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2233_ clknet_leaf_233_clk booth_b20_m42 VGND VGND VPWR VPWR pp_row62_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_57_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_51_2 c$358 c$360 c$362 VGND VGND VPWR VPWR c$1342 s$1343 sky130_fd_sc_hd__fa_1
Xfanout1470 net18 VGND VGND VPWR VPWR net1470 sky130_fd_sc_hd__buf_6
XFILLER_94_941 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1481 net1482 VGND VGND VPWR VPWR net1481 sky130_fd_sc_hd__buf_4
XFILLER_39_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2164_ clknet_leaf_29_clk booth_b26_m34 VGND VGND VPWR VPWR pp_row60_13 sky130_fd_sc_hd__dfxtp_1
Xfanout1492 net1493 VGND VGND VPWR VPWR net1492 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_44_1 pp_row44_20 pp_row44_21 pp_row44_22 VGND VGND VPWR VPWR c$1256 s$1257
+ sky130_fd_sc_hd__fa_1
XFILLER_94_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1115_ clknet_leaf_47_clk booth_b4_m11 VGND VGND VPWR VPWR pp_row15_2 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$10 c$4170 s$4173 VGND VGND VPWR VPWR final_adder.$signal$22 final_adder.$signal$1100
+ sky130_fd_sc_hd__ha_1
XFILLER_66_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3250 t$6065 net1355 VGND VGND VPWR VPWR booth_b46_m46 sky130_fd_sc_hd__xor2_1
XFILLER_0_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2095_ clknet_leaf_88_clk booth_b26_m32 VGND VGND VPWR VPWR pp_row58_13 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_21_0 c$2810 c$2812 c$2814 VGND VGND VPWR VPWR c$3480 s$3481 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$21 c$4192 s$4195 VGND VGND VPWR VPWR final_adder.$signal$44 final_adder.$signal$1111
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_2_37_0 pp_row37_5 pp_row37_6 pp_row37_7 VGND VGND VPWR VPWR c$1170 s$1171
+ sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$32 c$4214 s$4217 VGND VGND VPWR VPWR final_adder.$signal$66 final_adder.$signal$1122
+ sky130_fd_sc_hd__ha_2
XU$$3261 net1652 net507 net1644 net780 VGND VGND VPWR VPWR t$6071 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$43 c$4236 s$4239 VGND VGND VPWR VPWR final_adder.$signal$88 final_adder.$signal$1133
+ sky130_fd_sc_hd__ha_1
XFILLER_0_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3272 t$6076 net1350 VGND VGND VPWR VPWR booth_b46_m57 sky130_fd_sc_hd__xor2_1
X_1046_ clknet_leaf_61_clk booth_b0_m7 VGND VGND VPWR VPWR pp_row7_0 sky130_fd_sc_hd__dfxtp_1
XU$$3283 net1540 net508 net1532 net781 VGND VGND VPWR VPWR t$6082 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$54 c$4258 s$4261 VGND VGND VPWR VPWR final_adder.$signal$110 final_adder.$signal$111
+ sky130_fd_sc_hd__ha_1
XU$$3294 net1791 net493 net1229 net766 VGND VGND VPWR VPWR t$6089 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$65 c$4280 s$4283 VGND VGND VPWR VPWR final_adder.$signal$132 final_adder.$signal$1155
+ sky130_fd_sc_hd__ha_2
XU$$2560 net1731 net555 net1722 net828 VGND VGND VPWR VPWR t$5713 sky130_fd_sc_hd__a22o_1
XFILLER_55_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$76 c$4302 s$4305 VGND VGND VPWR VPWR final_adder.$signal$154 final_adder.$signal$1166
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$87 c$4324 s$4327 VGND VGND VPWR VPWR final_adder.$signal$176 final_adder.$signal$1177
+ sky130_fd_sc_hd__ha_1
XFILLER_179_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$98 c$4346 s$4349 VGND VGND VPWR VPWR final_adder.$signal$198 final_adder.$signal$1188
+ sky130_fd_sc_hd__ha_1
XU$$2571 t$5718 net1411 VGND VGND VPWR VPWR booth_b36_m49 sky130_fd_sc_hd__xor2_1
XFILLER_94_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_154_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_154_clk
+ sky130_fd_sc_hd__clkbuf_16
XU$$2582 net1624 net557 net1616 net830 VGND VGND VPWR VPWR t$5724 sky130_fd_sc_hd__a22o_1
XU$$2593 t$5729 net1410 VGND VGND VPWR VPWR booth_b36_m60 sky130_fd_sc_hd__xor2_1
XFILLER_22_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1870 t$5360 net1465 VGND VGND VPWR VPWR booth_b26_m41 sky130_fd_sc_hd__xor2_1
XFILLER_22_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1881 net1703 net598 net1695 net871 VGND VGND VPWR VPWR t$5366 sky130_fd_sc_hd__a22o_1
XFILLER_21_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1892 t$5371 net1464 VGND VGND VPWR VPWR booth_b26_m52 sky130_fd_sc_hd__xor2_1
XFILLER_107_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1948_ clknet_leaf_78_clk booth_b4_m50 VGND VGND VPWR VPWR pp_row54_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_163_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_829 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1879_ clknet_leaf_70_clk booth_b46_m5 VGND VGND VPWR VPWR pp_row51_23 sky130_fd_sc_hd__dfxtp_1
XFILLER_163_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_89_3 pp_row89_9 pp_row89_10 pp_row89_11 VGND VGND VPWR VPWR c$1016 s$1017
+ sky130_fd_sc_hd__fa_1
XFILLER_27_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_66_2 s$2369 s$2371 s$2373 VGND VGND VPWR VPWR c$3090 s$3091 sky130_fd_sc_hd__fa_1
XFILLER_135_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_59_1 c$2306 c$2308 s$2311 VGND VGND VPWR VPWR c$3046 s$3047 sky130_fd_sc_hd__fa_1
XFILLER_88_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$500 final_adder.p_new$506 final_adder.p_new$502 VGND VGND VPWR VPWR
+ final_adder.p_new$628 sky130_fd_sc_hd__and2_1
Xdadda_fa_7_36_0 s$3543 c$3966 s$3969 VGND VGND VPWR VPWR c$4224 s$4225 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$511 final_adder.p_new$514 final_adder.g_new$523 final_adder.g_new$515
+ VGND VGND VPWR VPWR final_adder.g_new$639 sky130_fd_sc_hd__a21o_1
XFILLER_85_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$522 final_adder.p_new$534 final_adder.p_new$526 VGND VGND VPWR VPWR
+ final_adder.p_new$650 sky130_fd_sc_hd__and2_1
XTAP_3804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$533 final_adder.p_new$536 final_adder.g_new$545 final_adder.g_new$537
+ VGND VGND VPWR VPWR final_adder.g_new$661 sky130_fd_sc_hd__a21o_1
XTAP_3815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$544 final_adder.p_new$556 final_adder.p_new$548 VGND VGND VPWR VPWR
+ final_adder.p_new$672 sky130_fd_sc_hd__and2_1
XTAP_3826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$555 final_adder.p_new$558 final_adder.g_new$567 final_adder.g_new$559
+ VGND VGND VPWR VPWR final_adder.g_new$683 sky130_fd_sc_hd__a21o_1
XTAP_3837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$405 t$4611 net1280 VGND VGND VPWR VPWR booth_b4_m62 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$566 final_adder.p_new$578 final_adder.p_new$570 VGND VGND VPWR VPWR
+ final_adder.p_new$694 sky130_fd_sc_hd__and2_1
XFILLER_151_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$577 final_adder.p_new$580 final_adder.g_new$589 final_adder.g_new$581
+ VGND VGND VPWR VPWR final_adder.g_new$705 sky130_fd_sc_hd__a21o_1
XU$$416 net61 net1275 VGND VGND VPWR VPWR sel_1$4618 sky130_fd_sc_hd__xor2_1
XTAP_3859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$427 net1676 net430 net1564 net712 VGND VGND VPWR VPWR t$4624 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$588 final_adder.p_new$600 final_adder.p_new$592 VGND VGND VPWR VPWR
+ final_adder.p_new$716 sky130_fd_sc_hd__and2_1
XU$$438 t$4629 net1245 VGND VGND VPWR VPWR booth_b6_m10 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$599 final_adder.p_new$602 final_adder.g_new$611 final_adder.g_new$603
+ VGND VGND VPWR VPWR final_adder.g_new$727 sky130_fd_sc_hd__a21o_1
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$449 net1170 net429 net1161 net711 VGND VGND VPWR VPWR t$4635 sky130_fd_sc_hd__a22o_1
XFILLER_71_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_145_clk clknet_5_25__leaf_clk VGND VGND VPWR VPWR clknet_leaf_145_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_12_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_61_1 c$1450 c$1452 c$1454 VGND VGND VPWR VPWR c$2328 s$2329 sky130_fd_sc_hd__fa_1
XFILLER_192_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_54_0 s$437 c$1362 c$1364 VGND VGND VPWR VPWR c$2270 s$2271 sky130_fd_sc_hd__fa_1
XFILLER_134_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$950 net1551 net395 net1543 net661 VGND VGND VPWR VPWR t$4890 sky130_fd_sc_hd__a22o_1
XFILLER_63_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1100 notblock$4965\[2\] net8 net1188 t$4966 notblock$4965\[0\] VGND VGND VPWR
+ VPWR sel_0$4967 sky130_fd_sc_hd__a32o_2
XFILLER_189_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$961 net1189 VGND VGND VPWR VPWR notblock$4895\[2\] sky130_fd_sc_hd__inv_1
XU$$972 t$4902 net1183 VGND VGND VPWR VPWR booth_b14_m3 sky130_fd_sc_hd__xor2_1
XU$$1111 t$4973 net1009 VGND VGND VPWR VPWR booth_b16_m4 sky130_fd_sc_hd__xor2_1
XU$$1122 net1494 net643 net1219 net916 VGND VGND VPWR VPWR t$4979 sky130_fd_sc_hd__a22o_1
XU$$983 net1505 net387 net1496 net653 VGND VGND VPWR VPWR t$4908 sky130_fd_sc_hd__a22o_1
XU$$994 t$4913 net1183 VGND VGND VPWR VPWR booth_b14_m14 sky130_fd_sc_hd__xor2_1
XU$$1133 t$4984 net1006 VGND VGND VPWR VPWR booth_b16_m15 sky130_fd_sc_hd__xor2_1
XFILLER_90_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1144 net1115 net645 net1106 net918 VGND VGND VPWR VPWR t$4990 sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_136_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_136_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_189_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1155 t$4995 net1006 VGND VGND VPWR VPWR booth_b16_m26 sky130_fd_sc_hd__xor2_1
XU$$1166 net1015 net644 net998 net917 VGND VGND VPWR VPWR t$5001 sky130_fd_sc_hd__a22o_1
XU$$1177 t$5006 net1010 VGND VGND VPWR VPWR booth_b16_m37 sky130_fd_sc_hd__xor2_1
XFILLER_176_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1188 net1738 net648 net1730 net921 VGND VGND VPWR VPWR t$5012 sky130_fd_sc_hd__a22o_1
XU$$1199 t$5017 net1014 VGND VGND VPWR VPWR booth_b16_m48 sky130_fd_sc_hd__xor2_1
X_1802_ clknet_leaf_219_clk booth_b16_m33 VGND VGND VPWR VPWR pp_row49_8 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_7_111_0 s$3843 c$4116 s$4119 VGND VGND VPWR VPWR c$4374 s$4375 sky130_fd_sc_hd__fa_1
XFILLER_129_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1733_ clknet_leaf_24_clk booth_b46_m0 VGND VGND VPWR VPWR pp_row46_23 sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_99_2 pp_row99_6 pp_row99_7 pp_row99_8 VGND VGND VPWR VPWR c$1918 s$1919
+ sky130_fd_sc_hd__fa_1
XFILLER_7_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1664_ clknet_leaf_24_clk booth_b20_m24 VGND VGND VPWR VPWR pp_row44_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_116_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_76_1 s$3147 s$3149 s$3151 VGND VGND VPWR VPWR c$3702 s$3703 sky130_fd_sc_hd__fa_2
XFILLER_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0615_ clknet_leaf_195_clk net238 VGND VGND VPWR VPWR pp_row83_24 sky130_fd_sc_hd__dfxtp_1
XFILLER_153_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1595_ clknet_leaf_5_clk booth_b34_m7 VGND VGND VPWR VPWR pp_row41_17 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_69_0 c$3098 c$3100 c$3102 VGND VGND VPWR VPWR c$3672 s$3673 sky130_fd_sc_hd__fa_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout707 sel_1$6578 VGND VGND VPWR VPWR net707 sky130_fd_sc_hd__buf_4
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0546_ clknet_leaf_171_clk booth_b42_m39 VGND VGND VPWR VPWR pp_row81_13 sky130_fd_sc_hd__dfxtp_1
Xfanout718 net719 VGND VGND VPWR VPWR net718 sky130_fd_sc_hd__buf_4
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout729 net731 VGND VGND VPWR VPWR net729 sky130_fd_sc_hd__buf_4
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0477_ clknet_leaf_129_clk booth_b58_m57 VGND VGND VPWR VPWR pp_row115_4 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_68_8 s$137 s$139 s$141 VGND VGND VPWR VPWR c$688 s$689 sky130_fd_sc_hd__fa_1
XFILLER_26_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2216_ clknet_leaf_133_clk booth_b48_m62 VGND VGND VPWR VPWR pp_row110_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_67_996 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2147_ clknet_leaf_87_clk booth_b58_m1 VGND VGND VPWR VPWR pp_row59_29 sky130_fd_sc_hd__dfxtp_1
XFILLER_38_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2078_ clknet_leaf_85_clk booth_b56_m1 VGND VGND VPWR VPWR pp_row57_28 sky130_fd_sc_hd__dfxtp_1
XU$$3080 net1046 net510 net1030 net783 VGND VGND VPWR VPWR t$5979 sky130_fd_sc_hd__a22o_1
Xdadda_fa_6_8_0 c$3424 c$3426 s$3429 VGND VGND VPWR VPWR c$3912 s$3913 sky130_fd_sc_hd__fa_1
XU$$3091 t$5984 net1360 VGND VGND VPWR VPWR booth_b44_m35 sky130_fd_sc_hd__xor2_1
XFILLER_35_882 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1029_ clknet_leaf_248_clk net190 VGND VGND VPWR VPWR pp_row3_2 sky130_fd_sc_hd__dfxtp_4
Xclkbuf_leaf_127_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_127_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_50_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2390 t$5626 net1422 VGND VGND VPWR VPWR booth_b34_m27 sky130_fd_sc_hd__xor2_1
XFILLER_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_71_0 s$1589 c$2398 c$2400 VGND VGND VPWR VPWR c$3116 s$3117 sky130_fd_sc_hd__fa_1
Xdadda_fa_1_87_0 pp_row87_0 pp_row87_1 pp_row87_2 VGND VGND VPWR VPWR c$990 s$991
+ sky130_fd_sc_hd__fa_1
XFILLER_103_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$330 final_adder.p_new$332 final_adder.p_new$330 VGND VGND VPWR VPWR
+ final_adder.p_new$458 sky130_fd_sc_hd__and2_1
XTAP_4346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$341 final_adder.p_new$340 final_adder.g_new$343 final_adder.g_new$341
+ VGND VGND VPWR VPWR final_adder.g_new$469 sky130_fd_sc_hd__a21o_1
XTAP_4368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$352 final_adder.p_new$354 final_adder.p_new$352 VGND VGND VPWR VPWR
+ final_adder.p_new$480 sky130_fd_sc_hd__and2_1
XTAP_4379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$202 t$4508 net1385 VGND VGND VPWR VPWR booth_b2_m29 sky130_fd_sc_hd__xor2_1
XFILLER_57_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$363 final_adder.p_new$362 final_adder.g_new$365 final_adder.g_new$363
+ VGND VGND VPWR VPWR final_adder.g_new$491 sky130_fd_sc_hd__a21o_1
XTAP_3645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$374 final_adder.p_new$376 final_adder.p_new$374 VGND VGND VPWR VPWR
+ final_adder.p_new$502 sky130_fd_sc_hd__and2_1
XU$$213 net982 net619 net973 net892 VGND VGND VPWR VPWR t$4514 sky130_fd_sc_hd__a22o_1
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$224 t$4519 net1385 VGND VGND VPWR VPWR booth_b2_m40 sky130_fd_sc_hd__xor2_1
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$385 final_adder.p_new$386 final_adder.g_new$391 final_adder.g_new$387
+ VGND VGND VPWR VPWR final_adder.g_new$513 sky130_fd_sc_hd__a21o_1
XFILLER_17_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$396 final_adder.p_new$402 final_adder.p_new$398 VGND VGND VPWR VPWR
+ final_adder.p_new$524 sky130_fd_sc_hd__and2_1
XU$$235 net1711 net621 net1703 net894 VGND VGND VPWR VPWR t$4525 sky130_fd_sc_hd__a22o_1
XU$$246 t$4530 net1392 VGND VGND VPWR VPWR booth_b2_m51 sky130_fd_sc_hd__xor2_1
XTAP_3678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$257 net1604 net621 net1595 net894 VGND VGND VPWR VPWR t$4536 sky130_fd_sc_hd__a22o_1
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$268 t$4541 net1388 VGND VGND VPWR VPWR booth_b2_m62 sky130_fd_sc_hd__xor2_1
XFILLER_72_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$279 net45 net1388 VGND VGND VPWR VPWR sel_1$4548 sky130_fd_sc_hd__xor2_4
XTAP_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_118_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_118_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_913 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$7 t$4410 net1574 VGND VGND VPWR VPWR booth_b0_m0 sky130_fd_sc_hd__xor2_1
Xdadda_fa_6_86_0 c$3736 c$3738 s$3741 VGND VGND VPWR VPWR c$4068 s$4069 sky130_fd_sc_hd__fa_1
XFILLER_5_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0400_ clknet_leaf_127_clk booth_b62_m52 VGND VGND VPWR VPWR pp_row114_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_171_1022 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1380_ clknet_leaf_42_clk booth_b16_m16 VGND VGND VPWR VPWR pp_row32_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_110_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0331_ clknet_leaf_224_clk booth_b38_m36 VGND VGND VPWR VPWR pp_row74_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_95_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0262_ clknet_leaf_210_clk booth_b32_m40 VGND VGND VPWR VPWR pp_row72_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_64_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2001_ clknet_leaf_62_clk booth_b38_m17 VGND VGND VPWR VPWR pp_row55_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_36_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0193_ clknet_leaf_146_clk booth_b28_m42 VGND VGND VPWR VPWR pp_row70_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_75_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_109_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_109_clk
+ sky130_fd_sc_hd__clkbuf_16
XU$$780 t$4803 net1416 VGND VGND VPWR VPWR booth_b10_m44 sky130_fd_sc_hd__xor2_1
XU$$791 net1681 net408 net1656 net674 VGND VGND VPWR VPWR t$4809 sky130_fd_sc_hd__a22o_1
XFILLER_56_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1716_ clknet_leaf_138_clk booth_b54_m52 VGND VGND VPWR VPWR pp_row106_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_172_551 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1647_ clknet_leaf_5_clk booth_b36_m7 VGND VGND VPWR VPWR pp_row43_18 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_80_7 pp_row80_21 pp_row80_22 pp_row80_23 VGND VGND VPWR VPWR c$902 s$903
+ sky130_fd_sc_hd__fa_1
XFILLER_99_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout504 net509 VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__clkbuf_4
Xfanout515 net516 VGND VGND VPWR VPWR net515 sky130_fd_sc_hd__buf_4
XFILLER_113_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1578_ clknet_leaf_243_clk booth_b4_m37 VGND VGND VPWR VPWR pp_row41_2 sky130_fd_sc_hd__dfxtp_1
Xfanout526 sel_0$5877 VGND VGND VPWR VPWR net526 sky130_fd_sc_hd__clkbuf_8
Xdadda_fa_1_73_6 pp_row73_27 pp_row73_28 pp_row73_29 VGND VGND VPWR VPWR c$774 s$775
+ sky130_fd_sc_hd__fa_1
XFILLER_98_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout537 net538 VGND VGND VPWR VPWR net537 sky130_fd_sc_hd__clkbuf_8
Xfanout548 net550 VGND VGND VPWR VPWR net548 sky130_fd_sc_hd__buf_4
XFILLER_58_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout559 sel_0$5667 VGND VGND VPWR VPWR net559 sky130_fd_sc_hd__buf_6
X_0529_ clknet_leaf_159_clk booth_b64_m16 VGND VGND VPWR VPWR pp_row80_25 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_66_5 pp_row66_33 c$96 c$98 VGND VGND VPWR VPWR c$646 s$647 sky130_fd_sc_hd__fa_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_59_4 pp_row59_23 pp_row59_24 pp_row59_25 VGND VGND VPWR VPWR c$518 s$519
+ sky130_fd_sc_hd__fa_1
XFILLER_27_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_29_2 s$2073 s$2075 s$2077 VGND VGND VPWR VPWR c$2868 s$2869 sky130_fd_sc_hd__fa_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_835 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4506 net1601 sel_0$6647 net1592 net696 VGND VGND VPWR VPWR t$6707 sky130_fd_sc_hd__a22o_1
XU$$4517 t$6712 net1879 VGND VGND VPWR VPWR booth_b64_m63 sky130_fd_sc_hd__xor2_1
XTAP_4121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_579 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3805 net1686 net474 net1661 net747 VGND VGND VPWR VPWR t$6349 sky130_fd_sc_hd__a22o_1
XFILLER_92_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_ha_3_18_2 pp_row18_6 pp_row18_7 VGND VGND VPWR VPWR c$1990 s$1991 sky130_fd_sc_hd__ha_1
XFILLER_92_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3816 t$6354 net1306 VGND VGND VPWR VPWR booth_b54_m55 sky130_fd_sc_hd__xor2_1
XU$$3827 net1554 net469 net1545 net742 VGND VGND VPWR VPWR t$6360 sky130_fd_sc_hd__a22o_1
XTAP_4176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$160 final_adder.$signal$1184 final_adder.$signal$1185 VGND VGND VPWR
+ VPWR final_adder.p_new$288 sky130_fd_sc_hd__and2_1
XTAP_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_944 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3838 net1292 VGND VGND VPWR VPWR notblock$6365\[2\] sky130_fd_sc_hd__inv_1
XTAP_4187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3849 t$6372 net1291 VGND VGND VPWR VPWR booth_b56_m3 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$171 final_adder.$signal$1175 final_adder.$signal$170 final_adder.$signal$172
+ VGND VGND VPWR VPWR final_adder.g_new$299 sky130_fd_sc_hd__a21o_1
XTAP_4198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_31_2 c$1096 c$1098 s$1101 VGND VGND VPWR VPWR c$2090 s$2091 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$182 final_adder.$signal$1162 final_adder.$signal$1163 VGND VGND VPWR
+ VPWR final_adder.p_new$310 sky130_fd_sc_hd__and2_1
XTAP_3464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$193 final_adder.$signal$1153 final_adder.$signal$126 final_adder.$signal$128
+ VGND VGND VPWR VPWR final_adder.g_new$321 sky130_fd_sc_hd__a21o_1
XFILLER_166_1113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_420 net511 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_24_1 pp_row24_8 pp_row24_9 pp_row24_10 VGND VGND VPWR VPWR c$2032 s$2033
+ sky130_fd_sc_hd__fa_1
XANTENNA_431 net713 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_442 net986 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_453 net1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_464 net1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_17_0 pp_row17_0 pp_row17_1 pp_row17_2 VGND VGND VPWR VPWR c$1982 s$1983
+ sky130_fd_sc_hd__fa_1
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0880_ clknet_leaf_194_clk net250 VGND VGND VPWR VPWR pp_row94_19 sky130_fd_sc_hd__dfxtp_2
XFILLER_9_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1501_ clknet_leaf_244_clk net187 VGND VGND VPWR VPWR pp_row37_19 sky130_fd_sc_hd__dfxtp_2
XFILLER_5_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2481_ clknet_leaf_147_clk notsign$4614 VGND VGND VPWR VPWR pp_row69_0 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_83_5 s$945 s$947 s$949 VGND VGND VPWR VPWR c$1732 s$1733 sky130_fd_sc_hd__fa_1
X_1432_ clknet_leaf_63_clk booth_b32_m2 VGND VGND VPWR VPWR pp_row34_16 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_76_4 s$821 s$823 s$825 VGND VGND VPWR VPWR c$1646 s$1647 sky130_fd_sc_hd__fa_1
XFILLER_96_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1363_ clknet_leaf_9_clk booth_b18_m13 VGND VGND VPWR VPWR pp_row31_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_95_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_69_3 c$688 s$691 s$693 VGND VGND VPWR VPWR c$1560 s$1561 sky130_fd_sc_hd__fa_1
XFILLER_110_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0314_ clknet_leaf_200_clk booth_b64_m9 VGND VGND VPWR VPWR pp_row73_28 sky130_fd_sc_hd__dfxtp_1
X_1294_ clknet_leaf_119_clk booth_b60_m43 VGND VGND VPWR VPWR pp_row103_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_39_1 s$2925 s$2927 s$2929 VGND VGND VPWR VPWR c$3554 s$3555 sky130_fd_sc_hd__fa_2
XFILLER_23_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0245_ clknet_leaf_145_clk booth_b60_m11 VGND VGND VPWR VPWR pp_row71_27 sky130_fd_sc_hd__dfxtp_1
XFILLER_48_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0176_ clknet_leaf_99_clk booth_b60_m9 VGND VGND VPWR VPWR pp_row69_28 sky130_fd_sc_hd__dfxtp_1
XFILLER_110_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_1074 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_113_1 s$3369 s$3371 s$3373 VGND VGND VPWR VPWR c$3850 s$3851 sky130_fd_sc_hd__fa_1
XFILLER_176_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_106_0 c$3320 c$3322 c$3324 VGND VGND VPWR VPWR c$3820 s$3821 sky130_fd_sc_hd__fa_1
XFILLER_191_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4415_1828 VGND VGND VPWR VPWR U$$4415_1828/HI net1828 sky130_fd_sc_hd__conb_1
Xdadda_fa_1_71_3 pp_row71_21 pp_row71_22 pp_row71_23 VGND VGND VPWR VPWR c$732 s$733
+ sky130_fd_sc_hd__fa_1
XFILLER_8_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_64_2 pp_row64_24 pp_row64_25 pp_row64_26 VGND VGND VPWR VPWR c$604 s$605
+ sky130_fd_sc_hd__fa_1
XFILLER_115_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout389 net392 VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_4_41_1 c$2162 c$2164 s$2167 VGND VGND VPWR VPWR c$2938 s$2939 sky130_fd_sc_hd__fa_1
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1078 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_57_1 pp_row57_11 pp_row57_12 pp_row57_13 VGND VGND VPWR VPWR c$476 s$477
+ sky130_fd_sc_hd__fa_1
XFILLER_189_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_34_0 s$1145 c$2102 c$2104 VGND VGND VPWR VPWR c$2894 s$2895 sky130_fd_sc_hd__fa_1
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_86_3 s$1763 s$1765 s$1767 VGND VGND VPWR VPWR c$2532 s$2533 sky130_fd_sc_hd__fa_1
XFILLER_184_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_79_2 c$1672 s$1675 s$1677 VGND VGND VPWR VPWR c$2474 s$2475 sky130_fd_sc_hd__fa_1
XFILLER_104_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_49_0 c$3588 c$3590 s$3593 VGND VGND VPWR VPWR c$3994 s$3995 sky130_fd_sc_hd__fa_1
XU$$4303 net1085 net420 net1077 net702 VGND VGND VPWR VPWR t$6604 sky130_fd_sc_hd__a22o_1
XU$$4314 t$6609 net1259 VGND VGND VPWR VPWR booth_b62_m30 sky130_fd_sc_hd__xor2_1
XU$$4325 net980 net424 net971 net706 VGND VGND VPWR VPWR t$6615 sky130_fd_sc_hd__a22o_1
XU$$4336 t$6620 net1261 VGND VGND VPWR VPWR booth_b62_m41 sky130_fd_sc_hd__xor2_1
Xfanout890 net891 VGND VGND VPWR VPWR net890 sky130_fd_sc_hd__clkbuf_4
XU$$3602 net1163 net480 net1153 net753 VGND VGND VPWR VPWR t$6246 sky130_fd_sc_hd__a22o_1
XU$$4347 net1710 net423 net1702 net705 VGND VGND VPWR VPWR t$6626 sky130_fd_sc_hd__a22o_1
XU$$3613 t$6251 net1319 VGND VGND VPWR VPWR booth_b52_m22 sky130_fd_sc_hd__xor2_1
XU$$4358 t$6631 net1260 VGND VGND VPWR VPWR booth_b62_m52 sky130_fd_sc_hd__xor2_1
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3624 net1060 net477 net1051 net750 VGND VGND VPWR VPWR t$6257 sky130_fd_sc_hd__a22o_1
XFILLER_46_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4369 net1598 net420 net1589 net702 VGND VGND VPWR VPWR t$6637 sky130_fd_sc_hd__a22o_1
XU$$3635 t$6262 net1323 VGND VGND VPWR VPWR booth_b52_m33 sky130_fd_sc_hd__xor2_1
XU$$2901 net1509 net523 net1500 net796 VGND VGND VPWR VPWR t$5888 sky130_fd_sc_hd__a22o_1
XU$$3646 net953 net480 net945 net753 VGND VGND VPWR VPWR t$6268 sky130_fd_sc_hd__a22o_1
XTAP_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2912 t$5893 net1372 VGND VGND VPWR VPWR booth_b42_m14 sky130_fd_sc_hd__xor2_1
XU$$3657 t$6273 net1326 VGND VGND VPWR VPWR booth_b52_m44 sky130_fd_sc_hd__xor2_1
XFILLER_46_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3668 net1686 net482 net1661 net755 VGND VGND VPWR VPWR t$6279 sky130_fd_sc_hd__a22o_1
XU$$2923 net1136 net520 net1120 net793 VGND VGND VPWR VPWR t$5899 sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_108_2 s$2705 s$2707 s$2709 VGND VGND VPWR VPWR c$3342 s$3343 sky130_fd_sc_hd__fa_1
XTAP_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2934 t$5904 net1375 VGND VGND VPWR VPWR booth_b42_m25 sky130_fd_sc_hd__xor2_1
XFILLER_34_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3679 t$6284 net1322 VGND VGND VPWR VPWR booth_b52_m55 sky130_fd_sc_hd__xor2_1
XTAP_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2945 net1024 net519 net1016 net792 VGND VGND VPWR VPWR t$5910 sky130_fd_sc_hd__a22o_1
XTAP_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2956 t$5915 net1370 VGND VGND VPWR VPWR booth_b42_m36 sky130_fd_sc_hd__xor2_1
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2967 net1747 net521 net1739 net794 VGND VGND VPWR VPWR t$5921 sky130_fd_sc_hd__a22o_1
XANTENNA_250 net1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_261 net1674 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2978 t$5926 net1371 VGND VGND VPWR VPWR booth_b42_m47 sky130_fd_sc_hd__xor2_1
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2989 net1642 net523 net1637 net796 VGND VGND VPWR VPWR t$5932 sky130_fd_sc_hd__a22o_1
XFILLER_60_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_272 net1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_283 pp_row46_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_294 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1981_ clknet_leaf_78_clk booth_b2_m53 VGND VGND VPWR VPWR pp_row55_1 sky130_fd_sc_hd__dfxtp_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0932_ clknet_leaf_130_clk notsign$6434 VGND VGND VPWR VPWR pp_row121_0 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_40_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_140_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0863_ clknet_leaf_105_clk booth_b36_m58 VGND VGND VPWR VPWR pp_row94_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_158_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0794_ clknet_leaf_93_clk booth_b30_m61 VGND VGND VPWR VPWR pp_row91_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_177_1050 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1083 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_81_2 c$896 c$898 c$900 VGND VGND VPWR VPWR c$1702 s$1703 sky130_fd_sc_hd__fa_1
XFILLER_103_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2464_ clknet_leaf_94_clk booth_b38_m30 VGND VGND VPWR VPWR pp_row68_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_138_1067 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_74_1 c$766 c$768 c$770 VGND VGND VPWR VPWR c$1616 s$1617 sky130_fd_sc_hd__fa_1
X_1415_ clknet_leaf_40_clk booth_b2_m32 VGND VGND VPWR VPWR pp_row34_1 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_51_0 c$2990 c$2992 c$2994 VGND VGND VPWR VPWR c$3600 s$3601 sky130_fd_sc_hd__fa_1
X_2395_ clknet_leaf_96_clk booth_b44_m22 VGND VGND VPWR VPWR pp_row66_22 sky130_fd_sc_hd__dfxtp_1
XFILLER_60_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_67_0 s$131 c$636 c$638 VGND VGND VPWR VPWR c$1530 s$1531 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$907 final_adder.$signal$1198 final_adder.g_new$983 final_adder.$signal$218
+ VGND VGND VPWR VPWR final_adder.g_new$1035 sky130_fd_sc_hd__a21o_1
X_1346_ clknet_leaf_3_clk booth_b24_m6 VGND VGND VPWR VPWR pp_row30_12 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$918 final_adder.$signal$1176 final_adder.g_new$1005 final_adder.$signal$174
+ VGND VGND VPWR VPWR final_adder.g_new$1046 sky130_fd_sc_hd__a21o_1
XFILLER_84_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_985 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$929 final_adder.$signal$1154 final_adder.g_new$931 final_adder.$signal$130
+ VGND VGND VPWR VPWR final_adder.g_new$1057 sky130_fd_sc_hd__a21o_1
XFILLER_68_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1277_ clknet_leaf_9_clk net1458 VGND VGND VPWR VPWR pp_row26_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_84_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0228_ clknet_leaf_153_clk booth_b30_m41 VGND VGND VPWR VPWR pp_row71_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_51_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_31_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_138_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_96_2 s$2609 s$2611 s$2613 VGND VGND VPWR VPWR c$3270 s$3271 sky130_fd_sc_hd__fa_1
XFILLER_193_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_89_1 c$2546 c$2548 s$2551 VGND VGND VPWR VPWR c$3226 s$3227 sky130_fd_sc_hd__fa_1
XFILLER_133_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_66_0 s$3663 c$4026 s$4029 VGND VGND VPWR VPWR c$4284 s$4285 sky130_fd_sc_hd__fa_1
XFILLER_105_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1107 net1110 VGND VGND VPWR VPWR net1107 sky130_fd_sc_hd__clkbuf_8
Xfanout1118 net77 VGND VGND VPWR VPWR net1118 sky130_fd_sc_hd__buf_4
XFILLER_120_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_98_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_98_clk sky130_fd_sc_hd__clkbuf_16
Xfanout1129 net76 VGND VGND VPWR VPWR net1129 sky130_fd_sc_hd__buf_4
XU$$2208 net1676 net571 net1561 net844 VGND VGND VPWR VPWR t$5534 sky130_fd_sc_hd__a22o_1
XU$$2219 t$5539 net1430 VGND VGND VPWR VPWR booth_b32_m10 sky130_fd_sc_hd__xor2_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1507 net1491 VGND VGND VPWR VPWR notblock$5175\[0\] sky130_fd_sc_hd__inv_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1518 t$5181 net1475 VGND VGND VPWR VPWR booth_b22_m2 sky130_fd_sc_hd__xor2_1
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1529 net1511 net610 net1503 net883 VGND VGND VPWR VPWR t$5187 sky130_fd_sc_hd__a22o_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_22_clk clknet_5_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_184_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_91_1 c$1810 c$1812 c$1814 VGND VGND VPWR VPWR c$2568 s$2569 sky130_fd_sc_hd__fa_1
XFILLER_6_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_84_0 s$965 c$1722 c$1724 VGND VGND VPWR VPWR c$2510 s$2511 sky130_fd_sc_hd__fa_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_89_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_89_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_78_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1630 net1632 VGND VGND VPWR VPWR net1630 sky130_fd_sc_hd__buf_4
X_1200_ clknet_leaf_49_clk booth_b0_m22 VGND VGND VPWR VPWR pp_row22_0 sky130_fd_sc_hd__dfxtp_1
X_2180_ clknet_leaf_218_clk booth_b54_m6 VGND VGND VPWR VPWR pp_row60_27 sky130_fd_sc_hd__dfxtp_1
XFILLER_78_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1641 net112 VGND VGND VPWR VPWR net1641 sky130_fd_sc_hd__buf_4
Xfanout1652 net1653 VGND VGND VPWR VPWR net1652 sky130_fd_sc_hd__buf_4
XU$$4100 t$6499 net1284 VGND VGND VPWR VPWR booth_b58_m60 sky130_fd_sc_hd__xor2_1
Xfanout1663 net1667 VGND VGND VPWR VPWR net1663 sky130_fd_sc_hd__buf_6
XFILLER_66_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4111 net57 VGND VGND VPWR VPWR notblock$6505\[1\] sky130_fd_sc_hd__inv_1
XU$$4122 net87 net434 net98 net716 VGND VGND VPWR VPWR t$6512 sky130_fd_sc_hd__a22o_1
Xfanout1674 net109 VGND VGND VPWR VPWR net1674 sky130_fd_sc_hd__buf_4
XU$$4133 t$6517 net1269 VGND VGND VPWR VPWR booth_b60_m8 sky130_fd_sc_hd__xor2_1
Xfanout1685 net108 VGND VGND VPWR VPWR net1685 sky130_fd_sc_hd__buf_4
X_1131_ clknet_leaf_11_clk booth_b14_m2 VGND VGND VPWR VPWR pp_row16_7 sky130_fd_sc_hd__dfxtp_1
XU$$4144 net1196 net434 net1177 net716 VGND VGND VPWR VPWR t$6523 sky130_fd_sc_hd__a22o_1
Xfanout1696 net1697 VGND VGND VPWR VPWR net1696 sky130_fd_sc_hd__buf_4
XU$$4155 t$6528 net1267 VGND VGND VPWR VPWR booth_b60_m19 sky130_fd_sc_hd__xor2_1
XU$$3410 net1600 net499 net1591 net772 VGND VGND VPWR VPWR t$6147 sky130_fd_sc_hd__a22o_1
XU$$4166 net1085 net436 net1077 net718 VGND VGND VPWR VPWR t$6534 sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_46_5 s$295 s$297 s$299 VGND VGND VPWR VPWR c$1288 s$1289 sky130_fd_sc_hd__fa_1
Xdadda_fa_4_113_0 pp_row113_6 pp_row113_7 pp_row113_8 VGND VGND VPWR VPWR c$3368 s$3369
+ sky130_fd_sc_hd__fa_1
XU$$3421 t$6152 net1345 VGND VGND VPWR VPWR booth_b48_m63 sky130_fd_sc_hd__xor2_1
XFILLER_168_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3432 t$6159 net1329 VGND VGND VPWR VPWR booth_b50_m0 sky130_fd_sc_hd__xor2_1
XU$$4177 t$6539 net1270 VGND VGND VPWR VPWR booth_b60_m30 sky130_fd_sc_hd__xor2_1
XU$$4188 net979 net438 net970 net720 VGND VGND VPWR VPWR t$6545 sky130_fd_sc_hd__a22o_1
X_1062_ clknet_leaf_51_clk booth_b2_m7 VGND VGND VPWR VPWR pp_row9_1 sky130_fd_sc_hd__dfxtp_1
XU$$3443 net1566 net492 net1525 net765 VGND VGND VPWR VPWR t$6165 sky130_fd_sc_hd__a22o_1
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4199 t$6550 net1271 VGND VGND VPWR VPWR booth_b60_m41 sky130_fd_sc_hd__xor2_1
XU$$3454 t$6170 net1329 VGND VGND VPWR VPWR booth_b50_m11 sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_39_4 pp_row39_20 c$216 c$218 VGND VGND VPWR VPWR c$1202 s$1203 sky130_fd_sc_hd__fa_1
XU$$3465 net1163 net488 net1153 net761 VGND VGND VPWR VPWR t$6176 sky130_fd_sc_hd__a22o_1
XU$$2720 t$5794 net1400 VGND VGND VPWR VPWR booth_b38_m55 sky130_fd_sc_hd__xor2_1
XFILLER_20_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2731 net1557 net548 net1550 net821 VGND VGND VPWR VPWR t$5800 sky130_fd_sc_hd__a22o_1
XU$$3476 t$6181 net1329 VGND VGND VPWR VPWR booth_b50_m22 sky130_fd_sc_hd__xor2_1
XU$$3487 net1060 net485 net1051 net758 VGND VGND VPWR VPWR t$6187 sky130_fd_sc_hd__a22o_1
XU$$2742 net1378 VGND VGND VPWR VPWR notblock$5805\[2\] sky130_fd_sc_hd__inv_1
XTAP_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2753 t$5812 net1376 VGND VGND VPWR VPWR booth_b40_m3 sky130_fd_sc_hd__xor2_1
XU$$3498 t$6192 net1331 VGND VGND VPWR VPWR booth_b50_m33 sky130_fd_sc_hd__xor2_1
XTAP_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2764 net1506 net536 net1497 net809 VGND VGND VPWR VPWR t$5818 sky130_fd_sc_hd__a22o_1
XU$$2775 t$5823 net1381 VGND VGND VPWR VPWR booth_b40_m14 sky130_fd_sc_hd__xor2_1
XU$$2786 net1132 net535 net1116 net808 VGND VGND VPWR VPWR t$5829 sky130_fd_sc_hd__a22o_1
XU$$2797 t$5834 net1381 VGND VGND VPWR VPWR booth_b40_m25 sky130_fd_sc_hd__xor2_1
XFILLER_33_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1964_ clknet_leaf_63_clk booth_b30_m24 VGND VGND VPWR VPWR pp_row54_15 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_13_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_119_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0915_ clknet_leaf_104_clk booth_b56_m40 VGND VGND VPWR VPWR pp_row96_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_174_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1895_ clknet_leaf_65_clk booth_b20_m32 VGND VGND VPWR VPWR pp_row52_10 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_99_0 c$3278 c$3280 c$3282 VGND VGND VPWR VPWR c$3792 s$3793 sky130_fd_sc_hd__fa_1
XFILLER_179_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0846_ clknet_leaf_105_clk booth_b42_m51 VGND VGND VPWR VPWR pp_row93_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_134_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0777_ clknet_leaf_181_clk net149 VGND VGND VPWR VPWR pp_row118_7 sky130_fd_sc_hd__dfxtp_2
XFILLER_143_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2447_ clknet_leaf_128_clk booth_b48_m64 VGND VGND VPWR VPWR pp_row112_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_69_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$704 final_adder.p_new$728 final_adder.p_new$712 VGND VGND VPWR VPWR
+ final_adder.p_new$832 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$715 final_adder.p_new$722 final_adder.g_new$739 final_adder.g_new$723
+ VGND VGND VPWR VPWR final_adder.g_new$843 sky130_fd_sc_hd__a21o_1
XFILLER_69_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2378_ clknet_leaf_83_clk booth_b16_m50 VGND VGND VPWR VPWR pp_row66_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_96_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$737 final_adder.p_new$744 final_adder.g_new$383 final_adder.g_new$745
+ VGND VGND VPWR VPWR final_adder.g_new$865 sky130_fd_sc_hd__a21o_2
XFILLER_29_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$748 final_adder.p_new$796 final_adder.p_new$764 VGND VGND VPWR VPWR
+ final_adder.p_new$876 sky130_fd_sc_hd__and2_1
X_1329_ clknet_leaf_4_clk booth_b24_m5 VGND VGND VPWR VPWR pp_row29_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_112_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$759 final_adder.p_new$774 final_adder.g_new$807 final_adder.g_new$775
+ VGND VGND VPWR VPWR final_adder.g_new$887 sky130_fd_sc_hd__a21o_1
XFILLER_186_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$609 t$4716 net1239 VGND VGND VPWR VPWR booth_b8_m27 sky130_fd_sc_hd__xor2_1
XFILLER_83_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_108_1 pp_row108_5 pp_row108_6 pp_row108_7 VGND VGND VPWR VPWR c$2704 s$2705
+ sky130_fd_sc_hd__fa_1
XFILLER_133_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput290 net290 VGND VGND VPWR VPWR o[14] sky130_fd_sc_hd__buf_2
XFILLER_181_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_49_3 s$1319 s$1321 s$1323 VGND VGND VPWR VPWR c$2236 s$2237 sky130_fd_sc_hd__fa_1
XU$$4467_1854 VGND VGND VPWR VPWR U$$4467_1854/HI net1854 sky130_fd_sc_hd__conb_1
XFILLER_90_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2005 t$5429 net1455 VGND VGND VPWR VPWR booth_b28_m40 sky130_fd_sc_hd__xor2_1
XU$$2016 net1711 net586 net1703 net859 VGND VGND VPWR VPWR t$5435 sky130_fd_sc_hd__a22o_1
XU$$2027 t$5440 net1454 VGND VGND VPWR VPWR booth_b28_m51 sky130_fd_sc_hd__xor2_1
XU$$2038 net1605 net590 net1597 net863 VGND VGND VPWR VPWR t$5446 sky130_fd_sc_hd__a22o_1
XU$$1304 t$5071 net1666 VGND VGND VPWR VPWR booth_b18_m32 sky130_fd_sc_hd__xor2_1
XU$$2049 t$5451 net1456 VGND VGND VPWR VPWR booth_b28_m62 sky130_fd_sc_hd__xor2_1
XFILLER_16_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1315 net957 net638 net949 net911 VGND VGND VPWR VPWR t$5077 sky130_fd_sc_hd__a22o_1
XFILLER_188_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1326 t$5082 net1663 VGND VGND VPWR VPWR booth_b18_m43 sky130_fd_sc_hd__xor2_1
XU$$1337 net1692 net642 net1680 net915 VGND VGND VPWR VPWR t$5088 sky130_fd_sc_hd__a22o_1
XU$$1348 t$5093 net1669 VGND VGND VPWR VPWR booth_b18_m54 sky130_fd_sc_hd__xor2_1
XFILLER_71_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1359 net1581 net641 net1552 net914 VGND VGND VPWR VPWR t$5099 sky130_fd_sc_hd__a22o_1
XFILLER_71_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_903 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0700_ clknet_leaf_174_clk booth_b32_m55 VGND VGND VPWR VPWR pp_row87_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_156_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1680_ clknet_leaf_24_clk booth_b0_m45 VGND VGND VPWR VPWR pp_row45_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_183_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0631_ clknet_leaf_178_clk booth_b48_m36 VGND VGND VPWR VPWR pp_row84_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0562_ clknet_leaf_186_clk booth_b22_m60 VGND VGND VPWR VPWR pp_row82_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_140_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2301_ clknet_leaf_198_clk booth_b8_m56 VGND VGND VPWR VPWR pp_row64_4 sky130_fd_sc_hd__dfxtp_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0493_ clknet_leaf_161_clk booth_b52_m27 VGND VGND VPWR VPWR pp_row79_19 sky130_fd_sc_hd__dfxtp_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2232_ clknet_leaf_233_clk booth_b18_m44 VGND VGND VPWR VPWR pp_row62_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_2_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_2_51_3 c$364 s$367 s$369 VGND VGND VPWR VPWR c$1344 s$1345 sky130_fd_sc_hd__fa_1
Xfanout1460 net1462 VGND VGND VPWR VPWR net1460 sky130_fd_sc_hd__buf_6
Xfanout1471 net1472 VGND VGND VPWR VPWR net1471 sky130_fd_sc_hd__buf_4
XFILLER_78_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1482 net1483 VGND VGND VPWR VPWR net1482 sky130_fd_sc_hd__buf_4
X_2163_ clknet_leaf_30_clk booth_b24_m36 VGND VGND VPWR VPWR pp_row60_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_94_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1493 net14 VGND VGND VPWR VPWR net1493 sky130_fd_sc_hd__buf_8
XFILLER_39_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_44_2 pp_row44_23 pp_row44_24 c$254 VGND VGND VPWR VPWR c$1258 s$1259 sky130_fd_sc_hd__fa_1
XFILLER_66_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1114_ clknet_leaf_13_clk booth_b2_m13 VGND VGND VPWR VPWR pp_row15_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$11 c$4172 s$4175 VGND VGND VPWR VPWR final_adder.$signal$24 final_adder.$signal$1101
+ sky130_fd_sc_hd__ha_1
XU$$3240 t$6060 net1351 VGND VGND VPWR VPWR booth_b46_m41 sky130_fd_sc_hd__xor2_1
X_2094_ clknet_leaf_143_clk booth_b48_m61 VGND VGND VPWR VPWR pp_row109_2 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_21_1 s$2817 s$2819 s$2821 VGND VGND VPWR VPWR c$3482 s$3483 sky130_fd_sc_hd__fa_1
XU$$3251 net1708 net507 net1700 net780 VGND VGND VPWR VPWR t$6066 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$22 c$4194 s$4197 VGND VGND VPWR VPWR final_adder.$signal$46 final_adder.$signal$1112
+ sky130_fd_sc_hd__ha_2
XU$$3262 t$6071 net1355 VGND VGND VPWR VPWR booth_b46_m52 sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_37_1 pp_row37_8 pp_row37_9 pp_row37_10 VGND VGND VPWR VPWR c$1172 s$1173
+ sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$33 c$4216 s$4219 VGND VGND VPWR VPWR final_adder.$signal$68 final_adder.$signal$1123
+ sky130_fd_sc_hd__ha_1
XU$$3273 net1602 net507 net1593 net780 VGND VGND VPWR VPWR t$6077 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$44 c$4238 s$4241 VGND VGND VPWR VPWR final_adder.$signal$90 final_adder.$signal$1134
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$55 c$4260 s$4263 VGND VGND VPWR VPWR final_adder.$signal$112 final_adder.$signal$113
+ sky130_fd_sc_hd__ha_1
XFILLER_0_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1045_ clknet_leaf_248_clk net223 VGND VGND VPWR VPWR pp_row6_5 sky130_fd_sc_hd__dfxtp_4
XU$$3284 t$6082 net1356 VGND VGND VPWR VPWR booth_b46_m63 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$66 c$4282 s$4285 VGND VGND VPWR VPWR final_adder.$signal$134 final_adder.$signal$1156
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_5_14_0 c$2768 c$2770 c$2772 VGND VGND VPWR VPWR c$3452 s$3453 sky130_fd_sc_hd__fa_2
XU$$2550 net950 net555 net942 net828 VGND VGND VPWR VPWR t$5708 sky130_fd_sc_hd__a22o_1
XU$$3295 t$6089 net1338 VGND VGND VPWR VPWR booth_b48_m0 sky130_fd_sc_hd__xor2_1
XU$$2561 t$5713 net1409 VGND VGND VPWR VPWR booth_b36_m44 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$77 c$4304 s$4307 VGND VGND VPWR VPWR final_adder.$signal$156 final_adder.$signal$1167
+ sky130_fd_sc_hd__ha_1
XU$$2572 net1680 net556 net1655 net829 VGND VGND VPWR VPWR t$5719 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$88 c$4326 s$4329 VGND VGND VPWR VPWR final_adder.$signal$178 final_adder.$signal$1178
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$99 c$4348 s$4351 VGND VGND VPWR VPWR final_adder.$signal$200 final_adder.$signal$1189
+ sky130_fd_sc_hd__ha_1
XFILLER_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2583 t$5724 net1410 VGND VGND VPWR VPWR booth_b36_m55 sky130_fd_sc_hd__xor2_1
XFILLER_146_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2594 net1557 net558 net1550 net831 VGND VGND VPWR VPWR t$5730 sky130_fd_sc_hd__a22o_1
XU$$1860 t$5355 net1459 VGND VGND VPWR VPWR booth_b26_m36 sky130_fd_sc_hd__xor2_1
XFILLER_107_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1871 net1747 net600 net1739 net873 VGND VGND VPWR VPWR t$5361 sky130_fd_sc_hd__a22o_1
XU$$1882 t$5366 net1464 VGND VGND VPWR VPWR booth_b26_m47 sky130_fd_sc_hd__xor2_1
XU$$1893 net1639 net598 net1631 net871 VGND VGND VPWR VPWR t$5372 sky130_fd_sc_hd__a22o_1
XFILLER_9_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1947_ clknet_leaf_78_clk booth_b2_m52 VGND VGND VPWR VPWR pp_row54_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_159_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1878_ clknet_leaf_70_clk booth_b44_m7 VGND VGND VPWR VPWR pp_row51_22 sky130_fd_sc_hd__dfxtp_1
XFILLER_174_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0829_ clknet_leaf_108_clk booth_b54_m38 VGND VGND VPWR VPWR pp_row92_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_1_40_3 pp_row40_9 pp_row40_10 VGND VGND VPWR VPWR c$234 s$235 sky130_fd_sc_hd__ha_1
Xdadda_fa_4_59_2 s$2313 s$2315 s$2317 VGND VGND VPWR VPWR c$3048 s$3049 sky130_fd_sc_hd__fa_1
XFILLER_130_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$501 final_adder.p_new$502 final_adder.g_new$507 final_adder.g_new$503
+ VGND VGND VPWR VPWR final_adder.g_new$629 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$512 final_adder.p_new$524 final_adder.p_new$516 VGND VGND VPWR VPWR
+ final_adder.p_new$640 sky130_fd_sc_hd__and2_1
XFILLER_28_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$523 final_adder.p_new$526 final_adder.g_new$535 final_adder.g_new$527
+ VGND VGND VPWR VPWR final_adder.g_new$651 sky130_fd_sc_hd__a21o_1
XTAP_3805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_4_10_1 pp_row10_3 pp_row10_4 VGND VGND VPWR VPWR c$2756 s$2757 sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$534 final_adder.p_new$546 final_adder.p_new$538 VGND VGND VPWR VPWR
+ final_adder.p_new$662 sky130_fd_sc_hd__and2_1
XTAP_3816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$545 final_adder.p_new$548 final_adder.g_new$557 final_adder.g_new$549
+ VGND VGND VPWR VPWR final_adder.g_new$673 sky130_fd_sc_hd__a21o_1
XTAP_3827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_29_0 s$3515 c$3952 s$3955 VGND VGND VPWR VPWR c$4210 s$4211 sky130_fd_sc_hd__fa_2
XFILLER_84_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$556 final_adder.p_new$568 final_adder.p_new$560 VGND VGND VPWR VPWR
+ final_adder.p_new$684 sky130_fd_sc_hd__and2_1
XTAP_3838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$406 net1539 net534 net1531 net807 VGND VGND VPWR VPWR t$4612 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$567 final_adder.p_new$570 final_adder.g_new$579 final_adder.g_new$571
+ VGND VGND VPWR VPWR final_adder.g_new$695 sky130_fd_sc_hd__a21o_1
XTAP_3849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$417 net1806 net429 net1231 net711 VGND VGND VPWR VPWR t$4619 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$578 final_adder.p_new$590 final_adder.p_new$582 VGND VGND VPWR VPWR
+ final_adder.p_new$706 sky130_fd_sc_hd__and2_1
XFILLER_151_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$428 t$4624 net1248 VGND VGND VPWR VPWR booth_b6_m5 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$589 final_adder.p_new$592 final_adder.g_new$601 final_adder.g_new$593
+ VGND VGND VPWR VPWR final_adder.g_new$717 sky130_fd_sc_hd__a21o_1
XFILLER_56_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$439 net1221 net427 net1211 net709 VGND VGND VPWR VPWR t$4630 sky130_fd_sc_hd__a22o_1
XFILLER_25_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4497_1869 VGND VGND VPWR VPWR U$$4497_1869/HI net1869 sky130_fd_sc_hd__conb_1
XFILLER_138_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_61_2 c$1456 s$1459 s$1461 VGND VGND VPWR VPWR c$2330 s$2331 sky130_fd_sc_hd__fa_1
XFILLER_121_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_54_1 c$1366 c$1368 c$1370 VGND VGND VPWR VPWR c$2272 s$2273 sky130_fd_sc_hd__fa_1
XFILLER_0_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_31_0 c$3516 c$3518 s$3521 VGND VGND VPWR VPWR c$3958 s$3959 sky130_fd_sc_hd__fa_1
Xdadda_fa_3_47_0 s$315 c$1278 c$1280 VGND VGND VPWR VPWR c$2214 s$2215 sky130_fd_sc_hd__fa_1
XFILLER_85_74 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_997 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$940 net1615 net399 net1607 net665 VGND VGND VPWR VPWR t$4885 sky130_fd_sc_hd__a22o_1
XU$$951 t$4890 net1316 VGND VGND VPWR VPWR booth_b12_m61 sky130_fd_sc_hd__xor2_1
XU$$1101 net8 net1188 VGND VGND VPWR VPWR sel_1$4968 sky130_fd_sc_hd__xor2_4
XU$$962 net1189 notblock$4895\[1\] VGND VGND VPWR VPWR t$4896 sky130_fd_sc_hd__and2_1
XFILLER_63_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$973 net933 net387 net1672 net653 VGND VGND VPWR VPWR t$4903 sky130_fd_sc_hd__a22o_1
XU$$1112 net1676 net646 net1564 net919 VGND VGND VPWR VPWR t$4974 sky130_fd_sc_hd__a22o_1
XFILLER_189_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1123 t$4979 net1008 VGND VGND VPWR VPWR booth_b16_m10 sky130_fd_sc_hd__xor2_1
XU$$984 t$4908 net1185 VGND VGND VPWR VPWR booth_b14_m9 sky130_fd_sc_hd__xor2_1
XFILLER_188_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$995 net1173 net385 net1164 net651 VGND VGND VPWR VPWR t$4914 sky130_fd_sc_hd__a22o_1
XU$$1134 net1166 net645 net1157 net918 VGND VGND VPWR VPWR t$4985 sky130_fd_sc_hd__a22o_1
XU$$1145 t$4990 net1009 VGND VGND VPWR VPWR booth_b16_m21 sky130_fd_sc_hd__xor2_1
XU$$1156 net1064 net648 net1056 net921 VGND VGND VPWR VPWR t$4996 sky130_fd_sc_hd__a22o_1
XFILLER_189_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1167 t$5001 net1007 VGND VGND VPWR VPWR booth_b16_m32 sky130_fd_sc_hd__xor2_1
XU$$1178 net961 net645 net955 net918 VGND VGND VPWR VPWR t$5007 sky130_fd_sc_hd__a22o_1
XFILLER_188_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1189 t$5012 net1008 VGND VGND VPWR VPWR booth_b16_m43 sky130_fd_sc_hd__xor2_1
XFILLER_148_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1801_ clknet_leaf_219_clk booth_b14_m35 VGND VGND VPWR VPWR pp_row49_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_157_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_7_104_0 s$3815 c$4102 s$4105 VGND VGND VPWR VPWR c$4360 s$4361 sky130_fd_sc_hd__fa_1
XFILLER_156_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1732_ clknet_leaf_24_clk booth_b44_m2 VGND VGND VPWR VPWR pp_row46_22 sky130_fd_sc_hd__dfxtp_1
XFILLER_117_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1663_ clknet_leaf_24_clk booth_b18_m26 VGND VGND VPWR VPWR pp_row44_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_144_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_99_3 pp_row99_9 pp_row99_10 pp_row99_11 VGND VGND VPWR VPWR c$1920 s$1921
+ sky130_fd_sc_hd__fa_1
XFILLER_171_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0614_ clknet_leaf_189_clk booth_b64_m19 VGND VGND VPWR VPWR pp_row83_23 sky130_fd_sc_hd__dfxtp_1
X_1594_ clknet_leaf_110_clk booth_b58_m47 VGND VGND VPWR VPWR pp_row105_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_125_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_5_69_1 s$3105 s$3107 s$3109 VGND VGND VPWR VPWR c$3674 s$3675 sky130_fd_sc_hd__fa_1
Xfanout708 net709 VGND VGND VPWR VPWR net708 sky130_fd_sc_hd__buf_4
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0545_ clknet_leaf_167_clk booth_b40_m41 VGND VGND VPWR VPWR pp_row81_12 sky130_fd_sc_hd__dfxtp_1
Xfanout719 net723 VGND VGND VPWR VPWR net719 sky130_fd_sc_hd__buf_4
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0476_ clknet_leaf_193_clk booth_b22_m57 VGND VGND VPWR VPWR pp_row79_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_100_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1042 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2215_ clknet_leaf_29_clk booth_b52_m9 VGND VGND VPWR VPWR pp_row61_26 sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1290 net55 VGND VGND VPWR VPWR net1290 sky130_fd_sc_hd__buf_6
X_2146_ clknet_leaf_31_clk booth_b56_m3 VGND VGND VPWR VPWR pp_row59_28 sky130_fd_sc_hd__dfxtp_1
XFILLER_27_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3070 net1087 net511 net1078 net784 VGND VGND VPWR VPWR t$5974 sky130_fd_sc_hd__a22o_1
X_2077_ clknet_leaf_82_clk booth_b54_m3 VGND VGND VPWR VPWR pp_row57_27 sky130_fd_sc_hd__dfxtp_1
XU$$3081 t$5979 net1357 VGND VGND VPWR VPWR booth_b44_m30 sky130_fd_sc_hd__xor2_1
XU$$3092 net976 net513 net967 net786 VGND VGND VPWR VPWR t$5985 sky130_fd_sc_hd__a22o_1
X_1028_ clknet_leaf_61_clk booth_b2_m1 VGND VGND VPWR VPWR pp_row3_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_35_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2380 t$5621 net1424 VGND VGND VPWR VPWR booth_b34_m22 sky130_fd_sc_hd__xor2_1
XU$$2391 net1062 net565 net1053 net838 VGND VGND VPWR VPWR t$5627 sky130_fd_sc_hd__a22o_1
XFILLER_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1690 net1131 net603 net1115 net876 VGND VGND VPWR VPWR t$5269 sky130_fd_sc_hd__a22o_1
XFILLER_136_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_71_1 c$2402 c$2404 s$2407 VGND VGND VPWR VPWR c$3118 s$3119 sky130_fd_sc_hd__fa_1
Xdadda_fa_1_87_1 pp_row87_3 pp_row87_4 pp_row87_5 VGND VGND VPWR VPWR c$992 s$993
+ sky130_fd_sc_hd__fa_2
XFILLER_1_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1081 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_64_0 s$1505 c$2342 c$2344 VGND VGND VPWR VPWR c$3074 s$3075 sky130_fd_sc_hd__fa_1
XFILLER_7_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$320 final_adder.p_new$322 final_adder.p_new$320 VGND VGND VPWR VPWR
+ final_adder.p_new$448 sky130_fd_sc_hd__and2_1
XTAP_4347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$331 final_adder.p_new$330 final_adder.g_new$333 final_adder.g_new$331
+ VGND VGND VPWR VPWR final_adder.g_new$459 sky130_fd_sc_hd__a21o_1
XFILLER_57_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$342 final_adder.p_new$344 final_adder.p_new$342 VGND VGND VPWR VPWR
+ final_adder.p_new$470 sky130_fd_sc_hd__and2_1
XTAP_3624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$353 final_adder.p_new$352 final_adder.g_new$355 final_adder.g_new$353
+ VGND VGND VPWR VPWR final_adder.g_new$481 sky130_fd_sc_hd__a21o_1
XTAP_4369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$203 net1039 net620 net1024 net893 VGND VGND VPWR VPWR t$4509 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$364 final_adder.p_new$366 final_adder.p_new$364 VGND VGND VPWR VPWR
+ final_adder.p_new$492 sky130_fd_sc_hd__and2_1
XFILLER_176_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$375 final_adder.p_new$374 final_adder.g_new$377 final_adder.g_new$375
+ VGND VGND VPWR VPWR final_adder.g_new$503 sky130_fd_sc_hd__a21o_1
XU$$214 t$4514 net1385 VGND VGND VPWR VPWR booth_b2_m35 sky130_fd_sc_hd__xor2_1
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$225 net924 net621 net1745 net894 VGND VGND VPWR VPWR t$4520 sky130_fd_sc_hd__a22o_1
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$386 final_adder.p_new$392 final_adder.p_new$388 VGND VGND VPWR VPWR
+ final_adder.p_new$514 sky130_fd_sc_hd__and2_1
XTAP_3668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$397 final_adder.p_new$398 final_adder.g_new$403 final_adder.g_new$399
+ VGND VGND VPWR VPWR final_adder.g_new$525 sky130_fd_sc_hd__a21o_1
XU$$236 t$4525 net1387 VGND VGND VPWR VPWR booth_b2_m46 sky130_fd_sc_hd__xor2_1
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$247 net1650 net626 net1642 net899 VGND VGND VPWR VPWR t$4531 sky130_fd_sc_hd__a22o_1
XTAP_3679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$258 t$4536 net1387 VGND VGND VPWR VPWR booth_b2_m57 sky130_fd_sc_hd__xor2_1
XFILLER_73_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1000 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$269 net1539 net626 net1531 net899 VGND VGND VPWR VPWR t$4542 sky130_fd_sc_hd__a22o_1
XTAP_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$8 net1232 net446 net1127 net688 VGND VGND VPWR VPWR t$4411 sky130_fd_sc_hd__a22o_1
XFILLER_139_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_969 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_0_76_1 pp_row76_3 pp_row76_4 VGND VGND VPWR VPWR c$198 s$199 sky130_fd_sc_hd__ha_1
Xdadda_fa_6_79_0 c$3708 c$3710 s$3713 VGND VGND VPWR VPWR c$4054 s$4055 sky130_fd_sc_hd__fa_1
XFILLER_126_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0330_ clknet_leaf_224_clk booth_b36_m38 VGND VGND VPWR VPWR pp_row74_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_121_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0261_ clknet_leaf_210_clk booth_b30_m42 VGND VGND VPWR VPWR pp_row72_12 sky130_fd_sc_hd__dfxtp_1
X_2000_ clknet_leaf_69_clk booth_b36_m19 VGND VGND VPWR VPWR pp_row55_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_64_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0192_ clknet_leaf_148_clk booth_b26_m44 VGND VGND VPWR VPWR pp_row70_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_35_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$770 t$4798 net1418 VGND VGND VPWR VPWR booth_b10_m39 sky130_fd_sc_hd__xor2_1
XU$$781 net1724 net404 net1715 net670 VGND VGND VPWR VPWR t$4804 sky130_fd_sc_hd__a22o_1
XFILLER_189_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$792 t$4809 net1419 VGND VGND VPWR VPWR booth_b10_m50 sky130_fd_sc_hd__xor2_1
XFILLER_90_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1715_ clknet_leaf_237_clk booth_b16_m30 VGND VGND VPWR VPWR pp_row46_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_117_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_81_0 c$3170 c$3172 c$3174 VGND VGND VPWR VPWR c$3720 s$3721 sky130_fd_sc_hd__fa_1
Xdadda_fa_2_97_0 pp_row97_0 pp_row97_1 pp_row97_2 VGND VGND VPWR VPWR c$1890 s$1891
+ sky130_fd_sc_hd__fa_1
XFILLER_145_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1646_ clknet_leaf_6_clk booth_b34_m9 VGND VGND VPWR VPWR pp_row43_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_144_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout505 net506 VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__buf_4
X_1577_ clknet_leaf_243_clk booth_b2_m39 VGND VGND VPWR VPWR pp_row41_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_141_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout516 net517 VGND VGND VPWR VPWR net516 sky130_fd_sc_hd__buf_4
Xfanout527 net530 VGND VGND VPWR VPWR net527 sky130_fd_sc_hd__buf_4
XFILLER_101_803 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_73_7 c$172 c$174 c$176 VGND VGND VPWR VPWR c$776 s$777 sky130_fd_sc_hd__fa_1
Xfanout538 net542 VGND VGND VPWR VPWR net538 sky130_fd_sc_hd__buf_4
X_0528_ clknet_leaf_159_clk booth_b62_m18 VGND VGND VPWR VPWR pp_row80_24 sky130_fd_sc_hd__dfxtp_1
Xfanout549 net550 VGND VGND VPWR VPWR net549 sky130_fd_sc_hd__buf_4
XFILLER_98_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_66_6 c$100 c$102 c$104 VGND VGND VPWR VPWR c$648 s$649 sky130_fd_sc_hd__fa_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0459_ clknet_leaf_157_clk booth_b44_m34 VGND VGND VPWR VPWR pp_row78_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_55_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_59_5 pp_row59_26 pp_row59_27 pp_row59_28 VGND VGND VPWR VPWR c$520 s$521
+ sky130_fd_sc_hd__fa_1
XFILLER_55_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2129_ clknet_leaf_29_clk booth_b24_m35 VGND VGND VPWR VPWR pp_row59_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_15_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_96_0 s$3783 c$4086 s$4089 VGND VGND VPWR VPWR c$4344 s$4345 sky130_fd_sc_hd__fa_1
XFILLER_22_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4390_1815 VGND VGND VPWR VPWR U$$4390_1815/HI net1815 sky130_fd_sc_hd__conb_1
XFILLER_155_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4507 t$6707 net1874 VGND VGND VPWR VPWR booth_b64_m58 sky130_fd_sc_hd__xor2_1
XTAP_4111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_111_0 c$3836 c$3838 s$3841 VGND VGND VPWR VPWR c$4118 s$4119 sky130_fd_sc_hd__fa_1
XTAP_4144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3806 t$6349 net1308 VGND VGND VPWR VPWR booth_b54_m50 sky130_fd_sc_hd__xor2_1
XTAP_4155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3817 net1616 net473 net1608 net746 VGND VGND VPWR VPWR t$6355 sky130_fd_sc_hd__a22o_1
XTAP_4166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$150 final_adder.$signal$1194 final_adder.$signal$1195 VGND VGND VPWR
+ VPWR final_adder.p_new$278 sky130_fd_sc_hd__and2_1
XTAP_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3828 t$6360 net1302 VGND VGND VPWR VPWR booth_b54_m61 sky130_fd_sc_hd__xor2_1
XTAP_4177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$161 final_adder.$signal$1185 final_adder.$signal$190 final_adder.$signal$192
+ VGND VGND VPWR VPWR final_adder.g_new$289 sky130_fd_sc_hd__a21o_1
XTAP_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3839 net1292 notblock$6365\[1\] VGND VGND VPWR VPWR t$6366 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$172 final_adder.$signal$1172 final_adder.$signal$1173 VGND VGND VPWR
+ VPWR final_adder.p_new$300 sky130_fd_sc_hd__and2_1
XTAP_4188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_31_3 s$1103 s$1105 s$1107 VGND VGND VPWR VPWR c$2092 s$2093 sky130_fd_sc_hd__fa_1
XFILLER_46_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$183 final_adder.$signal$1163 final_adder.$signal$146 final_adder.$signal$148
+ VGND VGND VPWR VPWR final_adder.g_new$311 sky130_fd_sc_hd__a21o_1
XTAP_3465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_410 net1732 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$194 final_adder.$signal$1150 final_adder.$signal$1151 VGND VGND VPWR
+ VPWR final_adder.p_new$322 sky130_fd_sc_hd__and2_1
XFILLER_166_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_421 net526 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_24_2 pp_row24_11 pp_row24_12 pp_row24_13 VGND VGND VPWR VPWR c$2034 s$2035
+ sky130_fd_sc_hd__fa_1
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_432 net745 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_443 net1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_454 net1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_917 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1500_ clknet_leaf_45_clk booth_b36_m1 VGND VGND VPWR VPWR pp_row37_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_126_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2480_ clknet_leaf_125_clk booth_b54_m58 VGND VGND VPWR VPWR pp_row112_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_181_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1431_ clknet_leaf_63_clk booth_b30_m4 VGND VGND VPWR VPWR pp_row34_15 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_76_5 s$827 s$829 s$831 VGND VGND VPWR VPWR c$1648 s$1649 sky130_fd_sc_hd__fa_1
XFILLER_96_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1362_ clknet_leaf_10_clk booth_b16_m15 VGND VGND VPWR VPWR pp_row31_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_122_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_69_4 s$695 s$697 s$699 VGND VGND VPWR VPWR c$1562 s$1563 sky130_fd_sc_hd__fa_2
X_0313_ clknet_leaf_201_clk booth_b62_m11 VGND VGND VPWR VPWR pp_row73_27 sky130_fd_sc_hd__dfxtp_1
XFILLER_96_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1293_ clknet_leaf_3_clk booth_b24_m3 VGND VGND VPWR VPWR pp_row27_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_55_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0244_ clknet_leaf_126_clk booth_b52_m61 VGND VGND VPWR VPWR pp_row113_2 sky130_fd_sc_hd__dfxtp_1
Xinput190 c[3] VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0175_ clknet_leaf_99_clk booth_b58_m11 VGND VGND VPWR VPWR pp_row69_27 sky130_fd_sc_hd__dfxtp_1
XFILLER_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_106_1 s$3327 s$3329 s$3331 VGND VGND VPWR VPWR c$3822 s$3823 sky130_fd_sc_hd__fa_1
XFILLER_133_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1629_ clknet_leaf_221_clk booth_b2_m41 VGND VGND VPWR VPWR pp_row43_1 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_71_4 pp_row71_24 pp_row71_25 pp_row71_26 VGND VGND VPWR VPWR c$734 s$735
+ sky130_fd_sc_hd__fa_1
XFILLER_143_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_64_3 pp_row64_27 pp_row64_28 pp_row64_29 VGND VGND VPWR VPWR c$606 s$607
+ sky130_fd_sc_hd__fa_1
XFILLER_115_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$5_1880 VGND VGND VPWR VPWR U$$5_1880/HI net1880 sky130_fd_sc_hd__conb_1
Xdadda_fa_4_41_2 s$2169 s$2171 s$2173 VGND VGND VPWR VPWR c$2940 s$2941 sky130_fd_sc_hd__fa_1
Xdadda_fa_1_57_2 pp_row57_14 pp_row57_15 pp_row57_16 VGND VGND VPWR VPWR c$478 s$479
+ sky130_fd_sc_hd__fa_1
XFILLER_100_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_34_1 c$2106 c$2108 s$2111 VGND VGND VPWR VPWR c$2896 s$2897 sky130_fd_sc_hd__fa_1
XFILLER_39_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_11_0 s$3443 c$3916 s$3919 VGND VGND VPWR VPWR c$4174 s$4175 sky130_fd_sc_hd__fa_1
Xdadda_fa_4_27_0 s$1073 c$2046 c$2048 VGND VGND VPWR VPWR c$2852 s$2853 sky130_fd_sc_hd__fa_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_0_60_4 pp_row60_12 pp_row60_13 VGND VGND VPWR VPWR c$48 s$49 sky130_fd_sc_hd__ha_1
Xdadda_fa_3_79_3 s$1679 s$1681 s$1683 VGND VGND VPWR VPWR c$2476 s$2477 sky130_fd_sc_hd__fa_1
XFILLER_96_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4304 t$6604 net1256 VGND VGND VPWR VPWR booth_b62_m25 sky130_fd_sc_hd__xor2_1
XFILLER_78_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4315 net1029 net422 net1021 net704 VGND VGND VPWR VPWR t$6610 sky130_fd_sc_hd__a22o_1
XU$$4326 t$6615 net1261 VGND VGND VPWR VPWR booth_b62_m36 sky130_fd_sc_hd__xor2_1
Xfanout880 net882 VGND VGND VPWR VPWR net880 sky130_fd_sc_hd__buf_6
XU$$4337 net1751 net424 net1743 net706 VGND VGND VPWR VPWR t$6621 sky130_fd_sc_hd__a22o_1
Xfanout891 sel_1$5178 VGND VGND VPWR VPWR net891 sky130_fd_sc_hd__buf_6
XU$$3603 t$6246 net1324 VGND VGND VPWR VPWR booth_b52_m17 sky130_fd_sc_hd__xor2_1
XU$$4348 t$6626 net1260 VGND VGND VPWR VPWR booth_b62_m47 sky130_fd_sc_hd__xor2_1
XU$$3614 net1102 net476 net1094 net749 VGND VGND VPWR VPWR t$6252 sky130_fd_sc_hd__a22o_1
XU$$4359 net1645 net423 net1636 net705 VGND VGND VPWR VPWR t$6632 sky130_fd_sc_hd__a22o_1
XFILLER_46_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3625 t$6257 net1321 VGND VGND VPWR VPWR booth_b52_m28 sky130_fd_sc_hd__xor2_1
XU$$3636 net995 net477 net984 net750 VGND VGND VPWR VPWR t$6263 sky130_fd_sc_hd__a22o_1
XU$$2902 t$5888 net1372 VGND VGND VPWR VPWR booth_b42_m9 sky130_fd_sc_hd__xor2_1
XU$$3647 t$6268 net1324 VGND VGND VPWR VPWR booth_b52_m39 sky130_fd_sc_hd__xor2_1
XFILLER_46_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2913 net1179 net526 net1170 net799 VGND VGND VPWR VPWR t$5894 sky130_fd_sc_hd__a22o_1
XTAP_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3658 net1726 net482 net1717 net755 VGND VGND VPWR VPWR t$6274 sky130_fd_sc_hd__a22o_1
XTAP_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3669 t$6279 net1328 VGND VGND VPWR VPWR booth_b52_m50 sky130_fd_sc_hd__xor2_1
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2924 t$5899 net1368 VGND VGND VPWR VPWR booth_b42_m20 sky130_fd_sc_hd__xor2_1
XU$$2935 net1078 net524 net1070 net797 VGND VGND VPWR VPWR t$5905 sky130_fd_sc_hd__a22o_1
XFILLER_33_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2946 t$5910 net1367 VGND VGND VPWR VPWR booth_b42_m31 sky130_fd_sc_hd__xor2_1
XTAP_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2957 net966 net521 net959 net794 VGND VGND VPWR VPWR t$5916 sky130_fd_sc_hd__a22o_1
XANTENNA_240 net1506 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2968 t$5921 net1369 VGND VGND VPWR VPWR booth_b42_m42 sky130_fd_sc_hd__xor2_1
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_251 net1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_262 net1723 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2979 net1697 net522 net1689 net795 VGND VGND VPWR VPWR t$5927 sky130_fd_sc_hd__a22o_1
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_273 net1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_284 s$4213 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_295 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1980_ clknet_leaf_78_clk booth_b0_m55 VGND VGND VPWR VPWR pp_row55_0 sky130_fd_sc_hd__dfxtp_1
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0931_ clknet_leaf_112_clk booth_b50_m47 VGND VGND VPWR VPWR pp_row97_9 sky130_fd_sc_hd__dfxtp_1
X_0862_ clknet_leaf_105_clk booth_b34_m60 VGND VGND VPWR VPWR pp_row94_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_174_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0793_ clknet_leaf_93_clk booth_b28_m63 VGND VGND VPWR VPWR pp_row91_1 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_248_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_248_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_81_3 c$902 c$904 s$907 VGND VGND VPWR VPWR c$1704 s$1705 sky130_fd_sc_hd__fa_1
XFILLER_177_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2463_ clknet_leaf_94_clk booth_b36_m32 VGND VGND VPWR VPWR pp_row68_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_114_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_717 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_74_2 c$772 c$774 c$776 VGND VGND VPWR VPWR c$1618 s$1619 sky130_fd_sc_hd__fa_1
X_1414_ clknet_leaf_40_clk booth_b0_m34 VGND VGND VPWR VPWR pp_row34_0 sky130_fd_sc_hd__dfxtp_1
X_2394_ clknet_leaf_96_clk booth_b42_m24 VGND VGND VPWR VPWR pp_row66_21 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_51_1 s$2997 s$2999 s$3001 VGND VGND VPWR VPWR c$3602 s$3603 sky130_fd_sc_hd__fa_1
Xdadda_fa_2_67_1 c$640 c$642 c$644 VGND VGND VPWR VPWR c$1532 s$1533 sky130_fd_sc_hd__fa_2
XFILLER_96_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$908 final_adder.$signal$1196 final_adder.g_new$985 final_adder.$signal$214
+ VGND VGND VPWR VPWR final_adder.g_new$1036 sky130_fd_sc_hd__a21o_1
X_1345_ clknet_leaf_3_clk booth_b22_m8 VGND VGND VPWR VPWR pp_row30_11 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_44_0 c$2948 c$2950 c$2952 VGND VGND VPWR VPWR c$3572 s$3573 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$919 final_adder.$signal$1174 final_adder.g_new$1007 final_adder.$signal$170
+ VGND VGND VPWR VPWR final_adder.g_new$1047 sky130_fd_sc_hd__a21o_1
XFILLER_111_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1276_ clknet_leaf_8_clk booth_b26_m0 VGND VGND VPWR VPWR pp_row26_13 sky130_fd_sc_hd__dfxtp_1
X_0227_ clknet_leaf_208_clk booth_b28_m43 VGND VGND VPWR VPWR pp_row71_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_36_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_239_clk clknet_5_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_239_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_192_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_89_2 s$2553 s$2555 s$2557 VGND VGND VPWR VPWR c$3228 s$3229 sky130_fd_sc_hd__fa_1
XFILLER_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_59_0 s$3635 c$4012 s$4015 VGND VGND VPWR VPWR c$4270 s$4271 sky130_fd_sc_hd__fa_1
XFILLER_161_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1108 net1110 VGND VGND VPWR VPWR net1108 sky130_fd_sc_hd__buf_4
XFILLER_160_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1119 net1120 VGND VGND VPWR VPWR net1119 sky130_fd_sc_hd__buf_6
XU$$2198_1773 VGND VGND VPWR VPWR U$$2198_1773/HI net1773 sky130_fd_sc_hd__conb_1
XFILLER_86_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_62_0 pp_row62_17 pp_row62_18 pp_row62_19 VGND VGND VPWR VPWR c$564 s$565
+ sky130_fd_sc_hd__fa_1
XFILLER_75_826 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2209 t$5534 net1432 VGND VGND VPWR VPWR booth_b32_m5 sky130_fd_sc_hd__xor2_1
XFILLER_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1508 net15 VGND VGND VPWR VPWR notblock$5175\[1\] sky130_fd_sc_hd__inv_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1519 net1031 net611 net932 net884 VGND VGND VPWR VPWR t$5182 sky130_fd_sc_hd__a22o_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_975 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_91_2 c$1816 s$1819 s$1821 VGND VGND VPWR VPWR c$2570 s$2571 sky130_fd_sc_hd__fa_1
XFILLER_100_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_84_1 c$1726 c$1728 c$1730 VGND VGND VPWR VPWR c$2512 s$2513 sky130_fd_sc_hd__fa_1
XFILLER_3_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_6_61_0 c$3636 c$3638 s$3641 VGND VGND VPWR VPWR c$4018 s$4019 sky130_fd_sc_hd__fa_1
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_77_0 s$851 c$1638 c$1640 VGND VGND VPWR VPWR c$2454 s$2455 sky130_fd_sc_hd__fa_1
XFILLER_97_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1620 net1621 VGND VGND VPWR VPWR net1620 sky130_fd_sc_hd__buf_4
Xfanout1631 net1632 VGND VGND VPWR VPWR net1631 sky130_fd_sc_hd__buf_6
Xfanout1642 net112 VGND VGND VPWR VPWR net1642 sky130_fd_sc_hd__clkbuf_4
Xfanout1653 net111 VGND VGND VPWR VPWR net1653 sky130_fd_sc_hd__clkbuf_4
XU$$4101 net1557 net453 net1549 net726 VGND VGND VPWR VPWR t$6500 sky130_fd_sc_hd__a22o_1
XFILLER_65_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4112 net1265 VGND VGND VPWR VPWR notblock$6505\[2\] sky130_fd_sc_hd__inv_1
Xfanout1664 net1666 VGND VGND VPWR VPWR net1664 sky130_fd_sc_hd__buf_6
Xfanout1675 net1678 VGND VGND VPWR VPWR net1675 sky130_fd_sc_hd__clkbuf_4
XU$$4123 t$6512 net1264 VGND VGND VPWR VPWR booth_b60_m3 sky130_fd_sc_hd__xor2_1
X_1130_ clknet_leaf_13_clk booth_b12_m4 VGND VGND VPWR VPWR pp_row16_6 sky130_fd_sc_hd__dfxtp_1
XU$$4134 net127 net438 net1502 net720 VGND VGND VPWR VPWR t$6518 sky130_fd_sc_hd__a22o_1
Xfanout1686 net108 VGND VGND VPWR VPWR net1686 sky130_fd_sc_hd__buf_2
XU$$3400 net1644 net499 net1636 net772 VGND VGND VPWR VPWR t$6142 sky130_fd_sc_hd__a22o_1
XU$$4145 t$6523 net1263 VGND VGND VPWR VPWR booth_b60_m14 sky130_fd_sc_hd__xor2_1
Xfanout1697 net106 VGND VGND VPWR VPWR net1697 sky130_fd_sc_hd__buf_6
XFILLER_66_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4156 net1136 net435 net1120 net717 VGND VGND VPWR VPWR t$6529 sky130_fd_sc_hd__a22o_1
XU$$3411 t$6147 net1345 VGND VGND VPWR VPWR booth_b48_m58 sky130_fd_sc_hd__xor2_1
XU$$3422 net1533 net499 net1792 net772 VGND VGND VPWR VPWR t$6153 sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_113_1 pp_row113_9 c$2732 c$2734 VGND VGND VPWR VPWR c$3370 s$3371 sky130_fd_sc_hd__fa_1
XU$$4167 t$6534 net1268 VGND VGND VPWR VPWR booth_b60_m25 sky130_fd_sc_hd__xor2_1
XU$$4178 net1029 net438 net1021 net720 VGND VGND VPWR VPWR t$6540 sky130_fd_sc_hd__a22o_1
XU$$3433 net1229 net484 net1124 net757 VGND VGND VPWR VPWR t$6160 sky130_fd_sc_hd__a22o_1
X_1061_ clknet_leaf_129_clk booth_b62_m60 VGND VGND VPWR VPWR pp_row122_3 sky130_fd_sc_hd__dfxtp_1
XU$$4189 t$6545 net1269 VGND VGND VPWR VPWR booth_b60_m36 sky130_fd_sc_hd__xor2_1
XU$$3444 t$6165 net1337 VGND VGND VPWR VPWR booth_b50_m6 sky130_fd_sc_hd__xor2_1
XFILLER_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2710 t$5789 net1397 VGND VGND VPWR VPWR booth_b38_m50 sky130_fd_sc_hd__xor2_1
XU$$3455 net1214 net487 net1205 net760 VGND VGND VPWR VPWR t$6171 sky130_fd_sc_hd__a22o_1
XU$$3466 t$6176 net1333 VGND VGND VPWR VPWR booth_b50_m17 sky130_fd_sc_hd__xor2_1
XU$$2721 net1618 net547 net1609 net820 VGND VGND VPWR VPWR t$5795 sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_106_0 s$1969 c$2678 c$2680 VGND VGND VPWR VPWR c$3326 s$3327 sky130_fd_sc_hd__fa_1
Xdadda_fa_2_39_5 c$220 s$223 s$225 VGND VGND VPWR VPWR c$1204 s$1205 sky130_fd_sc_hd__fa_1
XU$$2732 t$5800 net1400 VGND VGND VPWR VPWR booth_b38_m61 sky130_fd_sc_hd__xor2_1
XTAP_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3477 net1102 net484 net1090 net757 VGND VGND VPWR VPWR t$6182 sky130_fd_sc_hd__a22o_1
XTAP_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3488 t$6187 net1331 VGND VGND VPWR VPWR booth_b50_m28 sky130_fd_sc_hd__xor2_1
XU$$2743 net1378 notblock$5805\[1\] VGND VGND VPWR VPWR t$5806 sky130_fd_sc_hd__and2_1
XTAP_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3499 net995 net485 net984 net758 VGND VGND VPWR VPWR t$6193 sky130_fd_sc_hd__a22o_1
XU$$2754 net934 net535 net1673 net808 VGND VGND VPWR VPWR t$5813 sky130_fd_sc_hd__a22o_1
XU$$2765 t$5818 net1377 VGND VGND VPWR VPWR booth_b40_m9 sky130_fd_sc_hd__xor2_1
XU$$2776 net1181 net539 net1172 net812 VGND VGND VPWR VPWR t$5824 sky130_fd_sc_hd__a22o_1
XU$$2787 t$5829 net1376 VGND VGND VPWR VPWR booth_b40_m20 sky130_fd_sc_hd__xor2_1
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2798 net1078 net542 net1070 net815 VGND VGND VPWR VPWR t$5835 sky130_fd_sc_hd__a22o_1
XFILLER_33_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1963_ clknet_leaf_63_clk booth_b28_m26 VGND VGND VPWR VPWR pp_row54_14 sky130_fd_sc_hd__dfxtp_1
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0914_ clknet_leaf_104_clk booth_b54_m42 VGND VGND VPWR VPWR pp_row96_12 sky130_fd_sc_hd__dfxtp_1
X_1894_ clknet_leaf_137_clk booth_b60_m47 VGND VGND VPWR VPWR pp_row107_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_175_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_99_1 s$3285 s$3287 s$3289 VGND VGND VPWR VPWR c$3794 s$3795 sky130_fd_sc_hd__fa_1
XFILLER_88_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0845_ clknet_leaf_105_clk booth_b40_m53 VGND VGND VPWR VPWR pp_row93_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0776_ clknet_leaf_141_clk booth_b40_m50 VGND VGND VPWR VPWR pp_row90_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_143_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2446_ clknet_leaf_90_clk booth_b6_m62 VGND VGND VPWR VPWR pp_row68_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_124_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2377_ clknet_leaf_83_clk booth_b14_m52 VGND VGND VPWR VPWR pp_row66_7 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$705 final_adder.p_new$712 final_adder.g_new$729 final_adder.g_new$713
+ VGND VGND VPWR VPWR final_adder.g_new$833 sky130_fd_sc_hd__a21o_1
XFILLER_111_761 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$716 final_adder.p_new$740 final_adder.p_new$724 VGND VGND VPWR VPWR
+ final_adder.p_new$844 sky130_fd_sc_hd__and2_1
XFILLER_25_1068 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$727 final_adder.p_new$734 final_adder.g_new$751 final_adder.g_new$735
+ VGND VGND VPWR VPWR final_adder.g_new$855 sky130_fd_sc_hd__a21o_2
X_1328_ clknet_leaf_4_clk booth_b22_m7 VGND VGND VPWR VPWR pp_row29_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_57_859 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$749 final_adder.p_new$764 final_adder.g_new$797 final_adder.g_new$765
+ VGND VGND VPWR VPWR final_adder.g_new$877 sky130_fd_sc_hd__a21o_1
XFILLER_56_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1259_ clknet_leaf_9_clk booth_b24_m1 VGND VGND VPWR VPWR pp_row25_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_71_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_88_0_1900 VGND VGND VPWR VPWR net1900 dadda_fa_1_88_0_1900/LO sky130_fd_sc_hd__conb_1
XFILLER_177_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_94_0 s$1865 c$2582 c$2584 VGND VGND VPWR VPWR c$3254 s$3255 sky130_fd_sc_hd__fa_1
XFILLER_193_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_108_2 pp_row108_8 pp_row108_9 pp_row108_10 VGND VGND VPWR VPWR c$2706
+ s$2707 sky130_fd_sc_hd__fa_1
XFILLER_165_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput280 net280 VGND VGND VPWR VPWR o[120] sky130_fd_sc_hd__buf_2
Xoutput291 net291 VGND VGND VPWR VPWR o[15] sky130_fd_sc_hd__buf_2
XFILLER_102_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2006 net930 net591 net1751 net864 VGND VGND VPWR VPWR t$5430 sky130_fd_sc_hd__a22o_1
XU$$2017 t$5435 net1450 VGND VGND VPWR VPWR booth_b28_m46 sky130_fd_sc_hd__xor2_1
XU$$2028 net1647 net589 net1639 net862 VGND VGND VPWR VPWR t$5441 sky130_fd_sc_hd__a22o_1
XU$$2039 t$5446 net1453 VGND VGND VPWR VPWR booth_b28_m57 sky130_fd_sc_hd__xor2_1
XU$$1305 net1000 net638 net992 net911 VGND VGND VPWR VPWR t$5072 sky130_fd_sc_hd__a22o_1
XFILLER_167_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1316 t$5077 net1666 VGND VGND VPWR VPWR booth_b18_m38 sky130_fd_sc_hd__xor2_1
XU$$1327 net1729 net636 net1720 net909 VGND VGND VPWR VPWR t$5083 sky130_fd_sc_hd__a22o_1
XFILLER_128_1023 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1338 t$5088 net1670 VGND VGND VPWR VPWR booth_b18_m49 sky130_fd_sc_hd__xor2_1
XU$$1349 net1620 net640 net1612 net913 VGND VGND VPWR VPWR t$5094 sky130_fd_sc_hd__a22o_1
XFILLER_15_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0630_ clknet_leaf_178_clk booth_b46_m38 VGND VGND VPWR VPWR pp_row84_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0561_ clknet_leaf_186_clk booth_b20_m62 VGND VGND VPWR VPWR pp_row82_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_180_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2300_ clknet_leaf_198_clk booth_b6_m58 VGND VGND VPWR VPWR pp_row64_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_125_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4515_1878 VGND VGND VPWR VPWR U$$4515_1878/HI net1878 sky130_fd_sc_hd__conb_1
XFILLER_97_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0492_ clknet_leaf_159_clk booth_b50_m29 VGND VGND VPWR VPWR pp_row79_18 sky130_fd_sc_hd__dfxtp_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2231_ clknet_leaf_233_clk booth_b16_m46 VGND VGND VPWR VPWR pp_row62_8 sky130_fd_sc_hd__dfxtp_1
Xfanout1450 net1456 VGND VGND VPWR VPWR net1450 sky130_fd_sc_hd__buf_6
XFILLER_79_995 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1461 net1462 VGND VGND VPWR VPWR net1461 sky130_fd_sc_hd__buf_2
Xdadda_fa_2_51_4 s$371 s$373 s$375 VGND VGND VPWR VPWR c$1346 s$1347 sky130_fd_sc_hd__fa_1
Xfanout1472 net1473 VGND VGND VPWR VPWR net1472 sky130_fd_sc_hd__clkbuf_4
X_2162_ clknet_leaf_214_clk booth_b22_m38 VGND VGND VPWR VPWR pp_row60_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1483 net1484 VGND VGND VPWR VPWR net1483 sky130_fd_sc_hd__buf_8
Xfanout1494 net1495 VGND VGND VPWR VPWR net1494 sky130_fd_sc_hd__buf_4
XFILLER_65_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1113_ clknet_leaf_13_clk booth_b0_m15 VGND VGND VPWR VPWR pp_row15_0 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_44_3 c$256 c$258 c$260 VGND VGND VPWR VPWR c$1260 s$1261 sky130_fd_sc_hd__fa_1
XFILLER_38_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3230 t$6055 net1351 VGND VGND VPWR VPWR booth_b46_m36 sky130_fd_sc_hd__xor2_1
X_2093_ clknet_leaf_149_clk booth_b24_m34 VGND VGND VPWR VPWR pp_row58_12 sky130_fd_sc_hd__dfxtp_1
XU$$3241 net1748 net504 net1740 net777 VGND VGND VPWR VPWR t$6061 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$12 c$4174 s$4177 VGND VGND VPWR VPWR final_adder.$signal$26 final_adder.$signal$1102
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$23 c$4196 s$4199 VGND VGND VPWR VPWR final_adder.$signal$48 final_adder.$signal$1113
+ sky130_fd_sc_hd__ha_2
XU$$3252 t$6066 net1355 VGND VGND VPWR VPWR booth_b46_m47 sky130_fd_sc_hd__xor2_1
XFILLER_19_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_37_2 pp_row37_11 pp_row37_12 pp_row37_13 VGND VGND VPWR VPWR c$1174 s$1175
+ sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$34 c$4218 s$4221 VGND VGND VPWR VPWR final_adder.$signal$70 final_adder.$signal$1124
+ sky130_fd_sc_hd__ha_1
XU$$3263 net1644 net508 net1635 net781 VGND VGND VPWR VPWR t$6072 sky130_fd_sc_hd__a22o_1
X_1044_ clknet_leaf_56_clk net1249 VGND VGND VPWR VPWR pp_row6_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3274 t$6077 net1356 VGND VGND VPWR VPWR booth_b46_m58 sky130_fd_sc_hd__xor2_1
XFILLER_0_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$45 c$4240 s$4243 VGND VGND VPWR VPWR final_adder.$signal$92 final_adder.$signal$1135
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$56 c$4262 s$4265 VGND VGND VPWR VPWR final_adder.$signal$114 final_adder.$signal$1146
+ sky130_fd_sc_hd__ha_1
XFILLER_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2540 net994 net555 net984 net828 VGND VGND VPWR VPWR t$5703 sky130_fd_sc_hd__a22o_1
XU$$3285 net1532 net504 net1790 net777 VGND VGND VPWR VPWR t$6083 sky130_fd_sc_hd__a22o_1
XU$$2551 t$5708 net1409 VGND VGND VPWR VPWR booth_b36_m39 sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_14_1 s$2775 s$2777 s$2779 VGND VGND VPWR VPWR c$3454 s$3455 sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$67 c$4284 s$4287 VGND VGND VPWR VPWR final_adder.$signal$136 final_adder.$signal$1157
+ sky130_fd_sc_hd__ha_1
XU$$3296 net1229 net493 net1125 net766 VGND VGND VPWR VPWR t$6090 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$78 c$4306 s$4309 VGND VGND VPWR VPWR final_adder.$signal$158 final_adder.$signal$1168
+ sky130_fd_sc_hd__ha_1
XU$$2562 net1723 net556 net1713 net829 VGND VGND VPWR VPWR t$5714 sky130_fd_sc_hd__a22o_1
XU$$2573 t$5719 net1408 VGND VGND VPWR VPWR booth_b36_m50 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$89 c$4328 s$4331 VGND VGND VPWR VPWR final_adder.$signal$180 final_adder.$signal$1179
+ sky130_fd_sc_hd__ha_2
XU$$2584 net1618 net557 net1609 net830 VGND VGND VPWR VPWR t$5725 sky130_fd_sc_hd__a22o_1
XU$$2595 t$5730 net1410 VGND VGND VPWR VPWR booth_b36_m61 sky130_fd_sc_hd__xor2_1
XFILLER_55_1039 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1850 t$5350 net1460 VGND VGND VPWR VPWR booth_b26_m31 sky130_fd_sc_hd__xor2_1
XU$$1861 net965 net598 net957 net871 VGND VGND VPWR VPWR t$5356 sky130_fd_sc_hd__a22o_1
XU$$1872 t$5361 net1465 VGND VGND VPWR VPWR booth_b26_m42 sky130_fd_sc_hd__xor2_1
XU$$1883 net1695 net598 net1687 net871 VGND VGND VPWR VPWR t$5367 sky130_fd_sc_hd__a22o_1
XU$$1894 t$5372 net1464 VGND VGND VPWR VPWR booth_b26_m53 sky130_fd_sc_hd__xor2_1
X_1946_ clknet_leaf_78_clk booth_b0_m54 VGND VGND VPWR VPWR pp_row54_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1877_ clknet_leaf_70_clk booth_b42_m9 VGND VGND VPWR VPWR pp_row51_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_147_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0828_ clknet_leaf_108_clk booth_b52_m40 VGND VGND VPWR VPWR pp_row92_13 sky130_fd_sc_hd__dfxtp_1
X_0759_ clknet_leaf_153_clk booth_b50_m39 VGND VGND VPWR VPWR pp_row89_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_89_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2429_ clknet_leaf_96_clk booth_b38_m29 VGND VGND VPWR VPWR pp_row67_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_130_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$513 final_adder.p_new$516 final_adder.g_new$525 final_adder.g_new$517
+ VGND VGND VPWR VPWR final_adder.g_new$641 sky130_fd_sc_hd__a21o_1
XFILLER_130_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$524 final_adder.p_new$536 final_adder.p_new$528 VGND VGND VPWR VPWR
+ final_adder.p_new$652 sky130_fd_sc_hd__and2_1
XTAP_3806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$535 final_adder.p_new$538 final_adder.g_new$547 final_adder.g_new$539
+ VGND VGND VPWR VPWR final_adder.g_new$663 sky130_fd_sc_hd__a21o_1
XTAP_3817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$546 final_adder.p_new$558 final_adder.p_new$550 VGND VGND VPWR VPWR
+ final_adder.p_new$674 sky130_fd_sc_hd__and2_1
XTAP_3828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$557 final_adder.p_new$560 final_adder.g_new$569 final_adder.g_new$561
+ VGND VGND VPWR VPWR final_adder.g_new$685 sky130_fd_sc_hd__a21o_1
XTAP_3839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$568 final_adder.p_new$580 final_adder.p_new$572 VGND VGND VPWR VPWR
+ final_adder.p_new$696 sky130_fd_sc_hd__and2_1
XU$$407 t$4612 net1281 VGND VGND VPWR VPWR booth_b4_m63 sky130_fd_sc_hd__xor2_1
XU$$418 t$4619 net1248 VGND VGND VPWR VPWR booth_b6_m0 sky130_fd_sc_hd__xor2_1
XFILLER_56_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$579 final_adder.p_new$582 final_adder.g_new$591 final_adder.g_new$583
+ VGND VGND VPWR VPWR final_adder.g_new$707 sky130_fd_sc_hd__a21o_1
XU$$429 net1564 net429 net1523 net711 VGND VGND VPWR VPWR t$4625 sky130_fd_sc_hd__a22o_1
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_16__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_5_16__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_113_0 pp_row113_0 pp_row113_1 pp_row113_2 VGND VGND VPWR VPWR c$2738 s$2739
+ sky130_fd_sc_hd__fa_1
XFILLER_153_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_61_3 s$1463 s$1465 s$1467 VGND VGND VPWR VPWR c$2332 s$2333 sky130_fd_sc_hd__fa_1
XFILLER_79_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_54_2 c$1372 s$1375 s$1377 VGND VGND VPWR VPWR c$2274 s$2275 sky130_fd_sc_hd__fa_1
XFILLER_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_47_1 c$1282 c$1284 c$1286 VGND VGND VPWR VPWR c$2216 s$2217 sky130_fd_sc_hd__fa_1
XFILLER_85_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_24_0 c$3488 c$3490 s$3493 VGND VGND VPWR VPWR c$3944 s$3945 sky130_fd_sc_hd__fa_1
XU$$930 net1656 net400 net1648 net666 VGND VGND VPWR VPWR t$4880 sky130_fd_sc_hd__a22o_1
XU$$941 t$4885 net1318 VGND VGND VPWR VPWR booth_b12_m56 sky130_fd_sc_hd__xor2_1
XU$$952 net1546 net395 net1538 net661 VGND VGND VPWR VPWR t$4891 sky130_fd_sc_hd__a22o_1
XU$$963 notblock$4895\[2\] net6 net1316 t$4896 notblock$4895\[0\] VGND VGND VPWR VPWR
+ sel_0$4897 sky130_fd_sc_hd__a32o_1
XU$$1102 net1755 net643 net1228 net916 VGND VGND VPWR VPWR t$4969 sky130_fd_sc_hd__a22o_1
XFILLER_44_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$974 t$4903 net1185 VGND VGND VPWR VPWR booth_b14_m4 sky130_fd_sc_hd__xor2_1
XU$$1113 t$4974 net1009 VGND VGND VPWR VPWR booth_b16_m5 sky130_fd_sc_hd__xor2_1
XU$$1124 net1219 net643 net1210 net916 VGND VGND VPWR VPWR t$4980 sky130_fd_sc_hd__a22o_1
XU$$985 net1496 net385 net1221 net651 VGND VGND VPWR VPWR t$4909 sky130_fd_sc_hd__a22o_1
XU$$996 t$4914 net1183 VGND VGND VPWR VPWR booth_b14_m15 sky130_fd_sc_hd__xor2_1
XU$$1135 t$4985 net1010 VGND VGND VPWR VPWR booth_b16_m16 sky130_fd_sc_hd__xor2_1
XU$$1146 net1106 net646 net1100 net919 VGND VGND VPWR VPWR t$4991 sky130_fd_sc_hd__a22o_1
XFILLER_188_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1157 t$4996 net1007 VGND VGND VPWR VPWR booth_b16_m27 sky130_fd_sc_hd__xor2_1
XU$$1168 net999 net644 net991 net917 VGND VGND VPWR VPWR t$5002 sky130_fd_sc_hd__a22o_1
Xdadda_ha_3_112_2 pp_row112_6 pp_row112_7 VGND VGND VPWR VPWR c$2736 s$2737 sky130_fd_sc_hd__ha_1
XFILLER_189_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1179 t$5007 net1010 VGND VGND VPWR VPWR booth_b16_m38 sky130_fd_sc_hd__xor2_1
XFILLER_188_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1800_ clknet_leaf_220_clk booth_b12_m37 VGND VGND VPWR VPWR pp_row49_6 sky130_fd_sc_hd__dfxtp_1
X_1731_ clknet_leaf_24_clk booth_b42_m4 VGND VGND VPWR VPWR pp_row46_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1015 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1075 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1662_ clknet_leaf_21_clk booth_b16_m28 VGND VGND VPWR VPWR pp_row44_8 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_99_4 pp_row99_12 pp_row99_13 pp_row99_14 VGND VGND VPWR VPWR c$1922 s$1923
+ sky130_fd_sc_hd__fa_2
XFILLER_176_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0613_ clknet_leaf_173_clk booth_b62_m21 VGND VGND VPWR VPWR pp_row83_22 sky130_fd_sc_hd__dfxtp_1
XFILLER_160_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1593_ clknet_leaf_6_clk booth_b32_m9 VGND VGND VPWR VPWR pp_row41_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_171_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0544_ clknet_leaf_126_clk booth_b54_m62 VGND VGND VPWR VPWR pp_row116_2 sky130_fd_sc_hd__dfxtp_1
Xfanout709 net710 VGND VGND VPWR VPWR net709 sky130_fd_sc_hd__buf_6
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0475_ clknet_leaf_186_clk booth_b20_m59 VGND VGND VPWR VPWR pp_row79_3 sky130_fd_sc_hd__dfxtp_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2214_ clknet_leaf_217_clk booth_b50_m11 VGND VGND VPWR VPWR pp_row61_25 sky130_fd_sc_hd__dfxtp_1
XFILLER_61_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1280 net1281 VGND VGND VPWR VPWR net1280 sky130_fd_sc_hd__buf_6
Xfanout1291 net1295 VGND VGND VPWR VPWR net1291 sky130_fd_sc_hd__buf_6
X_2145_ clknet_leaf_31_clk booth_b54_m5 VGND VGND VPWR VPWR pp_row59_27 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_42_0 pp_row42_14 pp_row42_15 pp_row42_16 VGND VGND VPWR VPWR c$1230 s$1231
+ sky130_fd_sc_hd__fa_1
XFILLER_27_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3060 net1137 net514 net1121 net787 VGND VGND VPWR VPWR t$5969 sky130_fd_sc_hd__a22o_1
XFILLER_82_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2076_ clknet_leaf_85_clk booth_b52_m5 VGND VGND VPWR VPWR pp_row57_26 sky130_fd_sc_hd__dfxtp_1
XU$$3071 t$5974 net1358 VGND VGND VPWR VPWR booth_b44_m25 sky130_fd_sc_hd__xor2_1
XU$$3082 net1027 net512 net1019 net785 VGND VGND VPWR VPWR t$5980 sky130_fd_sc_hd__a22o_1
X_1027_ clknet_leaf_120_clk booth_b42_m60 VGND VGND VPWR VPWR pp_row102_3 sky130_fd_sc_hd__dfxtp_1
XU$$3093 t$5985 net1360 VGND VGND VPWR VPWR booth_b44_m36 sky130_fd_sc_hd__xor2_1
XU$$2370 t$5616 net1423 VGND VGND VPWR VPWR booth_b34_m17 sky130_fd_sc_hd__xor2_1
XFILLER_34_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2381 net1100 net560 net1091 net833 VGND VGND VPWR VPWR t$5622 sky130_fd_sc_hd__a22o_1
XU$$2392 t$5627 net1425 VGND VGND VPWR VPWR booth_b34_m28 sky130_fd_sc_hd__xor2_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1680 net1175 net603 net1166 net876 VGND VGND VPWR VPWR t$5264 sky130_fd_sc_hd__a22o_1
XU$$1691 t$5269 net1467 VGND VGND VPWR VPWR booth_b24_m20 sky130_fd_sc_hd__xor2_1
XFILLER_22_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1929_ clknet_leaf_67_clk booth_b24_m29 VGND VGND VPWR VPWR pp_row53_12 sky130_fd_sc_hd__dfxtp_1
Xdadda_ha_1_88_4 pp_row88_12 pp_row88_13 VGND VGND VPWR VPWR c$1008 s$1009 sky130_fd_sc_hd__ha_1
XFILLER_107_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_71_2 s$2409 s$2411 s$2413 VGND VGND VPWR VPWR c$3120 s$3121 sky130_fd_sc_hd__fa_1
Xdadda_fa_1_87_2 pp_row87_6 pp_row87_7 pp_row87_8 VGND VGND VPWR VPWR c$994 s$995
+ sky130_fd_sc_hd__fa_1
XFILLER_104_845 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_64_1 c$2346 c$2348 s$2351 VGND VGND VPWR VPWR c$3076 s$3077 sky130_fd_sc_hd__fa_1
XFILLER_104_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_41_0 s$3563 c$3976 s$3979 VGND VGND VPWR VPWR c$4234 s$4235 sky130_fd_sc_hd__fa_2
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_57_0 s$1421 c$2286 c$2288 VGND VGND VPWR VPWR c$3032 s$3033 sky130_fd_sc_hd__fa_1
XTAP_4304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$310 final_adder.p_new$312 final_adder.p_new$310 VGND VGND VPWR VPWR
+ final_adder.p_new$438 sky130_fd_sc_hd__and2_1
XFILLER_162_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$321 final_adder.p_new$320 final_adder.g_new$323 final_adder.g_new$321
+ VGND VGND VPWR VPWR final_adder.g_new$449 sky130_fd_sc_hd__a21o_1
XTAP_4337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$332 final_adder.p_new$334 final_adder.p_new$332 VGND VGND VPWR VPWR
+ final_adder.p_new$460 sky130_fd_sc_hd__and2_1
XTAP_4359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$343 final_adder.p_new$342 final_adder.g_new$345 final_adder.g_new$343
+ VGND VGND VPWR VPWR final_adder.g_new$471 sky130_fd_sc_hd__a21o_1
XTAP_3625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$354 final_adder.p_new$356 final_adder.p_new$354 VGND VGND VPWR VPWR
+ final_adder.p_new$482 sky130_fd_sc_hd__and2_1
XTAP_3636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$204 t$4509 net1386 VGND VGND VPWR VPWR booth_b2_m30 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$365 final_adder.p_new$364 final_adder.g_new$367 final_adder.g_new$365
+ VGND VGND VPWR VPWR final_adder.g_new$493 sky130_fd_sc_hd__a21o_1
XTAP_3647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$376 final_adder.p_new$378 final_adder.p_new$376 VGND VGND VPWR VPWR
+ final_adder.p_new$504 sky130_fd_sc_hd__and2_1
XU$$215 net974 net625 net965 net898 VGND VGND VPWR VPWR t$4515 sky130_fd_sc_hd__a22o_1
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$226 t$4520 net1387 VGND VGND VPWR VPWR booth_b2_m41 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$387 final_adder.p_new$388 final_adder.g_new$393 final_adder.g_new$389
+ VGND VGND VPWR VPWR final_adder.g_new$515 sky130_fd_sc_hd__a21o_1
XTAP_3669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$398 final_adder.p_new$404 final_adder.p_new$400 VGND VGND VPWR VPWR
+ final_adder.p_new$526 sky130_fd_sc_hd__and2_1
XU$$237 net1706 net626 net1698 net899 VGND VGND VPWR VPWR t$4526 sky130_fd_sc_hd__a22o_1
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$248 t$4531 net1392 VGND VGND VPWR VPWR booth_b2_m52 sky130_fd_sc_hd__xor2_1
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$259 net1596 net622 net1587 net895 VGND VGND VPWR VPWR t$4537 sky130_fd_sc_hd__a22o_1
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1012 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$9 t$4411 net1574 VGND VGND VPWR VPWR booth_b0_m1 sky130_fd_sc_hd__xor2_1
XFILLER_138_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_0_75_0 pp_row75_0 pp_row75_1 pp_row75_2 VGND VGND VPWR VPWR c$192 s$193
+ sky130_fd_sc_hd__fa_1
X_0260_ clknet_leaf_210_clk booth_b28_m44 VGND VGND VPWR VPWR pp_row72_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_121_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0191_ clknet_leaf_148_clk booth_b24_m46 VGND VGND VPWR VPWR pp_row70_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_75_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$760 t$4793 net1413 VGND VGND VPWR VPWR booth_b10_m34 sky130_fd_sc_hd__xor2_1
XFILLER_23_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$771 net940 net403 net924 net669 VGND VGND VPWR VPWR t$4799 sky130_fd_sc_hd__a22o_1
XFILLER_91_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$782 t$4804 net1416 VGND VGND VPWR VPWR booth_b10_m45 sky130_fd_sc_hd__xor2_1
XU$$793 net1654 net403 net1646 net669 VGND VGND VPWR VPWR t$4810 sky130_fd_sc_hd__a22o_1
XFILLER_16_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1714_ clknet_leaf_237_clk booth_b14_m32 VGND VGND VPWR VPWR pp_row46_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_145_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_81_1 s$3177 s$3179 s$3181 VGND VGND VPWR VPWR c$3722 s$3723 sky130_fd_sc_hd__fa_1
Xdadda_fa_2_97_1 pp_row97_3 pp_row97_4 pp_row97_5 VGND VGND VPWR VPWR c$1892 s$1893
+ sky130_fd_sc_hd__fa_1
X_1645_ clknet_leaf_6_clk booth_b32_m11 VGND VGND VPWR VPWR pp_row43_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_74_0 c$3128 c$3130 c$3132 VGND VGND VPWR VPWR c$3692 s$3693 sky130_fd_sc_hd__fa_1
XFILLER_126_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1576_ clknet_leaf_243_clk booth_b0_m41 VGND VGND VPWR VPWR pp_row41_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout506 net509 VGND VGND VPWR VPWR net506 sky130_fd_sc_hd__clkbuf_4
Xfanout517 net518 VGND VGND VPWR VPWR net517 sky130_fd_sc_hd__clkbuf_8
Xdadda_fa_1_73_8 c$178 s$181 s$183 VGND VGND VPWR VPWR c$778 s$779 sky130_fd_sc_hd__fa_2
Xfanout528 net530 VGND VGND VPWR VPWR net528 sky130_fd_sc_hd__clkbuf_4
X_0527_ clknet_leaf_162_clk booth_b60_m20 VGND VGND VPWR VPWR pp_row80_23 sky130_fd_sc_hd__dfxtp_1
Xfanout539 net542 VGND VGND VPWR VPWR net539 sky130_fd_sc_hd__buf_4
XFILLER_101_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_66_7 c$106 s$109 s$111 VGND VGND VPWR VPWR c$650 s$651 sky130_fd_sc_hd__fa_1
X_0458_ clknet_leaf_157_clk booth_b42_m36 VGND VGND VPWR VPWR pp_row78_15 sky130_fd_sc_hd__dfxtp_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_59_6 pp_row59_29 pp_row59_30 c$24 VGND VGND VPWR VPWR c$522 s$523 sky130_fd_sc_hd__fa_1
XFILLER_66_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0389_ clknet_leaf_181_clk net157 VGND VGND VPWR VPWR pp_row125_3 sky130_fd_sc_hd__dfxtp_2
XFILLER_27_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2128_ clknet_leaf_26_clk booth_b22_m37 VGND VGND VPWR VPWR pp_row59_11 sky130_fd_sc_hd__dfxtp_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2059_ clknet_leaf_39_clk booth_b24_m33 VGND VGND VPWR VPWR pp_row57_12 sky130_fd_sc_hd__dfxtp_1
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_876 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_89_0 s$3755 c$4072 s$4075 VGND VGND VPWR VPWR c$4330 s$4331 sky130_fd_sc_hd__fa_2
XFILLER_136_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_92_0 net1902 pp_row92_1 pp_row92_2 VGND VGND VPWR VPWR c$1032 s$1033 sky130_fd_sc_hd__fa_1
XFILLER_150_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4508 net1589 sel_0$6647 net1580 net695 VGND VGND VPWR VPWR t$6708 sky130_fd_sc_hd__a22o_1
XTAP_4112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3807 net1660 net474 net1652 net747 VGND VGND VPWR VPWR t$6350 sky130_fd_sc_hd__a22o_1
XTAP_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$140 final_adder.$signal$1204 final_adder.$signal$1205 VGND VGND VPWR
+ VPWR final_adder.p_new$268 sky130_fd_sc_hd__and2_1
XFILLER_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3818 t$6355 net1306 VGND VGND VPWR VPWR booth_b54_m56 sky130_fd_sc_hd__xor2_1
XTAP_4167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$151 final_adder.$signal$1195 final_adder.$signal$210 final_adder.$signal$212
+ VGND VGND VPWR VPWR final_adder.g_new$279 sky130_fd_sc_hd__a21o_1
XTAP_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3829 net1549 net473 net1541 net746 VGND VGND VPWR VPWR t$6361 sky130_fd_sc_hd__a22o_1
XTAP_4178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_104_0 c$3808 c$3810 s$3813 VGND VGND VPWR VPWR c$4104 s$4105 sky130_fd_sc_hd__fa_1
XTAP_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$162 final_adder.$signal$1182 final_adder.$signal$1183 VGND VGND VPWR
+ VPWR final_adder.p_new$290 sky130_fd_sc_hd__and2_1
XTAP_4189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$173 final_adder.$signal$1173 final_adder.$signal$166 final_adder.$signal$168
+ VGND VGND VPWR VPWR final_adder.g_new$301 sky130_fd_sc_hd__a21o_1
XTAP_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$184 final_adder.$signal$1160 final_adder.$signal$1161 VGND VGND VPWR
+ VPWR final_adder.p_new$312 sky130_fd_sc_hd__and2_1
XTAP_3466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_400 net1631 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$195 final_adder.$signal$1151 final_adder.$signal$122 final_adder.$signal$124
+ VGND VGND VPWR VPWR final_adder.g_new$323 sky130_fd_sc_hd__a21o_1
XFILLER_73_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_411 net1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_422 net526 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_433 net754 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_444 net1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdadda_fa_3_24_3 pp_row24_14 c$1052 s$1055 VGND VGND VPWR VPWR c$2036 s$2037 sky130_fd_sc_hd__fa_1
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_455 net1588 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_91_0 c$3756 c$3758 s$3761 VGND VGND VPWR VPWR c$4078 s$4079 sky130_fd_sc_hd__fa_1
XFILLER_12_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_929 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1430_ clknet_leaf_63_clk booth_b28_m6 VGND VGND VPWR VPWR pp_row34_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_123_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1361_ clknet_leaf_10_clk booth_b14_m17 VGND VGND VPWR VPWR pp_row31_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_122_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_69_5 s$701 s$703 s$705 VGND VGND VPWR VPWR c$1564 s$1565 sky130_fd_sc_hd__fa_1
X_0312_ clknet_leaf_202_clk booth_b60_m13 VGND VGND VPWR VPWR pp_row73_26 sky130_fd_sc_hd__dfxtp_1
X_1292_ clknet_leaf_3_clk booth_b22_m5 VGND VGND VPWR VPWR pp_row27_11 sky130_fd_sc_hd__dfxtp_1
X_0243_ clknet_leaf_153_clk booth_b58_m13 VGND VGND VPWR VPWR pp_row71_26 sky130_fd_sc_hd__dfxtp_1
Xinput180 c[30] VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_1
Xinput191 c[40] VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_1
X_0174_ clknet_leaf_101_clk booth_b56_m13 VGND VGND VPWR VPWR pp_row69_26 sky130_fd_sc_hd__dfxtp_1
Xdadda_ha_0_78_0_1915 VGND VGND VPWR VPWR net1915 dadda_ha_0_78_0_1915/LO sky130_fd_sc_hd__conb_1
XFILLER_93_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$590 net1146 net409 net1138 net675 VGND VGND VPWR VPWR t$4707 sky130_fd_sc_hd__a22o_1
XFILLER_189_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1628_ clknet_leaf_121_clk booth_b64_m41 VGND VGND VPWR VPWR pp_row105_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_154_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1559_ clknet_leaf_7_clk booth_b16_m24 VGND VGND VPWR VPWR pp_row40_8 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_71_5 pp_row71_27 pp_row71_28 pp_row71_29 VGND VGND VPWR VPWR c$736 s$737
+ sky130_fd_sc_hd__fa_1
XFILLER_8_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_64_4 pp_row64_30 pp_row64_31 pp_row64_32 VGND VGND VPWR VPWR c$608 s$609
+ sky130_fd_sc_hd__fa_1
XFILLER_101_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_57_3 pp_row57_17 pp_row57_18 pp_row57_19 VGND VGND VPWR VPWR c$480 s$481
+ sky130_fd_sc_hd__fa_1
Xdadda_fa_4_34_2 s$2113 s$2115 s$2117 VGND VGND VPWR VPWR c$2898 s$2899 sky130_fd_sc_hd__fa_1
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_27_1 c$2050 c$2052 s$2055 VGND VGND VPWR VPWR c$2854 s$2855 sky130_fd_sc_hd__fa_1
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4305 net1077 net419 net1069 net701 VGND VGND VPWR VPWR t$6605 sky130_fd_sc_hd__a22o_1
XFILLER_77_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout870 net874 VGND VGND VPWR VPWR net870 sky130_fd_sc_hd__buf_6
XU$$4316 t$6610 net1259 VGND VGND VPWR VPWR booth_b62_m31 sky130_fd_sc_hd__xor2_1
XU$$4327 net971 net424 net963 net706 VGND VGND VPWR VPWR t$6616 sky130_fd_sc_hd__a22o_1
Xfanout881 net882 VGND VGND VPWR VPWR net881 sky130_fd_sc_hd__clkbuf_4
XFILLER_19_913 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4338 t$6621 net1262 VGND VGND VPWR VPWR booth_b62_m42 sky130_fd_sc_hd__xor2_1
Xfanout892 net895 VGND VGND VPWR VPWR net892 sky130_fd_sc_hd__buf_4
XFILLER_77_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3604 net1151 net479 net1142 net752 VGND VGND VPWR VPWR t$6247 sky130_fd_sc_hd__a22o_1
XU$$4349 net1702 net420 net1692 net702 VGND VGND VPWR VPWR t$6627 sky130_fd_sc_hd__a22o_1
XFILLER_18_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3615 t$6252 net1319 VGND VGND VPWR VPWR booth_b52_m23 sky130_fd_sc_hd__xor2_1
Xdadda_ha_3_16_1 pp_row16_3 pp_row16_4 VGND VGND VPWR VPWR c$1980 s$1981 sky130_fd_sc_hd__ha_1
XU$$3626 net1052 net477 net1044 net750 VGND VGND VPWR VPWR t$6258 sky130_fd_sc_hd__a22o_1
XTAP_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3637 t$6263 net1323 VGND VGND VPWR VPWR booth_b52_m34 sky130_fd_sc_hd__xor2_1
XTAP_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2903 net1500 net523 net1225 net796 VGND VGND VPWR VPWR t$5889 sky130_fd_sc_hd__a22o_1
XU$$3648 net945 net482 net929 net755 VGND VGND VPWR VPWR t$6269 sky130_fd_sc_hd__a22o_1
XU$$3659 t$6274 net1326 VGND VGND VPWR VPWR booth_b52_m45 sky130_fd_sc_hd__xor2_1
XU$$2914 t$5894 net1375 VGND VGND VPWR VPWR booth_b42_m15 sky130_fd_sc_hd__xor2_1
XTAP_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2925 net1120 net522 net1111 net795 VGND VGND VPWR VPWR t$5900 sky130_fd_sc_hd__a22o_1
XFILLER_93_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2936 t$5905 net1373 VGND VGND VPWR VPWR booth_b42_m26 sky130_fd_sc_hd__xor2_1
XTAP_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_193_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_193_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_18_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2947 net1022 net519 net1005 net792 VGND VGND VPWR VPWR t$5911 sky130_fd_sc_hd__a22o_1
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_22_0 pp_row22_2 pp_row22_3 pp_row22_4 VGND VGND VPWR VPWR c$2014 s$2015
+ sky130_fd_sc_hd__fa_1
XANTENNA_230 net1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2958 t$5916 net1370 VGND VGND VPWR VPWR booth_b42_m37 sky130_fd_sc_hd__xor2_1
XANTENNA_241 net1522 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2969 net1740 net521 net1732 net794 VGND VGND VPWR VPWR t$5922 sky130_fd_sc_hd__a22o_1
XANTENNA_252 net1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_263 net1723 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_274 net1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_285 s$4217 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_296 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0930_ clknet_leaf_111_clk booth_b48_m49 VGND VGND VPWR VPWR pp_row97_8 sky130_fd_sc_hd__dfxtp_1
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0861_ clknet_leaf_102_clk booth_b32_m62 VGND VGND VPWR VPWR pp_row94_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_146_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0792_ clknet_leaf_93_clk notsign$5384 VGND VGND VPWR VPWR pp_row91_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_173_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_873 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_81_4 s$909 s$911 s$913 VGND VGND VPWR VPWR c$1706 s$1707 sky130_fd_sc_hd__fa_1
X_2462_ clknet_leaf_95_clk booth_b34_m34 VGND VGND VPWR VPWR pp_row68_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_5_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_898 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1413_ clknet_leaf_244_clk net183 VGND VGND VPWR VPWR pp_row33_17 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_74_3 c$778 s$781 s$783 VGND VGND VPWR VPWR c$1620 s$1621 sky130_fd_sc_hd__fa_1
XFILLER_130_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2393_ clknet_leaf_96_clk booth_b40_m26 VGND VGND VPWR VPWR pp_row66_20 sky130_fd_sc_hd__dfxtp_1
XFILLER_111_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1344_ clknet_leaf_3_clk booth_b20_m10 VGND VGND VPWR VPWR pp_row30_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_96_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_67_2 c$646 c$648 c$650 VGND VGND VPWR VPWR c$1534 s$1535 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$909 final_adder.$signal$1194 final_adder.g_new$987 final_adder.$signal$210
+ VGND VGND VPWR VPWR final_adder.g_new$1037 sky130_fd_sc_hd__a21o_1
Xdadda_fa_5_44_1 s$2955 s$2957 s$2959 VGND VGND VPWR VPWR c$3574 s$3575 sky130_fd_sc_hd__fa_1
X_1275_ clknet_leaf_11_clk booth_b24_m2 VGND VGND VPWR VPWR pp_row26_12 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_37_0 c$2906 c$2908 c$2910 VGND VGND VPWR VPWR c$3544 s$3545 sky130_fd_sc_hd__fa_1
XFILLER_114_1080 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0226_ clknet_leaf_208_clk booth_b26_m45 VGND VGND VPWR VPWR pp_row71_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_64_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_184_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_184_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_64_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_111_0 c$3350 c$3352 c$3354 VGND VGND VPWR VPWR c$3840 s$3841 sky130_fd_sc_hd__fa_1
XFILLER_118_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1109 net1110 VGND VGND VPWR VPWR net1109 sky130_fd_sc_hd__buf_4
XFILLER_102_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_62_1 pp_row62_20 pp_row62_21 pp_row62_22 VGND VGND VPWR VPWR c$566 s$567
+ sky130_fd_sc_hd__fa_1
XFILLER_86_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_55_0 pp_row55_5 pp_row55_6 pp_row55_7 VGND VGND VPWR VPWR c$438 s$439
+ sky130_fd_sc_hd__fa_2
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_175_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_175_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1509 net1481 VGND VGND VPWR VPWR notblock$5175\[2\] sky130_fd_sc_hd__inv_1
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_818 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_91_3 s$1823 s$1825 s$1827 VGND VGND VPWR VPWR c$2572 s$2573 sky130_fd_sc_hd__fa_1
XFILLER_124_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_84_2 c$1732 s$1735 s$1737 VGND VGND VPWR VPWR c$2514 s$2515 sky130_fd_sc_hd__fa_1
XFILLER_136_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_864 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_77_1 c$1642 c$1644 c$1646 VGND VGND VPWR VPWR c$2456 s$2457 sky130_fd_sc_hd__fa_1
XFILLER_2_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_54_0 c$3608 c$3610 s$3613 VGND VGND VPWR VPWR c$4004 s$4005 sky130_fd_sc_hd__fa_1
XFILLER_33_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1610 net1611 VGND VGND VPWR VPWR net1610 sky130_fd_sc_hd__clkbuf_4
XFILLER_2_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1621 net1628 VGND VGND VPWR VPWR net1621 sky130_fd_sc_hd__buf_4
Xfanout1632 net113 VGND VGND VPWR VPWR net1632 sky130_fd_sc_hd__clkbuf_4
Xfanout1643 net1645 VGND VGND VPWR VPWR net1643 sky130_fd_sc_hd__buf_4
Xfanout1654 net1656 VGND VGND VPWR VPWR net1654 sky130_fd_sc_hd__buf_4
XU$$4102 t$6500 net1288 VGND VGND VPWR VPWR booth_b58_m61 sky130_fd_sc_hd__xor2_1
Xfanout1665 net1666 VGND VGND VPWR VPWR net1665 sky130_fd_sc_hd__clkbuf_4
XU$$4113 net1265 notblock$6505\[1\] VGND VGND VPWR VPWR t$6506 sky130_fd_sc_hd__and2_1
XU$$4124 net938 net438 net1677 net720 VGND VGND VPWR VPWR t$6513 sky130_fd_sc_hd__a22o_1
Xfanout1676 net1678 VGND VGND VPWR VPWR net1676 sky130_fd_sc_hd__buf_4
XFILLER_92_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4135 t$6518 net1269 VGND VGND VPWR VPWR booth_b60_m9 sky130_fd_sc_hd__xor2_1
Xfanout1687 net1689 VGND VGND VPWR VPWR net1687 sky130_fd_sc_hd__buf_4
XU$$3401 t$6142 net1346 VGND VGND VPWR VPWR booth_b48_m53 sky130_fd_sc_hd__xor2_1
Xfanout1698 net106 VGND VGND VPWR VPWR net1698 sky130_fd_sc_hd__buf_6
XU$$4146 net1177 net434 net1168 net716 VGND VGND VPWR VPWR t$6524 sky130_fd_sc_hd__a22o_1
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4157 t$6529 net1267 VGND VGND VPWR VPWR booth_b60_m20 sky130_fd_sc_hd__xor2_1
XU$$3412 net1591 net495 net1583 net768 VGND VGND VPWR VPWR t$6148 sky130_fd_sc_hd__a22o_1
X_1060_ clknet_leaf_120_clk booth_b48_m54 VGND VGND VPWR VPWR pp_row102_6 sky130_fd_sc_hd__dfxtp_1
XU$$4168 net1077 net436 net1069 net718 VGND VGND VPWR VPWR t$6535 sky130_fd_sc_hd__a22o_1
XU$$3423 t$6153 net1345 VGND VGND VPWR VPWR booth_b48_m64 sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_113_2 c$2736 s$2739 s$2741 VGND VGND VPWR VPWR c$3372 s$3373 sky130_fd_sc_hd__fa_1
XU$$4179 t$6540 net1269 VGND VGND VPWR VPWR booth_b60_m31 sky130_fd_sc_hd__xor2_1
XU$$3434 t$6160 net1329 VGND VGND VPWR VPWR booth_b50_m1 sky130_fd_sc_hd__xor2_1
XFILLER_93_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2700 t$5784 net1396 VGND VGND VPWR VPWR booth_b38_m45 sky130_fd_sc_hd__xor2_1
XFILLER_20_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3445 net1525 net492 net1517 net765 VGND VGND VPWR VPWR t$6166 sky130_fd_sc_hd__a22o_1
XU$$2711 net1656 net546 net1648 net819 VGND VGND VPWR VPWR t$5790 sky130_fd_sc_hd__a22o_1
XU$$3456 t$6171 net1332 VGND VGND VPWR VPWR booth_b50_m12 sky130_fd_sc_hd__xor2_1
XTAP_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3467 net1153 net488 net1145 net761 VGND VGND VPWR VPWR t$6177 sky130_fd_sc_hd__a22o_1
XU$$2722 t$5795 net1400 VGND VGND VPWR VPWR booth_b38_m56 sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_106_1 c$2682 c$2684 s$2687 VGND VGND VPWR VPWR c$3328 s$3329 sky130_fd_sc_hd__fa_1
XU$$2733 net1550 net548 net1542 net821 VGND VGND VPWR VPWR t$5801 sky130_fd_sc_hd__a22o_1
XU$$3478 t$6182 net1329 VGND VGND VPWR VPWR booth_b50_m23 sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_166_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_166_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2744 notblock$5805\[2\] net35 net1398 t$5806 notblock$5805\[0\] VGND VGND VPWR
+ VPWR sel_0$5807 sky130_fd_sc_hd__a32o_1
XU$$3489 net1051 net485 net1043 net758 VGND VGND VPWR VPWR t$6188 sky130_fd_sc_hd__a22o_1
XTAP_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2755 t$5813 net1376 VGND VGND VPWR VPWR booth_b40_m4 sky130_fd_sc_hd__xor2_1
XTAP_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2766 net1500 net539 net1225 net812 VGND VGND VPWR VPWR t$5819 sky130_fd_sc_hd__a22o_1
XFILLER_2_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2777 t$5824 net1381 VGND VGND VPWR VPWR booth_b40_m15 sky130_fd_sc_hd__xor2_1
XU$$2788 net1120 net536 net1111 net809 VGND VGND VPWR VPWR t$5830 sky130_fd_sc_hd__a22o_1
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2799 t$5835 net1381 VGND VGND VPWR VPWR booth_b40_m26 sky130_fd_sc_hd__xor2_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1962_ clknet_leaf_64_clk booth_b26_m28 VGND VGND VPWR VPWR pp_row54_13 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_7_127_0 c$3898 c$4148 s$4151 VGND VGND VPWR VPWR dadda_fa_7_127_0/COUT s$4407
+ sky130_fd_sc_hd__fa_1
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0913_ clknet_leaf_104_clk booth_b52_m44 VGND VGND VPWR VPWR pp_row96_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_147_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1893_ clknet_leaf_64_clk booth_b18_m34 VGND VGND VPWR VPWR pp_row52_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0844_ clknet_leaf_129_clk booth_b64_m55 VGND VGND VPWR VPWR pp_row119_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_128_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0775_ clknet_leaf_141_clk booth_b38_m52 VGND VGND VPWR VPWR pp_row90_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_115_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2445_ clknet_leaf_89_clk booth_b4_m64 VGND VGND VPWR VPWR pp_row68_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_64_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_72_0 s$179 c$726 c$728 VGND VGND VPWR VPWR c$1590 s$1591 sky130_fd_sc_hd__fa_1
XFILLER_25_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2376_ clknet_leaf_85_clk booth_b12_m54 VGND VGND VPWR VPWR pp_row66_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$706 final_adder.p_new$730 final_adder.p_new$714 VGND VGND VPWR VPWR
+ final_adder.p_new$834 sky130_fd_sc_hd__and2_1
XFILLER_111_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$717 final_adder.p_new$724 final_adder.g_new$741 final_adder.g_new$725
+ VGND VGND VPWR VPWR final_adder.g_new$845 sky130_fd_sc_hd__a21o_1
X_1327_ clknet_leaf_184_clk net133 VGND VGND VPWR VPWR pp_row103_14 sky130_fd_sc_hd__dfxtp_2
XFILLER_68_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1258_ clknet_leaf_9_clk booth_b22_m3 VGND VGND VPWR VPWR pp_row25_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_56_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_157_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_157_clk
+ sky130_fd_sc_hd__clkbuf_16
X_0209_ clknet_leaf_152_clk booth_b58_m12 VGND VGND VPWR VPWR pp_row70_27 sky130_fd_sc_hd__dfxtp_1
XFILLER_52_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1189_ clknet_leaf_49_clk booth_b4_m17 VGND VGND VPWR VPWR pp_row21_2 sky130_fd_sc_hd__dfxtp_1
XU$$3990 t$6444 net1282 VGND VGND VPWR VPWR booth_b58_m5 sky130_fd_sc_hd__xor2_1
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_94_1 c$2586 c$2588 s$2591 VGND VGND VPWR VPWR c$3256 s$3257 sky130_fd_sc_hd__fa_1
XFILLER_137_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_71_0 s$3683 c$4036 s$4039 VGND VGND VPWR VPWR c$4294 s$4295 sky130_fd_sc_hd__fa_1
XFILLER_146_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_87_0 s$1781 c$2526 c$2528 VGND VGND VPWR VPWR c$3212 s$3213 sky130_fd_sc_hd__fa_1
Xdadda_fa_3_108_3 pp_row108_11 pp_row108_12 c$1970 VGND VGND VPWR VPWR c$2708 s$2709
+ sky130_fd_sc_hd__fa_1
XFILLER_165_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput270 net270 VGND VGND VPWR VPWR o[111] sky130_fd_sc_hd__buf_2
Xoutput281 net281 VGND VGND VPWR VPWR o[121] sky130_fd_sc_hd__buf_2
Xoutput292 net292 VGND VGND VPWR VPWR o[16] sky130_fd_sc_hd__buf_2
XU$$2061_1771 VGND VGND VPWR VPWR U$$2061_1771/HI net1771 sky130_fd_sc_hd__conb_1
XFILLER_0_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3148_1788 VGND VGND VPWR VPWR U$$3148_1788/HI net1788 sky130_fd_sc_hd__conb_1
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2007 t$5430 net1455 VGND VGND VPWR VPWR booth_b28_m41 sky130_fd_sc_hd__xor2_1
XU$$2018 net1704 net589 net1696 net862 VGND VGND VPWR VPWR t$5436 sky130_fd_sc_hd__a22o_1
XU$$2029 t$5441 net1453 VGND VGND VPWR VPWR booth_b28_m52 sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_148_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_148_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_28_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1306 t$5072 net1666 VGND VGND VPWR VPWR booth_b18_m33 sky130_fd_sc_hd__xor2_1
XFILLER_74_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1317 net955 net638 net944 net911 VGND VGND VPWR VPWR t$5078 sky130_fd_sc_hd__a22o_1
XU$$1328 t$5083 net1663 VGND VGND VPWR VPWR booth_b18_m44 sky130_fd_sc_hd__xor2_1
XU$$1339 net1682 net642 net1657 net915 VGND VGND VPWR VPWR t$5089 sky130_fd_sc_hd__a22o_1
XFILLER_128_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_1068 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_935 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0560_ clknet_leaf_186_clk booth_b18_m64 VGND VGND VPWR VPWR pp_row82_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_125_876 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0491_ clknet_leaf_159_clk booth_b48_m31 VGND VGND VPWR VPWR pp_row79_17 sky130_fd_sc_hd__dfxtp_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2230_ clknet_leaf_233_clk booth_b14_m48 VGND VGND VPWR VPWR pp_row62_7 sky130_fd_sc_hd__dfxtp_1
Xfanout1440 net1443 VGND VGND VPWR VPWR net1440 sky130_fd_sc_hd__buf_8
XFILLER_39_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2161_ clknet_leaf_214_clk booth_b20_m40 VGND VGND VPWR VPWR pp_row60_10 sky130_fd_sc_hd__dfxtp_1
Xfanout1451 net1452 VGND VGND VPWR VPWR net1451 sky130_fd_sc_hd__buf_6
Xfanout1462 net20 VGND VGND VPWR VPWR net1462 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_51_5 s$377 s$379 s$381 VGND VGND VPWR VPWR c$1348 s$1349 sky130_fd_sc_hd__fa_2
Xfanout1473 net1474 VGND VGND VPWR VPWR net1473 sky130_fd_sc_hd__buf_6
Xfanout1484 net16 VGND VGND VPWR VPWR net1484 sky130_fd_sc_hd__buf_6
X_1112_ clknet_leaf_248_clk net162 VGND VGND VPWR VPWR pp_row14_9 sky130_fd_sc_hd__dfxtp_2
Xfanout1495 net1498 VGND VGND VPWR VPWR net1495 sky130_fd_sc_hd__buf_2
XFILLER_66_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_44_4 c$262 s$265 s$267 VGND VGND VPWR VPWR c$1262 s$1263 sky130_fd_sc_hd__fa_1
X_2092_ clknet_leaf_149_clk booth_b22_m36 VGND VGND VPWR VPWR pp_row58_11 sky130_fd_sc_hd__dfxtp_1
XU$$3220 t$6050 net1349 VGND VGND VPWR VPWR booth_b46_m31 sky130_fd_sc_hd__xor2_1
Xdadda_ha_6_3_0 pp_row3_0 pp_row3_1 VGND VGND VPWR VPWR c$3902 s$3903 sky130_fd_sc_hd__ha_1
XFILLER_24_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3231 net966 net503 net959 net776 VGND VGND VPWR VPWR t$6056 sky130_fd_sc_hd__a22o_1
XU$$3242 t$6061 net1350 VGND VGND VPWR VPWR booth_b46_m42 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$13 c$4176 s$4179 VGND VGND VPWR VPWR final_adder.$signal$28 final_adder.$signal$1103
+ sky130_fd_sc_hd__ha_1
XU$$3253 net1700 net507 net1693 net780 VGND VGND VPWR VPWR t$6067 sky130_fd_sc_hd__a22o_1
X_1043_ clknet_leaf_56_clk booth_b6_m0 VGND VGND VPWR VPWR pp_row6_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_94_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$24 c$4198 s$4201 VGND VGND VPWR VPWR final_adder.$signal$50 final_adder.$signal$1114
+ sky130_fd_sc_hd__ha_2
XU$$3264 t$6072 net1355 VGND VGND VPWR VPWR booth_b46_m53 sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_37_3 pp_row37_14 pp_row37_15 pp_row37_16 VGND VGND VPWR VPWR c$1176 s$1177
+ sky130_fd_sc_hd__fa_1
Xclkbuf_leaf_139_clk clknet_5_25__leaf_clk VGND VGND VPWR VPWR clknet_leaf_139_clk
+ sky130_fd_sc_hd__clkbuf_16
Xfinal_adder.U$$35 c$4220 s$4223 VGND VGND VPWR VPWR final_adder.$signal$72 final_adder.$signal$1125
+ sky130_fd_sc_hd__ha_1
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$46 c$4242 s$4245 VGND VGND VPWR VPWR final_adder.$signal$94 final_adder.$signal$1136
+ sky130_fd_sc_hd__ha_1
XU$$2530 net1050 net554 net1042 net827 VGND VGND VPWR VPWR t$5698 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$57 c$4264 s$4267 VGND VGND VPWR VPWR final_adder.$signal$116 final_adder.$signal$1147
+ sky130_fd_sc_hd__ha_1
XU$$3275 net1593 net507 net1585 net780 VGND VGND VPWR VPWR t$6078 sky130_fd_sc_hd__a22o_1
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2541 t$5703 net1409 VGND VGND VPWR VPWR booth_b36_m34 sky130_fd_sc_hd__xor2_1
XU$$3286 t$6083 net1350 VGND VGND VPWR VPWR booth_b46_m64 sky130_fd_sc_hd__xor2_1
XU$$2552 net942 net555 net926 net828 VGND VGND VPWR VPWR t$5709 sky130_fd_sc_hd__a22o_1
XU$$3297 t$6090 net1338 VGND VGND VPWR VPWR booth_b48_m1 sky130_fd_sc_hd__xor2_1
XFILLER_80_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$68 c$4286 s$4289 VGND VGND VPWR VPWR final_adder.$signal$138 final_adder.$signal$1158
+ sky130_fd_sc_hd__ha_1
XFILLER_146_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2563 t$5714 net1408 VGND VGND VPWR VPWR booth_b36_m45 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$79 c$4308 s$4311 VGND VGND VPWR VPWR final_adder.$signal$160 final_adder.$signal$1169
+ sky130_fd_sc_hd__ha_1
XU$$2574 net1655 net556 net1647 net829 VGND VGND VPWR VPWR t$5720 sky130_fd_sc_hd__a22o_1
XU$$1840 t$5345 net1461 VGND VGND VPWR VPWR booth_b26_m26 sky130_fd_sc_hd__xor2_1
XU$$2585 t$5725 net1410 VGND VGND VPWR VPWR booth_b36_m56 sky130_fd_sc_hd__xor2_1
XU$$2596 net1550 net558 net1542 net831 VGND VGND VPWR VPWR t$5731 sky130_fd_sc_hd__a22o_1
XFILLER_146_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1851 net1018 net597 net1001 net870 VGND VGND VPWR VPWR t$5351 sky130_fd_sc_hd__a22o_1
XU$$1862 t$5356 net1459 VGND VGND VPWR VPWR booth_b26_m37 sky130_fd_sc_hd__xor2_1
XU$$1873 net1741 net600 net1733 net873 VGND VGND VPWR VPWR t$5362 sky130_fd_sc_hd__a22o_1
XU$$1884 t$5367 net1459 VGND VGND VPWR VPWR booth_b26_m48 sky130_fd_sc_hd__xor2_1
XFILLER_166_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1895 net1631 net598 net1622 net871 VGND VGND VPWR VPWR t$5373 sky130_fd_sc_hd__a22o_1
X_1945_ clknet_leaf_231_clk net205 VGND VGND VPWR VPWR pp_row53_27 sky130_fd_sc_hd__dfxtp_4
XFILLER_148_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1876_ clknet_leaf_69_clk booth_b40_m11 VGND VGND VPWR VPWR pp_row51_20 sky130_fd_sc_hd__dfxtp_1
XFILLER_119_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0827_ clknet_leaf_108_clk booth_b50_m42 VGND VGND VPWR VPWR pp_row92_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_116_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1095 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0758_ clknet_leaf_153_clk booth_b48_m41 VGND VGND VPWR VPWR pp_row89_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_115_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0689_ clknet_leaf_168_clk booth_b58_m28 VGND VGND VPWR VPWR pp_row86_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_142_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2428_ clknet_leaf_96_clk booth_b36_m31 VGND VGND VPWR VPWR pp_row67_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_9_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$503 final_adder.p_new$504 final_adder.g_new$509 final_adder.g_new$505
+ VGND VGND VPWR VPWR final_adder.g_new$631 sky130_fd_sc_hd__a21o_4
XFILLER_97_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$514 final_adder.p_new$526 final_adder.p_new$518 VGND VGND VPWR VPWR
+ final_adder.p_new$642 sky130_fd_sc_hd__and2_1
XFILLER_29_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2359_ clknet_leaf_127_clk booth_b52_m59 VGND VGND VPWR VPWR pp_row111_3 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$525 final_adder.p_new$528 final_adder.g_new$537 final_adder.g_new$529
+ VGND VGND VPWR VPWR final_adder.g_new$653 sky130_fd_sc_hd__a21o_1
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$536 final_adder.p_new$548 final_adder.p_new$540 VGND VGND VPWR VPWR
+ final_adder.p_new$664 sky130_fd_sc_hd__and2_1
XFILLER_96_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$547 final_adder.p_new$550 final_adder.g_new$559 final_adder.g_new$551
+ VGND VGND VPWR VPWR final_adder.g_new$675 sky130_fd_sc_hd__a21o_1
XTAP_3829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$558 final_adder.p_new$570 final_adder.p_new$562 VGND VGND VPWR VPWR
+ final_adder.p_new$686 sky130_fd_sc_hd__and2_1
XFILLER_151_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$569 final_adder.p_new$572 final_adder.g_new$581 final_adder.g_new$573
+ VGND VGND VPWR VPWR final_adder.g_new$697 sky130_fd_sc_hd__a21o_1
XFILLER_72_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$408 net1531 net533 net1803 net806 VGND VGND VPWR VPWR t$4613 sky130_fd_sc_hd__a22o_1
XU$$419 net1231 net429 net1127 net711 VGND VGND VPWR VPWR t$4620 sky130_fd_sc_hd__a22o_1
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_607 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_113_1 pp_row113_3 pp_row113_4 pp_row113_5 VGND VGND VPWR VPWR c$2740 s$2741
+ sky130_fd_sc_hd__fa_1
XFILLER_109_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_106_0 pp_row106_5 pp_row106_6 pp_row106_7 VGND VGND VPWR VPWR c$2686 s$2687
+ sky130_fd_sc_hd__fa_1
XFILLER_69_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_900 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_54_3 s$1379 s$1381 s$1383 VGND VGND VPWR VPWR c$2276 s$2277 sky130_fd_sc_hd__fa_1
XFILLER_134_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_47_2 c$1288 s$1291 s$1293 VGND VGND VPWR VPWR c$2218 s$2219 sky130_fd_sc_hd__fa_1
XFILLER_78_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$920 net1715 net399 net1706 net665 VGND VGND VPWR VPWR t$4875 sky130_fd_sc_hd__a22o_1
XU$$931 t$4880 net1317 VGND VGND VPWR VPWR booth_b12_m51 sky130_fd_sc_hd__xor2_1
XFILLER_16_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$942 net1607 net399 net1599 net665 VGND VGND VPWR VPWR t$4886 sky130_fd_sc_hd__a22o_1
XU$$953 t$4891 net1316 VGND VGND VPWR VPWR booth_b12_m62 sky130_fd_sc_hd__xor2_1
XFILLER_62_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_6_17_0 c$3460 c$3462 s$3465 VGND VGND VPWR VPWR c$3930 s$3931 sky130_fd_sc_hd__fa_1
XU$$964 net6 net1317 VGND VGND VPWR VPWR sel_1$4898 sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_80_0_1896 VGND VGND VPWR VPWR net1896 dadda_fa_1_80_0_1896/LO sky130_fd_sc_hd__conb_1
XU$$1103 t$4969 net1006 VGND VGND VPWR VPWR booth_b16_m0 sky130_fd_sc_hd__xor2_1
XFILLER_62_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1114 net1564 net646 net1523 net919 VGND VGND VPWR VPWR t$4975 sky130_fd_sc_hd__a22o_1
XFILLER_188_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$975 net1676 net389 net1564 net655 VGND VGND VPWR VPWR t$4904 sky130_fd_sc_hd__a22o_1
XU$$1125 t$4980 net1006 VGND VGND VPWR VPWR booth_b16_m11 sky130_fd_sc_hd__xor2_1
XU$$986 t$4909 net1183 VGND VGND VPWR VPWR booth_b14_m10 sky130_fd_sc_hd__xor2_1
XU$$997 net1164 net385 net1155 net651 VGND VGND VPWR VPWR t$4915 sky130_fd_sc_hd__a22o_1
XU$$1136 net1161 net646 net1149 net919 VGND VGND VPWR VPWR t$4986 sky130_fd_sc_hd__a22o_1
XU$$1147 t$4991 net1009 VGND VGND VPWR VPWR booth_b16_m22 sky130_fd_sc_hd__xor2_1
XU$$1158 net1055 net647 net1047 net920 VGND VGND VPWR VPWR t$4997 sky130_fd_sc_hd__a22o_1
XFILLER_188_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1169 t$5002 net1007 VGND VGND VPWR VPWR booth_b16_m33 sky130_fd_sc_hd__xor2_1
XFILLER_188_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_782 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1730_ clknet_leaf_24_clk booth_b40_m6 VGND VGND VPWR VPWR pp_row46_20 sky130_fd_sc_hd__dfxtp_1
XFILLER_156_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1661_ clknet_leaf_124_clk booth_b44_m62 VGND VGND VPWR VPWR pp_row106_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_144_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0612_ clknet_leaf_173_clk booth_b60_m23 VGND VGND VPWR VPWR pp_row83_21 sky130_fd_sc_hd__dfxtp_1
X_1592_ clknet_leaf_5_clk booth_b30_m11 VGND VGND VPWR VPWR pp_row41_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_4_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0543_ clknet_leaf_170_clk booth_b38_m43 VGND VGND VPWR VPWR pp_row81_11 sky130_fd_sc_hd__dfxtp_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0474_ clknet_leaf_193_clk booth_b18_m61 VGND VGND VPWR VPWR pp_row79_2 sky130_fd_sc_hd__dfxtp_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2213_ clknet_leaf_217_clk booth_b48_m13 VGND VGND VPWR VPWR pp_row61_24 sky130_fd_sc_hd__dfxtp_1
XFILLER_66_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1270 net1271 VGND VGND VPWR VPWR net1270 sky130_fd_sc_hd__buf_6
XFILLER_61_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1281 net56 VGND VGND VPWR VPWR net1281 sky130_fd_sc_hd__buf_6
Xfanout1292 net1293 VGND VGND VPWR VPWR net1292 sky130_fd_sc_hd__buf_4
X_2144_ clknet_leaf_31_clk booth_b52_m7 VGND VGND VPWR VPWR pp_row59_26 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_42_1 pp_row42_17 pp_row42_18 pp_row42_19 VGND VGND VPWR VPWR c$1232 s$1233
+ sky130_fd_sc_hd__fa_1
XFILLER_82_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3050 net1176 net511 net1167 net784 VGND VGND VPWR VPWR t$5964 sky130_fd_sc_hd__a22o_1
X_2075_ clknet_leaf_32_clk booth_b50_m7 VGND VGND VPWR VPWR pp_row57_25 sky130_fd_sc_hd__dfxtp_1
XU$$3061 t$5969 net1362 VGND VGND VPWR VPWR booth_b44_m20 sky130_fd_sc_hd__xor2_1
XFILLER_35_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_35_0 pp_row35_2 pp_row35_3 pp_row35_4 VGND VGND VPWR VPWR c$1146 s$1147
+ sky130_fd_sc_hd__fa_1
XU$$3072 net1076 net513 net1068 net786 VGND VGND VPWR VPWR t$5975 sky130_fd_sc_hd__a22o_1
XU$$3083 t$5980 net1359 VGND VGND VPWR VPWR booth_b44_m31 sky130_fd_sc_hd__xor2_1
X_1026_ clknet_leaf_61_clk booth_b0_m3 VGND VGND VPWR VPWR pp_row3_0 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_5_22__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_5_22__leaf_clk sky130_fd_sc_hd__clkbuf_16
XU$$3094 net967 net512 net958 net785 VGND VGND VPWR VPWR t$5986 sky130_fd_sc_hd__a22o_1
XU$$2360 t$5611 net1420 VGND VGND VPWR VPWR booth_b34_m12 sky130_fd_sc_hd__xor2_1
XU$$2371 net1150 net563 net1144 net836 VGND VGND VPWR VPWR t$5617 sky130_fd_sc_hd__a22o_1
XFILLER_22_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2382 t$5622 net1421 VGND VGND VPWR VPWR booth_b34_m23 sky130_fd_sc_hd__xor2_1
XU$$2393 net1051 net562 net1043 net835 VGND VGND VPWR VPWR t$5628 sky130_fd_sc_hd__a22o_1
XFILLER_34_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1670 net1500 net605 net1225 net878 VGND VGND VPWR VPWR t$5259 sky130_fd_sc_hd__a22o_1
XU$$1681 t$5264 net1467 VGND VGND VPWR VPWR booth_b24_m15 sky130_fd_sc_hd__xor2_1
XU$$1692 net1116 net603 net1106 net876 VGND VGND VPWR VPWR t$5270 sky130_fd_sc_hd__a22o_1
X_1928_ clknet_leaf_69_clk booth_b22_m31 VGND VGND VPWR VPWR pp_row53_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1859_ clknet_leaf_79_clk booth_b10_m41 VGND VGND VPWR VPWR pp_row51_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1001 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_87_3 pp_row87_9 pp_row87_10 pp_row87_11 VGND VGND VPWR VPWR c$996 s$997
+ sky130_fd_sc_hd__fa_1
XFILLER_104_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_64_2 s$2353 s$2355 s$2357 VGND VGND VPWR VPWR c$3078 s$3079 sky130_fd_sc_hd__fa_1
XFILLER_162_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_57_1 c$2290 c$2292 s$2295 VGND VGND VPWR VPWR c$3034 s$3035 sky130_fd_sc_hd__fa_1
XTAP_4305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$300 final_adder.p_new$302 final_adder.p_new$300 VGND VGND VPWR VPWR
+ final_adder.p_new$428 sky130_fd_sc_hd__and2_1
XTAP_4327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_34_0 s$3535 c$3962 s$3965 VGND VGND VPWR VPWR c$4220 s$4221 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$311 final_adder.p_new$310 final_adder.g_new$313 final_adder.g_new$311
+ VGND VGND VPWR VPWR final_adder.g_new$439 sky130_fd_sc_hd__a21o_1
XTAP_4338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$322 final_adder.p_new$324 final_adder.p_new$322 VGND VGND VPWR VPWR
+ final_adder.p_new$450 sky130_fd_sc_hd__and2_1
XTAP_4349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$333 final_adder.p_new$332 final_adder.g_new$335 final_adder.g_new$333
+ VGND VGND VPWR VPWR final_adder.g_new$461 sky130_fd_sc_hd__a21o_1
XTAP_3615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$344 final_adder.p_new$346 final_adder.p_new$344 VGND VGND VPWR VPWR
+ final_adder.p_new$472 sky130_fd_sc_hd__and2_1
XFILLER_45_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$355 final_adder.p_new$354 final_adder.g_new$357 final_adder.g_new$355
+ VGND VGND VPWR VPWR final_adder.g_new$483 sky130_fd_sc_hd__a21o_1
XTAP_3637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$205 net1025 net623 net1017 net896 VGND VGND VPWR VPWR t$4510 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$366 final_adder.p_new$368 final_adder.p_new$366 VGND VGND VPWR VPWR
+ final_adder.p_new$494 sky130_fd_sc_hd__and2_1
XTAP_3648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$377 final_adder.p_new$376 final_adder.g_new$379 final_adder.g_new$377
+ VGND VGND VPWR VPWR final_adder.g_new$505 sky130_fd_sc_hd__a21o_1
XU$$216 t$4515 net1386 VGND VGND VPWR VPWR booth_b2_m36 sky130_fd_sc_hd__xor2_1
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$388 final_adder.p_new$394 final_adder.p_new$390 VGND VGND VPWR VPWR
+ final_adder.p_new$516 sky130_fd_sc_hd__and2_1
XU$$227 net1745 net622 net1737 net895 VGND VGND VPWR VPWR t$4521 sky130_fd_sc_hd__a22o_1
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$238 t$4526 net1392 VGND VGND VPWR VPWR booth_b2_m47 sky130_fd_sc_hd__xor2_1
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$399 final_adder.p_new$400 final_adder.g_new$405 final_adder.g_new$401
+ VGND VGND VPWR VPWR final_adder.g_new$527 sky130_fd_sc_hd__a21o_1
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$249 net1642 net626 net1637 net899 VGND VGND VPWR VPWR t$4532 sky130_fd_sc_hd__a22o_1
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4401_1821 VGND VGND VPWR VPWR U$$4401_1821/HI net1821 sky130_fd_sc_hd__conb_1
XFILLER_154_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_1011 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_0_75_1 pp_row75_3 pp_row75_4 pp_row75_5 VGND VGND VPWR VPWR c$194 s$195
+ sky130_fd_sc_hd__fa_1
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_52_0 s$401 c$1338 c$1340 VGND VGND VPWR VPWR c$2254 s$2255 sky130_fd_sc_hd__fa_2
Xdadda_fa_0_68_0 net1891 pp_row68_1 pp_row68_2 VGND VGND VPWR VPWR c$132 s$133 sky130_fd_sc_hd__fa_1
XFILLER_36_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0190_ clknet_leaf_148_clk booth_b22_m48 VGND VGND VPWR VPWR pp_row70_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_152_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$750 t$4788 net1415 VGND VGND VPWR VPWR booth_b10_m29 sky130_fd_sc_hd__xor2_1
XU$$761 net986 net406 net981 net672 VGND VGND VPWR VPWR t$4794 sky130_fd_sc_hd__a22o_1
XFILLER_32_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$772 t$4799 net1418 VGND VGND VPWR VPWR booth_b10_m40 sky130_fd_sc_hd__xor2_1
XU$$783 net1716 net407 net1707 net673 VGND VGND VPWR VPWR t$4805 sky130_fd_sc_hd__a22o_1
XU$$794 t$4810 net1418 VGND VGND VPWR VPWR booth_b10_m51 sky130_fd_sc_hd__xor2_1
XFILLER_56_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_70_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_70_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_17_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1713_ clknet_leaf_237_clk booth_b12_m34 VGND VGND VPWR VPWR pp_row46_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_117_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_97_2 pp_row97_6 pp_row97_7 pp_row97_8 VGND VGND VPWR VPWR c$1894 s$1895
+ sky130_fd_sc_hd__fa_1
X_1644_ clknet_leaf_6_clk booth_b30_m13 VGND VGND VPWR VPWR pp_row43_15 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_74_1 s$3135 s$3137 s$3139 VGND VGND VPWR VPWR c$3694 s$3695 sky130_fd_sc_hd__fa_2
XFILLER_126_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1575_ clknet_leaf_244_clk net191 VGND VGND VPWR VPWR pp_row40_22 sky130_fd_sc_hd__dfxtp_1
XFILLER_98_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_67_0 c$3086 c$3088 c$3090 VGND VGND VPWR VPWR c$3664 s$3665 sky130_fd_sc_hd__fa_1
Xfanout507 net508 VGND VGND VPWR VPWR net507 sky130_fd_sc_hd__buf_4
Xfanout518 sel_0$5947 VGND VGND VPWR VPWR net518 sky130_fd_sc_hd__buf_4
XFILLER_59_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout529 net530 VGND VGND VPWR VPWR net529 sky130_fd_sc_hd__buf_4
X_0526_ clknet_leaf_162_clk booth_b58_m22 VGND VGND VPWR VPWR pp_row80_22 sky130_fd_sc_hd__dfxtp_1
XFILLER_98_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_985 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_66_8 s$113 s$115 s$117 VGND VGND VPWR VPWR c$652 s$653 sky130_fd_sc_hd__fa_1
X_0457_ clknet_leaf_157_clk booth_b40_m38 VGND VGND VPWR VPWR pp_row78_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_59_7 c$26 c$28 c$30 VGND VGND VPWR VPWR c$524 s$525 sky130_fd_sc_hd__fa_1
XFILLER_132_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0388_ clknet_leaf_127_clk booth_b60_m54 VGND VGND VPWR VPWR pp_row114_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2127_ clknet_leaf_129_clk booth_b54_m55 VGND VGND VPWR VPWR pp_row109_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_148_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2058_ clknet_leaf_42_clk booth_b22_m35 VGND VGND VPWR VPWR pp_row57_11 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_6_6_0 pp_row6_5 c$3418 s$3421 VGND VGND VPWR VPWR c$3908 s$3909 sky130_fd_sc_hd__fa_1
XFILLER_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1009_ clknet_leaf_119_clk booth_b58_m43 VGND VGND VPWR VPWR pp_row101_11 sky130_fd_sc_hd__dfxtp_1
XU$$2190 t$5523 net1447 VGND VGND VPWR VPWR booth_b30_m64 sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_61_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_61_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_23_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3294_1791 VGND VGND VPWR VPWR U$$3294_1791/HI net1791 sky130_fd_sc_hd__conb_1
XFILLER_182_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_92_1 pp_row92_3 pp_row92_4 pp_row92_5 VGND VGND VPWR VPWR c$1034 s$1035
+ sky130_fd_sc_hd__fa_1
XFILLER_123_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_85_0 pp_row85_0 pp_row85_1 pp_row85_2 VGND VGND VPWR VPWR c$966 s$967
+ sky130_fd_sc_hd__fa_1
XFILLER_132_941 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4431_1836 VGND VGND VPWR VPWR U$$4431_1836/HI net1836 sky130_fd_sc_hd__conb_1
XFILLER_104_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4509 t$6708 net1875 VGND VGND VPWR VPWR booth_b64_m59 sky130_fd_sc_hd__xor2_1
XTAP_4124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3808 t$6350 net1307 VGND VGND VPWR VPWR booth_b54_m51 sky130_fd_sc_hd__xor2_1
XFILLER_18_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$130 final_adder.$signal$1214 final_adder.$signal$1215 VGND VGND VPWR
+ VPWR final_adder.p_new$258 sky130_fd_sc_hd__and2_1
XTAP_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3819 net1608 net473 net1600 net746 VGND VGND VPWR VPWR t$6356 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$141 final_adder.$signal$1205 final_adder.$signal$230 final_adder.$signal$232
+ VGND VGND VPWR VPWR final_adder.g_new$269 sky130_fd_sc_hd__a21o_1
XTAP_4168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$152 final_adder.$signal$1192 final_adder.$signal$1193 VGND VGND VPWR
+ VPWR final_adder.p_new$280 sky130_fd_sc_hd__and2_1
XTAP_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$163 final_adder.$signal$1183 final_adder.$signal$186 final_adder.$signal$188
+ VGND VGND VPWR VPWR final_adder.g_new$291 sky130_fd_sc_hd__a21o_1
XTAP_4179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$174 final_adder.$signal$1170 final_adder.$signal$1171 VGND VGND VPWR
+ VPWR final_adder.p_new$302 sky130_fd_sc_hd__and2_1
XTAP_3456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_401 net1639 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$185 final_adder.$signal$1161 final_adder.$signal$142 final_adder.$signal$144
+ VGND VGND VPWR VPWR final_adder.g_new$313 sky130_fd_sc_hd__a21o_1
XTAP_3467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$196 final_adder.$signal$1148 final_adder.$signal$1149 VGND VGND VPWR
+ VPWR final_adder.p_new$324 sky130_fd_sc_hd__and2_1
XANTENNA_412 net1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_423 net568 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdadda_ha_5_126_0 net1920 pp_row126_1 VGND VGND VPWR VPWR c$3898 s$3899 sky130_fd_sc_hd__ha_1
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_434 net760 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_445 net1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_456 net1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_52_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_52_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_186_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4399_1820 VGND VGND VPWR VPWR U$$4399_1820/HI net1820 sky130_fd_sc_hd__conb_1
XFILLER_40_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_84_0 c$3728 c$3730 s$3733 VGND VGND VPWR VPWR c$4064 s$4065 sky130_fd_sc_hd__fa_1
XFILLER_103_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1360_ clknet_leaf_110_clk booth_b44_m60 VGND VGND VPWR VPWR pp_row104_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_68_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0311_ clknet_leaf_128_clk booth_b64_m49 VGND VGND VPWR VPWR pp_row113_8 sky130_fd_sc_hd__dfxtp_1
X_1291_ clknet_leaf_2_clk booth_b20_m7 VGND VGND VPWR VPWR pp_row27_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_96_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0242_ clknet_leaf_153_clk booth_b56_m15 VGND VGND VPWR VPWR pp_row71_25 sky130_fd_sc_hd__dfxtp_1
Xinput170 c[21] VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_1
Xinput181 c[31] VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$134_1758 VGND VGND VPWR VPWR U$$134_1758/HI net1758 sky130_fd_sc_hd__conb_1
Xinput192 c[41] VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_1
X_0173_ clknet_leaf_101_clk booth_b54_m15 VGND VGND VPWR VPWR pp_row69_25 sky130_fd_sc_hd__dfxtp_1
XTAP_3990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$580 net1207 net413 net1199 net679 VGND VGND VPWR VPWR t$4702 sky130_fd_sc_hd__a22o_1
XU$$591 t$4707 net1235 VGND VGND VPWR VPWR booth_b8_m18 sky130_fd_sc_hd__xor2_1
XFILLER_51_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1000 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_43_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_43_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_189_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1627_ clknet_leaf_221_clk booth_b0_m43 VGND VGND VPWR VPWR pp_row43_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_99_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1558_ clknet_leaf_7_clk booth_b14_m26 VGND VGND VPWR VPWR pp_row40_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_59_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_71_6 pp_row71_30 c$154 c$156 VGND VGND VPWR VPWR c$738 s$739 sky130_fd_sc_hd__fa_1
X_0509_ clknet_leaf_173_clk booth_b28_m52 VGND VGND VPWR VPWR pp_row80_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_98_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_64_5 pp_row64_33 c$72 c$74 VGND VGND VPWR VPWR c$610 s$611 sky130_fd_sc_hd__fa_2
X_1489_ clknet_leaf_43_clk booth_b16_m21 VGND VGND VPWR VPWR pp_row37_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_101_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_57_4 pp_row57_20 pp_row57_21 pp_row57_22 VGND VGND VPWR VPWR c$482 s$483
+ sky130_fd_sc_hd__fa_1
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_27_2 s$2057 s$2059 s$2061 VGND VGND VPWR VPWR c$2856 s$2857 sky130_fd_sc_hd__fa_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_34_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_52_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_579 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_2_108_0_1917 VGND VGND VPWR VPWR net1917 dadda_ha_2_108_0_1917/LO sky130_fd_sc_hd__conb_1
XFILLER_2_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4306 t$6605 net1256 VGND VGND VPWR VPWR booth_b62_m26 sky130_fd_sc_hd__xor2_1
Xfanout860 net861 VGND VGND VPWR VPWR net860 sky130_fd_sc_hd__buf_4
Xfanout871 net873 VGND VGND VPWR VPWR net871 sky130_fd_sc_hd__buf_4
XFILLER_77_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4317 net1021 net422 net1004 net704 VGND VGND VPWR VPWR t$6611 sky130_fd_sc_hd__a22o_1
XFILLER_133_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout882 sel_1$5248 VGND VGND VPWR VPWR net882 sky130_fd_sc_hd__buf_6
XU$$4328 t$6616 net1261 VGND VGND VPWR VPWR booth_b62_m37 sky130_fd_sc_hd__xor2_1
Xfanout893 net895 VGND VGND VPWR VPWR net893 sky130_fd_sc_hd__clkbuf_4
XU$$4339 net1742 net424 net1734 net706 VGND VGND VPWR VPWR t$6622 sky130_fd_sc_hd__a22o_1
XFILLER_19_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3605 t$6247 net1320 VGND VGND VPWR VPWR booth_b52_m18 sky130_fd_sc_hd__xor2_1
XU$$3616 net1094 net476 net1086 net749 VGND VGND VPWR VPWR t$6253 sky130_fd_sc_hd__a22o_1
XU$$3627 t$6258 net1323 VGND VGND VPWR VPWR booth_b52_m29 sky130_fd_sc_hd__xor2_1
XTAP_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3638 net985 net477 net976 net750 VGND VGND VPWR VPWR t$6264 sky130_fd_sc_hd__a22o_1
XTAP_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2904 t$5889 net1372 VGND VGND VPWR VPWR booth_b42_m10 sky130_fd_sc_hd__xor2_1
XTAP_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3649 t$6269 net1326 VGND VGND VPWR VPWR booth_b52_m40 sky130_fd_sc_hd__xor2_1
XU$$2915 net1168 net520 net1159 net793 VGND VGND VPWR VPWR t$5895 sky130_fd_sc_hd__a22o_1
XU$$2926 t$5900 net1371 VGND VGND VPWR VPWR booth_b42_m21 sky130_fd_sc_hd__xor2_1
XTAP_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_220 net1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2937 net1070 net522 net1062 net795 VGND VGND VPWR VPWR t$5906 sky130_fd_sc_hd__a22o_1
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2948 t$5911 net1368 VGND VGND VPWR VPWR booth_b42_m32 sky130_fd_sc_hd__xor2_1
XFILLER_61_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_231 net1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2959 net958 net522 net951 net795 VGND VGND VPWR VPWR t$5917 sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_22_1 pp_row22_5 pp_row22_6 pp_row22_7 VGND VGND VPWR VPWR c$2016 s$2017
+ sky130_fd_sc_hd__fa_1
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_242 net1522 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_253 net1619 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_264 net1723 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_16
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_275 c$1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_286 sel_1$4968 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_297 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0860_ clknet_leaf_102_clk booth_b30_m64 VGND VGND VPWR VPWR pp_row94_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_173_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0791_ clknet_leaf_194_clk net246 VGND VGND VPWR VPWR pp_row90_21 sky130_fd_sc_hd__dfxtp_2
XFILLER_158_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2461_ clknet_leaf_95_clk booth_b32_m36 VGND VGND VPWR VPWR pp_row68_15 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_81_5 s$915 s$917 s$919 VGND VGND VPWR VPWR c$1708 s$1709 sky130_fd_sc_hd__fa_1
X_1412_ clknet_leaf_41_clk booth_b32_m1 VGND VGND VPWR VPWR pp_row33_16 sky130_fd_sc_hd__dfxtp_1
X_2392_ clknet_leaf_179_clk notsign$6574 VGND VGND VPWR VPWR pp_row125_0 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_74_4 s$785 s$787 s$789 VGND VGND VPWR VPWR c$1622 s$1623 sky130_fd_sc_hd__fa_1
X_1343_ clknet_leaf_3_clk booth_b18_m12 VGND VGND VPWR VPWR pp_row30_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_110_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_67_3 c$652 s$655 s$657 VGND VGND VPWR VPWR c$1536 s$1537 sky130_fd_sc_hd__fa_1
X_1274_ clknet_leaf_11_clk booth_b22_m4 VGND VGND VPWR VPWR pp_row26_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_37_1 s$2913 s$2915 s$2917 VGND VGND VPWR VPWR c$3546 s$3547 sky130_fd_sc_hd__fa_1
X_0225_ clknet_leaf_208_clk booth_b24_m47 VGND VGND VPWR VPWR pp_row71_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_37_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_16_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_189_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_111_1 s$3357 s$3359 s$3361 VGND VGND VPWR VPWR c$3842 s$3843 sky130_fd_sc_hd__fa_1
XFILLER_146_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0989_ clknet_leaf_118_clk booth_b52_m48 VGND VGND VPWR VPWR pp_row100_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_104_0 c$3308 c$3310 c$3312 VGND VGND VPWR VPWR c$3812 s$3813 sky130_fd_sc_hd__fa_1
XFILLER_118_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_62_2 pp_row62_23 pp_row62_24 pp_row62_25 VGND VGND VPWR VPWR c$568 s$569
+ sky130_fd_sc_hd__fa_1
XFILLER_170_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_55_1 pp_row55_8 pp_row55_9 pp_row55_10 VGND VGND VPWR VPWR c$440 s$441
+ sky130_fd_sc_hd__fa_1
Xdadda_fa_4_32_0 s$1121 c$2086 c$2088 VGND VGND VPWR VPWR c$2882 s$2883 sky130_fd_sc_hd__fa_1
XFILLER_28_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_48_0 pp_row48_0 pp_row48_1 pp_row48_2 VGND VGND VPWR VPWR c$316 s$317
+ sky130_fd_sc_hd__fa_1
XFILLER_55_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_84_3 s$1739 s$1741 s$1743 VGND VGND VPWR VPWR c$2516 s$2517 sky130_fd_sc_hd__fa_1
XFILLER_163_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_77_2 c$1648 s$1651 s$1653 VGND VGND VPWR VPWR c$2458 s$2459 sky130_fd_sc_hd__fa_1
XFILLER_112_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_876 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1600 net1602 VGND VGND VPWR VPWR net1600 sky130_fd_sc_hd__buf_4
Xfanout1611 net116 VGND VGND VPWR VPWR net1611 sky130_fd_sc_hd__clkbuf_4
Xfanout1622 net1628 VGND VGND VPWR VPWR net1622 sky130_fd_sc_hd__clkbuf_8
Xfanout1633 net1637 VGND VGND VPWR VPWR net1633 sky130_fd_sc_hd__clkbuf_8
Xfanout1644 net1645 VGND VGND VPWR VPWR net1644 sky130_fd_sc_hd__buf_4
Xdadda_fa_6_47_0 c$3580 c$3582 s$3585 VGND VGND VPWR VPWR c$3990 s$3991 sky130_fd_sc_hd__fa_1
Xfanout1655 net1656 VGND VGND VPWR VPWR net1655 sky130_fd_sc_hd__clkbuf_8
XU$$4103 net1548 net453 net1540 net726 VGND VGND VPWR VPWR t$6501 sky130_fd_sc_hd__a22o_1
XFILLER_78_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4114 notblock$6505\[2\] net57 net1284 t$6506 notblock$6505\[0\] VGND VGND VPWR
+ VPWR sel_0$6507 sky130_fd_sc_hd__a32o_1
Xfanout1666 net1667 VGND VGND VPWR VPWR net1666 sky130_fd_sc_hd__buf_6
XU$$4125 t$6513 net1269 VGND VGND VPWR VPWR booth_b60_m4 sky130_fd_sc_hd__xor2_1
XFILLER_93_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1677 net1678 VGND VGND VPWR VPWR net1677 sky130_fd_sc_hd__buf_6
Xfanout1688 net1689 VGND VGND VPWR VPWR net1688 sky130_fd_sc_hd__buf_6
XU$$4136 net1498 net437 net1223 net719 VGND VGND VPWR VPWR t$6519 sky130_fd_sc_hd__a22o_1
Xfanout690 net691 VGND VGND VPWR VPWR net690 sky130_fd_sc_hd__buf_4
XU$$4147 t$6524 net1263 VGND VGND VPWR VPWR booth_b60_m15 sky130_fd_sc_hd__xor2_1
XU$$3402 net1636 net499 net1626 net772 VGND VGND VPWR VPWR t$6143 sky130_fd_sc_hd__a22o_1
Xfanout1699 net106 VGND VGND VPWR VPWR net1699 sky130_fd_sc_hd__clkbuf_2
XU$$3413 t$6148 net1340 VGND VGND VPWR VPWR booth_b48_m59 sky130_fd_sc_hd__xor2_1
XU$$4158 net1119 net436 net1112 net718 VGND VGND VPWR VPWR t$6530 sky130_fd_sc_hd__a22o_1
XU$$4169 t$6535 net1268 VGND VGND VPWR VPWR booth_b60_m26 sky130_fd_sc_hd__xor2_1
XU$$3424 net1345 VGND VGND VPWR VPWR notsign$6154 sky130_fd_sc_hd__inv_1
XU$$3435 net1129 net488 net1037 net761 VGND VGND VPWR VPWR t$6161 sky130_fd_sc_hd__a22o_1
XU$$2701 net1713 net545 net1704 net818 VGND VGND VPWR VPWR t$5785 sky130_fd_sc_hd__a22o_1
Xclkbuf_5_3__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_5_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XU$$3446 t$6166 net1337 VGND VGND VPWR VPWR booth_b50_m7 sky130_fd_sc_hd__xor2_1
XU$$3457 net1205 net484 net1196 net757 VGND VGND VPWR VPWR t$6172 sky130_fd_sc_hd__a22o_1
XU$$2712 t$5790 net1397 VGND VGND VPWR VPWR booth_b38_m51 sky130_fd_sc_hd__xor2_1
XTAP_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2723 net1611 net547 net1603 net820 VGND VGND VPWR VPWR t$5796 sky130_fd_sc_hd__a22o_1
XFILLER_92_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_106_2 s$2689 s$2691 s$2693 VGND VGND VPWR VPWR c$3330 s$3331 sky130_fd_sc_hd__fa_1
XU$$3468 t$6177 net1333 VGND VGND VPWR VPWR booth_b50_m18 sky130_fd_sc_hd__xor2_1
XTAP_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2734 t$5801 net1401 VGND VGND VPWR VPWR booth_b38_m62 sky130_fd_sc_hd__xor2_1
XU$$3479 net1090 net484 net1082 net757 VGND VGND VPWR VPWR t$6183 sky130_fd_sc_hd__a22o_1
XU$$4483_1862 VGND VGND VPWR VPWR U$$4483_1862/HI net1862 sky130_fd_sc_hd__conb_1
XTAP_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2745 net35 net1398 VGND VGND VPWR VPWR sel_1$5808 sky130_fd_sc_hd__xor2_1
XU$$2756 net1672 net536 net1562 net809 VGND VGND VPWR VPWR t$5814 sky130_fd_sc_hd__a22o_1
XTAP_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2767 t$5819 net1381 VGND VGND VPWR VPWR booth_b40_m10 sky130_fd_sc_hd__xor2_1
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2778 net1172 net539 net1163 net812 VGND VGND VPWR VPWR t$5825 sky130_fd_sc_hd__a22o_1
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2789 t$5830 net1377 VGND VGND VPWR VPWR booth_b40_m21 sky130_fd_sc_hd__xor2_1
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1961_ clknet_leaf_138_clk booth_b48_m60 VGND VGND VPWR VPWR pp_row108_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1090 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0912_ clknet_leaf_104_clk booth_b50_m46 VGND VGND VPWR VPWR pp_row96_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_159_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1892_ clknet_leaf_64_clk booth_b16_m36 VGND VGND VPWR VPWR pp_row52_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0843_ clknet_leaf_106_clk booth_b38_m55 VGND VGND VPWR VPWR pp_row93_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0774_ clknet_leaf_141_clk booth_b36_m54 VGND VGND VPWR VPWR pp_row90_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_6_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2444_ clknet_leaf_198_clk net220 VGND VGND VPWR VPWR pp_row67_33 sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_5_clk clknet_5_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_64_1020 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_72_1 c$730 c$732 c$734 VGND VGND VPWR VPWR c$1592 s$1593 sky130_fd_sc_hd__fa_1
XFILLER_69_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2375_ clknet_leaf_85_clk booth_b10_m56 VGND VGND VPWR VPWR pp_row66_5 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_65_0 s$107 c$600 c$602 VGND VGND VPWR VPWR c$1506 s$1507 sky130_fd_sc_hd__fa_2
XFILLER_151_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$707 final_adder.p_new$714 final_adder.g_new$731 final_adder.g_new$715
+ VGND VGND VPWR VPWR final_adder.g_new$835 sky130_fd_sc_hd__a21o_1
X_1326_ clknet_leaf_1_clk booth_b20_m9 VGND VGND VPWR VPWR pp_row29_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$718 final_adder.p_new$742 final_adder.p_new$726 VGND VGND VPWR VPWR
+ final_adder.p_new$846 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$729 final_adder.p_new$736 final_adder.g_new$753 final_adder.g_new$737
+ VGND VGND VPWR VPWR final_adder.g_new$857 sky130_fd_sc_hd__a21o_2
XFILLER_57_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1257_ clknet_leaf_11_clk booth_b20_m5 VGND VGND VPWR VPWR pp_row25_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_37_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0208_ clknet_leaf_151_clk booth_b56_m14 VGND VGND VPWR VPWR pp_row70_26 sky130_fd_sc_hd__dfxtp_1
XFILLER_37_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1188_ clknet_leaf_49_clk booth_b2_m19 VGND VGND VPWR VPWR pp_row21_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_52_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3980 t$6439 net1287 VGND VGND VPWR VPWR booth_b58_m0 sky130_fd_sc_hd__xor2_1
XU$$3991 net1566 net458 net1525 net731 VGND VGND VPWR VPWR t$6445 sky130_fd_sc_hd__a22o_1
XFILLER_52_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1915_1768 VGND VGND VPWR VPWR U$$1915_1768/HI net1768 sky130_fd_sc_hd__conb_1
XFILLER_193_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_94_2 s$2593 s$2595 s$2597 VGND VGND VPWR VPWR c$3258 s$3259 sky130_fd_sc_hd__fa_1
XFILLER_192_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_939 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_87_1 c$2530 c$2532 s$2535 VGND VGND VPWR VPWR c$3214 s$3215 sky130_fd_sc_hd__fa_1
XFILLER_106_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_64_0 s$3655 c$4022 s$4025 VGND VGND VPWR VPWR c$4280 s$4281 sky130_fd_sc_hd__fa_1
XFILLER_134_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput260 net260 VGND VGND VPWR VPWR o[102] sky130_fd_sc_hd__buf_2
XFILLER_161_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput271 net271 VGND VGND VPWR VPWR o[112] sky130_fd_sc_hd__buf_2
XFILLER_0_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput282 net282 VGND VGND VPWR VPWR o[122] sky130_fd_sc_hd__buf_2
Xoutput293 net293 VGND VGND VPWR VPWR o[17] sky130_fd_sc_hd__buf_2
XFILLER_0_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2008 net1751 net591 net1743 net864 VGND VGND VPWR VPWR t$5431 sky130_fd_sc_hd__a22o_1
XU$$2019 t$5436 net1454 VGND VGND VPWR VPWR booth_b28_m47 sky130_fd_sc_hd__xor2_1
XU$$1307 net992 net637 net987 net910 VGND VGND VPWR VPWR t$5073 sky130_fd_sc_hd__a22o_1
XFILLER_15_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1318 t$5078 net1666 VGND VGND VPWR VPWR booth_b18_m39 sky130_fd_sc_hd__xor2_1
XFILLER_167_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1329 net1721 net640 net1712 net913 VGND VGND VPWR VPWR t$5084 sky130_fd_sc_hd__a22o_1
XFILLER_167_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$280_1783 VGND VGND VPWR VPWR U$$280_1783/HI net1783 sky130_fd_sc_hd__conb_1
XFILLER_11_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_82_0 s$937 c$1698 c$1700 VGND VGND VPWR VPWR c$2494 s$2495 sky130_fd_sc_hd__fa_1
XFILLER_124_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0490_ clknet_leaf_159_clk booth_b46_m33 VGND VGND VPWR VPWR pp_row79_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_140_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_964 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1430 net1431 VGND VGND VPWR VPWR net1430 sky130_fd_sc_hd__buf_6
Xfanout1441 net1442 VGND VGND VPWR VPWR net1441 sky130_fd_sc_hd__buf_6
Xfanout1452 net1456 VGND VGND VPWR VPWR net1452 sky130_fd_sc_hd__buf_8
X_2160_ clknet_leaf_136_clk booth_b60_m49 VGND VGND VPWR VPWR pp_row109_8 sky130_fd_sc_hd__dfxtp_1
Xfanout1463 net1465 VGND VGND VPWR VPWR net1463 sky130_fd_sc_hd__clkbuf_8
XFILLER_120_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1474 net18 VGND VGND VPWR VPWR net1474 sky130_fd_sc_hd__buf_8
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1485 net1486 VGND VGND VPWR VPWR net1485 sky130_fd_sc_hd__buf_6
XFILLER_4_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1111_ clknet_leaf_15_clk net1185 VGND VGND VPWR VPWR pp_row14_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_120_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1496 net1498 VGND VGND VPWR VPWR net1496 sky130_fd_sc_hd__buf_4
XFILLER_24_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3210 t$6045 net1348 VGND VGND VPWR VPWR booth_b46_m26 sky130_fd_sc_hd__xor2_1
XFILLER_66_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2091_ clknet_leaf_37_clk booth_b20_m38 VGND VGND VPWR VPWR pp_row58_10 sky130_fd_sc_hd__dfxtp_1
XU$$3221 net1019 net503 net1002 net776 VGND VGND VPWR VPWR t$6051 sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_44_5 s$269 s$271 s$273 VGND VGND VPWR VPWR c$1264 s$1265 sky130_fd_sc_hd__fa_1
Xdadda_fa_4_111_0 pp_row111_9 pp_row111_10 c$2718 VGND VGND VPWR VPWR c$3356 s$3357
+ sky130_fd_sc_hd__fa_1
XU$$3232 t$6056 net1351 VGND VGND VPWR VPWR booth_b46_m37 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$14 c$4178 s$4181 VGND VGND VPWR VPWR final_adder.$signal$30 final_adder.$signal$1104
+ sky130_fd_sc_hd__ha_1
X_1042_ clknet_leaf_64_clk booth_b4_m2 VGND VGND VPWR VPWR pp_row6_2 sky130_fd_sc_hd__dfxtp_1
XU$$3243 net1740 net504 net1732 net777 VGND VGND VPWR VPWR t$6062 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$25 c$4200 s$4203 VGND VGND VPWR VPWR final_adder.$signal$52 final_adder.$signal$1115
+ sky130_fd_sc_hd__ha_1
XU$$3254 t$6067 net1355 VGND VGND VPWR VPWR booth_b46_m48 sky130_fd_sc_hd__xor2_1
XFILLER_0_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3265 net1635 net508 net1626 net781 VGND VGND VPWR VPWR t$6073 sky130_fd_sc_hd__a22o_1
XU$$2520 net1090 net553 net1082 net826 VGND VGND VPWR VPWR t$5693 sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_37_4 pp_row37_17 pp_row37_18 pp_row37_19 VGND VGND VPWR VPWR c$1178 s$1179
+ sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$36 c$4222 s$4225 VGND VGND VPWR VPWR final_adder.$signal$74 final_adder.$signal$1126
+ sky130_fd_sc_hd__ha_1
XU$$2531 t$5698 net1407 VGND VGND VPWR VPWR booth_b36_m29 sky130_fd_sc_hd__xor2_1
XU$$3276 t$6078 net1356 VGND VGND VPWR VPWR booth_b46_m59 sky130_fd_sc_hd__xor2_1
XFILLER_94_1024 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$47 c$4244 s$4247 VGND VGND VPWR VPWR final_adder.$signal$96 final_adder.$signal$1137
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$58 c$4266 s$4269 VGND VGND VPWR VPWR final_adder.$signal$118 final_adder.$signal$1148
+ sky130_fd_sc_hd__ha_1
XFILLER_34_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2542 net984 net555 net975 net828 VGND VGND VPWR VPWR t$5704 sky130_fd_sc_hd__a22o_1
XU$$3287 net1356 VGND VGND VPWR VPWR notsign$6084 sky130_fd_sc_hd__inv_1
Xfinal_adder.U$$69 c$4288 s$4291 VGND VGND VPWR VPWR final_adder.$signal$140 final_adder.$signal$1159
+ sky130_fd_sc_hd__ha_1
XU$$2553 t$5709 net1409 VGND VGND VPWR VPWR booth_b36_m40 sky130_fd_sc_hd__xor2_1
XU$$3298 net1125 net493 net1034 net766 VGND VGND VPWR VPWR t$6091 sky130_fd_sc_hd__a22o_1
XFILLER_181_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2564 net1713 net556 net1704 net829 VGND VGND VPWR VPWR t$5715 sky130_fd_sc_hd__a22o_1
XU$$2575 t$5720 net1408 VGND VGND VPWR VPWR booth_b36_m51 sky130_fd_sc_hd__xor2_1
XU$$1830 t$5340 net1459 VGND VGND VPWR VPWR booth_b26_m21 sky130_fd_sc_hd__xor2_1
XU$$2586 net1611 net557 net1599 net830 VGND VGND VPWR VPWR t$5726 sky130_fd_sc_hd__a22o_1
XU$$1841 net1066 net596 net1057 net869 VGND VGND VPWR VPWR t$5346 sky130_fd_sc_hd__a22o_1
XFILLER_22_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2597 t$5731 net1411 VGND VGND VPWR VPWR booth_b36_m62 sky130_fd_sc_hd__xor2_1
XFILLER_181_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1852 t$5351 net1462 VGND VGND VPWR VPWR booth_b26_m32 sky130_fd_sc_hd__xor2_1
XU$$1863 net961 net597 net955 net870 VGND VGND VPWR VPWR t$5357 sky130_fd_sc_hd__a22o_1
XU$$1874 t$5362 net1465 VGND VGND VPWR VPWR booth_b26_m43 sky130_fd_sc_hd__xor2_1
XU$$1885 net1687 net598 net1679 net871 VGND VGND VPWR VPWR t$5368 sky130_fd_sc_hd__a22o_1
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1896 t$5373 net1463 VGND VGND VPWR VPWR booth_b26_m54 sky130_fd_sc_hd__xor2_1
X_1944_ clknet_leaf_78_clk booth_b52_m1 VGND VGND VPWR VPWR pp_row53_26 sky130_fd_sc_hd__dfxtp_1
XFILLER_148_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1875_ clknet_leaf_69_clk booth_b38_m13 VGND VGND VPWR VPWR pp_row51_19 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_97_0 c$3266 c$3268 c$3270 VGND VGND VPWR VPWR c$3784 s$3785 sky130_fd_sc_hd__fa_1
XFILLER_163_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0826_ clknet_leaf_108_clk booth_b48_m44 VGND VGND VPWR VPWR pp_row92_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0757_ clknet_leaf_160_clk booth_b46_m43 VGND VGND VPWR VPWR pp_row89_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_127_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0688_ clknet_leaf_131_clk booth_b64_m53 VGND VGND VPWR VPWR pp_row117_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_131_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2427_ clknet_leaf_98_clk booth_b34_m33 VGND VGND VPWR VPWR pp_row67_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_130_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2358_ clknet_leaf_77_clk booth_b46_m19 VGND VGND VPWR VPWR pp_row65_23 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$515 final_adder.p_new$518 final_adder.g_new$527 final_adder.g_new$519
+ VGND VGND VPWR VPWR final_adder.g_new$643 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$526 final_adder.p_new$538 final_adder.p_new$530 VGND VGND VPWR VPWR
+ final_adder.p_new$654 sky130_fd_sc_hd__and2_1
XTAP_3808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$537 final_adder.p_new$540 final_adder.g_new$549 final_adder.g_new$541
+ VGND VGND VPWR VPWR final_adder.g_new$665 sky130_fd_sc_hd__a21o_1
XFILLER_28_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1309_ clknet_leaf_3_clk booth_b22_m6 VGND VGND VPWR VPWR pp_row28_11 sky130_fd_sc_hd__dfxtp_1
XU$$4386_1811 VGND VGND VPWR VPWR U$$4386_1811/HI net1811 sky130_fd_sc_hd__conb_1
Xfinal_adder.U$$548 final_adder.p_new$560 final_adder.p_new$552 VGND VGND VPWR VPWR
+ final_adder.p_new$676 sky130_fd_sc_hd__and2_1
XFILLER_84_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2289_ clknet_leaf_214_clk booth_b52_m11 VGND VGND VPWR VPWR pp_row63_26 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$559 final_adder.p_new$562 final_adder.g_new$571 final_adder.g_new$563
+ VGND VGND VPWR VPWR final_adder.g_new$687 sky130_fd_sc_hd__a21o_1
XU$$409 t$4613 net1280 VGND VGND VPWR VPWR booth_b4_m64 sky130_fd_sc_hd__xor2_1
XFILLER_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_106_1 pp_row106_8 pp_row106_9 pp_row106_10 VGND VGND VPWR VPWR c$2688
+ s$2689 sky130_fd_sc_hd__fa_1
XFILLER_122_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_127_0 pp_row127_0 pp_row127_1 pp_row127_2 VGND VGND VPWR VPWR dadda_fa_6_127_0/COUT
+ s$4151 sky130_fd_sc_hd__fa_1
XFILLER_76_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3011_1786 VGND VGND VPWR VPWR U$$3011_1786/HI net1786 sky130_fd_sc_hd__conb_1
XFILLER_48_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_47_3 s$1295 s$1297 s$1299 VGND VGND VPWR VPWR c$2220 s$2221 sky130_fd_sc_hd__fa_1
XFILLER_47_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$910 net931 net397 net1752 net663 VGND VGND VPWR VPWR t$4870 sky130_fd_sc_hd__a22o_1
XFILLER_16_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$921 t$4875 net1314 VGND VGND VPWR VPWR booth_b12_m46 sky130_fd_sc_hd__xor2_1
XFILLER_169_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$932 net1649 net399 net1641 net665 VGND VGND VPWR VPWR t$4881 sky130_fd_sc_hd__a22o_1
XFILLER_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$943 t$4886 net1318 VGND VGND VPWR VPWR booth_b12_m57 sky130_fd_sc_hd__xor2_1
XU$$954 net1535 net395 net1527 net661 VGND VGND VPWR VPWR t$4892 sky130_fd_sc_hd__a22o_1
XFILLER_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1104 net1228 net644 net1123 net917 VGND VGND VPWR VPWR t$4970 sky130_fd_sc_hd__a22o_1
XU$$965 net1889 net387 net1228 net653 VGND VGND VPWR VPWR t$4899 sky130_fd_sc_hd__a22o_1
XU$$976 t$4904 net1187 VGND VGND VPWR VPWR booth_b14_m5 sky130_fd_sc_hd__xor2_1
XU$$1115 t$4975 net1009 VGND VGND VPWR VPWR booth_b16_m6 sky130_fd_sc_hd__xor2_1
XFILLER_141_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1126 net1210 net643 net1201 net916 VGND VGND VPWR VPWR t$4981 sky130_fd_sc_hd__a22o_1
XU$$987 net1220 net385 net1210 net651 VGND VGND VPWR VPWR t$4910 sky130_fd_sc_hd__a22o_1
XU$$1137 t$4986 net1009 VGND VGND VPWR VPWR booth_b16_m17 sky130_fd_sc_hd__xor2_1
XU$$998 t$4915 net1183 VGND VGND VPWR VPWR booth_b14_m16 sky130_fd_sc_hd__xor2_1
XU$$1148 net1099 net643 net1089 net916 VGND VGND VPWR VPWR t$4992 sky130_fd_sc_hd__a22o_1
XU$$1159 t$4997 net1007 VGND VGND VPWR VPWR booth_b16_m28 sky130_fd_sc_hd__xor2_1
XFILLER_70_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1022 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1660_ clknet_leaf_21_clk booth_b14_m30 VGND VGND VPWR VPWR pp_row44_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0611_ clknet_leaf_179_clk booth_b64_m62 VGND VGND VPWR VPWR pp_row126_2 sky130_fd_sc_hd__dfxtp_1
X_1591_ clknet_leaf_5_clk booth_b28_m13 VGND VGND VPWR VPWR pp_row41_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_125_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0542_ clknet_leaf_170_clk booth_b36_m45 VGND VGND VPWR VPWR pp_row81_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_140_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_791 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0473_ clknet_leaf_193_clk booth_b16_m63 VGND VGND VPWR VPWR pp_row79_1 sky130_fd_sc_hd__dfxtp_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2212_ clknet_leaf_217_clk booth_b46_m15 VGND VGND VPWR VPWR pp_row61_23 sky130_fd_sc_hd__dfxtp_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1260 net1261 VGND VGND VPWR VPWR net1260 sky130_fd_sc_hd__buf_6
XFILLER_66_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1271 net1272 VGND VGND VPWR VPWR net1271 sky130_fd_sc_hd__buf_6
XFILLER_38_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2143_ clknet_leaf_219_clk booth_b50_m9 VGND VGND VPWR VPWR pp_row59_25 sky130_fd_sc_hd__dfxtp_1
Xfanout1282 net55 VGND VGND VPWR VPWR net1282 sky130_fd_sc_hd__buf_6
XFILLER_61_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1293 net1294 VGND VGND VPWR VPWR net1293 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_42_2 pp_row42_20 pp_row42_21 pp_row42_22 VGND VGND VPWR VPWR c$1234 s$1235
+ sky130_fd_sc_hd__fa_1
XFILLER_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3040 net1501 net514 net1226 net787 VGND VGND VPWR VPWR t$5959 sky130_fd_sc_hd__a22o_1
XFILLER_66_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2074_ clknet_leaf_32_clk booth_b48_m9 VGND VGND VPWR VPWR pp_row57_24 sky130_fd_sc_hd__dfxtp_1
XU$$3051 t$5964 net1358 VGND VGND VPWR VPWR booth_b44_m15 sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_35_1 pp_row35_5 pp_row35_6 pp_row35_7 VGND VGND VPWR VPWR c$1148 s$1149
+ sky130_fd_sc_hd__fa_1
XU$$3062 net1121 net514 net1113 net787 VGND VGND VPWR VPWR t$5970 sky130_fd_sc_hd__a22o_1
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1025_ clknet_leaf_249_clk net179 VGND VGND VPWR VPWR pp_row2_3 sky130_fd_sc_hd__dfxtp_4
XU$$3073 t$5975 net1360 VGND VGND VPWR VPWR booth_b44_m26 sky130_fd_sc_hd__xor2_1
XU$$3084 net1019 net512 net1002 net785 VGND VGND VPWR VPWR t$5981 sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_12_0 pp_row12_8 c$2758 c$2760 VGND VGND VPWR VPWR c$3444 s$3445 sky130_fd_sc_hd__fa_1
XU$$2350 t$5606 net1420 VGND VGND VPWR VPWR booth_b34_m7 sky130_fd_sc_hd__xor2_1
XU$$3095 t$5986 net1359 VGND VGND VPWR VPWR booth_b44_m37 sky130_fd_sc_hd__xor2_1
XU$$2361 net1202 net560 net1193 net833 VGND VGND VPWR VPWR t$5612 sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_28_0 pp_row28_0 pp_row28_1 pp_row28_2 VGND VGND VPWR VPWR c$1074 s$1075
+ sky130_fd_sc_hd__fa_1
XU$$2372 t$5617 net1423 VGND VGND VPWR VPWR booth_b34_m18 sky130_fd_sc_hd__xor2_1
XFILLER_35_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2383 net1092 net563 net1084 net836 VGND VGND VPWR VPWR t$5623 sky130_fd_sc_hd__a22o_1
XFILLER_22_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2394 t$5628 net1422 VGND VGND VPWR VPWR booth_b34_m29 sky130_fd_sc_hd__xor2_1
XU$$1660 net1671 net602 net1560 net875 VGND VGND VPWR VPWR t$5254 sky130_fd_sc_hd__a22o_1
XU$$1671 t$5259 net1469 VGND VGND VPWR VPWR booth_b24_m10 sky130_fd_sc_hd__xor2_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1682 net1164 net603 net1155 net876 VGND VGND VPWR VPWR t$5265 sky130_fd_sc_hd__a22o_1
XFILLER_148_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1693 t$5270 net1467 VGND VGND VPWR VPWR booth_b24_m21 sky130_fd_sc_hd__xor2_1
XFILLER_30_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1927_ clknet_leaf_184_clk net137 VGND VGND VPWR VPWR pp_row107_12 sky130_fd_sc_hd__dfxtp_2
XFILLER_163_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1858_ clknet_leaf_78_clk booth_b8_m43 VGND VGND VPWR VPWR pp_row51_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0809_ clknet_leaf_97_clk booth_b58_m33 VGND VGND VPWR VPWR pp_row91_16 sky130_fd_sc_hd__dfxtp_1
X_1789_ clknet_leaf_221_clk booth_b46_m2 VGND VGND VPWR VPWR pp_row48_23 sky130_fd_sc_hd__dfxtp_1
XFILLER_157_1040 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_87_4 pp_row87_12 pp_row87_13 pp_row87_14 VGND VGND VPWR VPWR c$998 s$999
+ sky130_fd_sc_hd__fa_1
XFILLER_118_1013 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_57_2 s$2297 s$2299 s$2301 VGND VGND VPWR VPWR c$3036 s$3037 sky130_fd_sc_hd__fa_1
XTAP_4306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$301 final_adder.p_new$300 final_adder.g_new$303 final_adder.g_new$301
+ VGND VGND VPWR VPWR final_adder.g_new$429 sky130_fd_sc_hd__a21o_1
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$312 final_adder.p_new$314 final_adder.p_new$312 VGND VGND VPWR VPWR
+ final_adder.p_new$440 sky130_fd_sc_hd__and2_1
XTAP_4328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$323 final_adder.p_new$322 final_adder.g_new$325 final_adder.g_new$323
+ VGND VGND VPWR VPWR final_adder.g_new$451 sky130_fd_sc_hd__a21o_1
XFILLER_29_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$334 final_adder.p_new$336 final_adder.p_new$334 VGND VGND VPWR VPWR
+ final_adder.p_new$462 sky130_fd_sc_hd__and2_1
XTAP_3616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$345 final_adder.p_new$344 final_adder.g_new$347 final_adder.g_new$345
+ VGND VGND VPWR VPWR final_adder.g_new$473 sky130_fd_sc_hd__a21o_1
XTAP_3627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_27_0 s$3507 c$3948 s$3951 VGND VGND VPWR VPWR c$4206 s$4207 sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$356 final_adder.p_new$358 final_adder.p_new$356 VGND VGND VPWR VPWR
+ final_adder.p_new$484 sky130_fd_sc_hd__and2_1
XTAP_3638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_220_clk clknet_5_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_220_clk
+ sky130_fd_sc_hd__clkbuf_16
XU$$206 t$4510 net1389 VGND VGND VPWR VPWR booth_b2_m31 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$367 final_adder.p_new$366 final_adder.g_new$369 final_adder.g_new$367
+ VGND VGND VPWR VPWR final_adder.g_new$495 sky130_fd_sc_hd__a21o_1
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$378 final_adder.p_new$380 final_adder.p_new$378 VGND VGND VPWR VPWR
+ final_adder.p_new$506 sky130_fd_sc_hd__and2_1
XU$$217 net968 net625 net957 net898 VGND VGND VPWR VPWR t$4516 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$389 final_adder.p_new$390 final_adder.g_new$395 final_adder.g_new$391
+ VGND VGND VPWR VPWR final_adder.g_new$517 sky130_fd_sc_hd__a21o_1
XU$$228 t$4521 net1388 VGND VGND VPWR VPWR booth_b2_m42 sky130_fd_sc_hd__xor2_1
XFILLER_72_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$239 net1695 net621 net1687 net894 VGND VGND VPWR VPWR t$4527 sky130_fd_sc_hd__a22o_1
XFILLER_44_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2609_1779 VGND VGND VPWR VPWR U$$2609_1779/HI net1779 sky130_fd_sc_hd__conb_1
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_1050 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1023 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_52_1 c$1342 c$1344 c$1346 VGND VGND VPWR VPWR c$2256 s$2257 sky130_fd_sc_hd__fa_1
XFILLER_0_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_0_68_1 pp_row68_3 pp_row68_4 pp_row68_5 VGND VGND VPWR VPWR c$134 s$135
+ sky130_fd_sc_hd__fa_1
XFILLER_48_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_45_0 s$287 c$1254 c$1256 VGND VGND VPWR VPWR c$2198 s$2199 sky130_fd_sc_hd__fa_1
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_211_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_211_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_152_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$740 t$4783 net1414 VGND VGND VPWR VPWR booth_b10_m24 sky130_fd_sc_hd__xor2_1
XU$$751 net1040 net402 net1024 net668 VGND VGND VPWR VPWR t$4789 sky130_fd_sc_hd__a22o_1
XFILLER_17_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$762 t$4794 net1416 VGND VGND VPWR VPWR booth_b10_m35 sky130_fd_sc_hd__xor2_1
XU$$773 net931 net407 net1749 net673 VGND VGND VPWR VPWR t$4800 sky130_fd_sc_hd__a22o_1
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$784 t$4805 net1419 VGND VGND VPWR VPWR booth_b10_m46 sky130_fd_sc_hd__xor2_1
XFILLER_188_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$795 net1646 net403 net1638 net669 VGND VGND VPWR VPWR t$4811 sky130_fd_sc_hd__a22o_1
XFILLER_17_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_2_98_5 pp_row98_15 pp_row98_16 VGND VGND VPWR VPWR c$1912 s$1913 sky130_fd_sc_hd__ha_1
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1712_ clknet_leaf_236_clk booth_b10_m36 VGND VGND VPWR VPWR pp_row46_5 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_7_102_0 s$3807 c$4098 s$4101 VGND VGND VPWR VPWR c$4356 s$4357 sky130_fd_sc_hd__fa_1
XFILLER_129_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1 c$1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1643_ clknet_leaf_6_clk booth_b28_m15 VGND VGND VPWR VPWR pp_row43_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_133_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_97_3 pp_row97_9 pp_row97_10 pp_row97_11 VGND VGND VPWR VPWR c$1896 s$1897
+ sky130_fd_sc_hd__fa_1
XFILLER_99_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1574_ clknet_leaf_21_clk net1376 VGND VGND VPWR VPWR pp_row40_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_141_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_67_1 s$3093 s$3095 s$3097 VGND VGND VPWR VPWR c$3666 s$3667 sky130_fd_sc_hd__fa_1
X_0525_ clknet_leaf_162_clk booth_b56_m24 VGND VGND VPWR VPWR pp_row80_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_112_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout508 net509 VGND VGND VPWR VPWR net508 sky130_fd_sc_hd__buf_4
Xfanout519 net520 VGND VGND VPWR VPWR net519 sky130_fd_sc_hd__buf_4
XFILLER_63_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0456_ clknet_leaf_158_clk booth_b38_m40 VGND VGND VPWR VPWR pp_row78_13 sky130_fd_sc_hd__dfxtp_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0387_ clknet_leaf_196_clk booth_b26_m50 VGND VGND VPWR VPWR pp_row76_8 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_59_8 s$33 s$35 s$37 VGND VGND VPWR VPWR c$526 s$527 sky130_fd_sc_hd__fa_2
Xclkbuf_leaf_202_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_202_clk
+ sky130_fd_sc_hd__clkbuf_16
Xfanout1090 net1093 VGND VGND VPWR VPWR net1090 sky130_fd_sc_hd__buf_6
XFILLER_82_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2126_ clknet_leaf_217_clk booth_b20_m39 VGND VGND VPWR VPWR pp_row59_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_67_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2057_ clknet_leaf_36_clk booth_b20_m37 VGND VGND VPWR VPWR pp_row57_10 sky130_fd_sc_hd__dfxtp_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_106_0 net1907 pp_row106_1 pp_row106_2 VGND VGND VPWR VPWR c$1966 s$1967
+ sky130_fd_sc_hd__fa_1
X_1008_ clknet_leaf_117_clk booth_b56_m45 VGND VGND VPWR VPWR pp_row101_10 sky130_fd_sc_hd__dfxtp_1
XU$$2180 t$5518 net1445 VGND VGND VPWR VPWR booth_b30_m59 sky130_fd_sc_hd__xor2_1
XU$$2191 net1447 VGND VGND VPWR VPWR notsign$5524 sky130_fd_sc_hd__inv_1
XFILLER_23_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1490 net1606 net632 net1596 net905 VGND VGND VPWR VPWR t$5166 sky130_fd_sc_hd__a22o_1
XFILLER_109_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_85_1 pp_row85_3 pp_row85_4 pp_row85_5 VGND VGND VPWR VPWR c$968 s$969
+ sky130_fd_sc_hd__fa_1
XFILLER_132_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_62_0 s$1481 c$2326 c$2328 VGND VGND VPWR VPWR c$3062 s$3063 sky130_fd_sc_hd__fa_1
Xdadda_fa_1_78_0 pp_row78_2 pp_row78_3 pp_row78_4 VGND VGND VPWR VPWR c$852 s$853
+ sky130_fd_sc_hd__fa_1
XFILLER_103_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$120 c$4390 s$4393 VGND VGND VPWR VPWR final_adder.$signal$242 final_adder.$signal$1210
+ sky130_fd_sc_hd__ha_2
Xfinal_adder.U$$131 final_adder.$signal$1215 final_adder.$signal$250 final_adder.$signal$252
+ VGND VGND VPWR VPWR final_adder.g_new$259 sky130_fd_sc_hd__a21o_1
XTAP_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3809 net1651 net473 net1643 net746 VGND VGND VPWR VPWR t$6351 sky130_fd_sc_hd__a22o_1
XTAP_4158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$142 final_adder.$signal$1202 final_adder.$signal$1203 VGND VGND VPWR
+ VPWR final_adder.p_new$270 sky130_fd_sc_hd__and2_1
XTAP_4169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$153 final_adder.$signal$1193 final_adder.$signal$206 final_adder.$signal$208
+ VGND VGND VPWR VPWR final_adder.g_new$281 sky130_fd_sc_hd__a21o_1
XTAP_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$164 final_adder.$signal$1180 final_adder.$signal$1181 VGND VGND VPWR
+ VPWR final_adder.p_new$292 sky130_fd_sc_hd__and2_1
XFILLER_174_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$175 final_adder.$signal$1171 final_adder.$signal$162 final_adder.$signal$164
+ VGND VGND VPWR VPWR final_adder.g_new$303 sky130_fd_sc_hd__a21o_1
XTAP_3457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$186 final_adder.$signal$1158 final_adder.$signal$1159 VGND VGND VPWR
+ VPWR final_adder.p_new$314 sky130_fd_sc_hd__and2_1
XANTENNA_402 net1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$197 final_adder.$signal$1149 final_adder.$signal$118 final_adder.$signal$120
+ VGND VGND VPWR VPWR final_adder.g_new$325 sky130_fd_sc_hd__a21o_1
XANTENNA_413 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_424 net592 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_435 net760 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_446 net1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_457 net1619 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_77_0 c$3700 c$3702 s$3705 VGND VGND VPWR VPWR c$4050 s$4051 sky130_fd_sc_hd__fa_1
XFILLER_123_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0310_ clknet_leaf_202_clk booth_b58_m15 VGND VGND VPWR VPWR pp_row73_25 sky130_fd_sc_hd__dfxtp_1
X_1290_ clknet_leaf_2_clk booth_b18_m9 VGND VGND VPWR VPWR pp_row27_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0241_ clknet_leaf_153_clk booth_b54_m17 VGND VGND VPWR VPWR pp_row71_24 sky130_fd_sc_hd__dfxtp_1
XFILLER_48_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput160 c[12] VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput171 c[22] VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_1
XFILLER_110_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput182 c[32] VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_1
Xinput193 c[42] VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__clkbuf_1
XFILLER_110_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0172_ clknet_leaf_101_clk booth_b52_m17 VGND VGND VPWR VPWR pp_row69_24 sky130_fd_sc_hd__dfxtp_1
XFILLER_64_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4447_1844 VGND VGND VPWR VPWR U$$4447_1844/HI net1844 sky130_fd_sc_hd__conb_1
XTAP_3980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$570 net1513 net410 net1505 net676 VGND VGND VPWR VPWR t$4697 sky130_fd_sc_hd__a22o_1
XFILLER_189_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$581 t$4702 net1240 VGND VGND VPWR VPWR booth_b8_m13 sky130_fd_sc_hd__xor2_1
XU$$592 net1138 net409 net1130 net675 VGND VGND VPWR VPWR t$4708 sky130_fd_sc_hd__a22o_1
XFILLER_108_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_104_0_1906 VGND VGND VPWR VPWR net1906 dadda_fa_2_104_0_1906/LO sky130_fd_sc_hd__conb_1
XFILLER_173_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_95_0 pp_row95_3 pp_row95_4 pp_row95_5 VGND VGND VPWR VPWR c$1866 s$1867
+ sky130_fd_sc_hd__fa_1
XFILLER_145_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1626_ clknet_leaf_236_clk net193 VGND VGND VPWR VPWR pp_row42_23 sky130_fd_sc_hd__dfxtp_1
XFILLER_126_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1557_ clknet_leaf_9_clk booth_b12_m28 VGND VGND VPWR VPWR pp_row40_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_87_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_71_7 c$158 c$160 c$162 VGND VGND VPWR VPWR c$740 s$741 sky130_fd_sc_hd__fa_1
XFILLER_115_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0508_ clknet_leaf_173_clk booth_b26_m54 VGND VGND VPWR VPWR pp_row80_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_59_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1488_ clknet_leaf_43_clk booth_b14_m23 VGND VGND VPWR VPWR pp_row37_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_115_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_64_6 c$76 c$78 c$80 VGND VGND VPWR VPWR c$612 s$613 sky130_fd_sc_hd__fa_1
XFILLER_74_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0439_ clknet_leaf_154_clk booth_b62_m15 VGND VGND VPWR VPWR pp_row77_25 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_57_5 pp_row57_23 pp_row57_24 pp_row57_25 VGND VGND VPWR VPWR c$484 s$485
+ sky130_fd_sc_hd__fa_1
XFILLER_67_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2109_ clknet_leaf_85_clk booth_b52_m6 VGND VGND VPWR VPWR pp_row58_26 sky130_fd_sc_hd__dfxtp_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_94_0 s$3775 c$4082 s$4085 VGND VGND VPWR VPWR c$4340 s$4341 sky130_fd_sc_hd__fa_1
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_975 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout850 net856 VGND VGND VPWR VPWR net850 sky130_fd_sc_hd__clkbuf_4
Xfanout861 net865 VGND VGND VPWR VPWR net861 sky130_fd_sc_hd__buf_6
XU$$4307 net1070 net418 net1062 net700 VGND VGND VPWR VPWR t$6606 sky130_fd_sc_hd__a22o_1
Xfanout872 net873 VGND VGND VPWR VPWR net872 sky130_fd_sc_hd__clkbuf_4
XU$$4318 t$6611 net1259 VGND VGND VPWR VPWR booth_b62_m32 sky130_fd_sc_hd__xor2_1
XU$$4329 net963 net424 net953 net706 VGND VGND VPWR VPWR t$6617 sky130_fd_sc_hd__a22o_1
Xfanout883 net885 VGND VGND VPWR VPWR net883 sky130_fd_sc_hd__buf_4
Xfanout894 net895 VGND VGND VPWR VPWR net894 sky130_fd_sc_hd__buf_4
XFILLER_46_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3606 net1142 net476 net1136 net749 VGND VGND VPWR VPWR t$6248 sky130_fd_sc_hd__a22o_1
XFILLER_92_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3617 t$6253 net1319 VGND VGND VPWR VPWR booth_b52_m24 sky130_fd_sc_hd__xor2_1
XTAP_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3628 net1043 net477 net1027 net750 VGND VGND VPWR VPWR t$6259 sky130_fd_sc_hd__a22o_1
XFILLER_133_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3639 t$6264 net1321 VGND VGND VPWR VPWR booth_b52_m35 sky130_fd_sc_hd__xor2_1
XTAP_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2905 net1225 net523 net1218 net796 VGND VGND VPWR VPWR t$5890 sky130_fd_sc_hd__a22o_1
XTAP_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2916 t$5895 net1368 VGND VGND VPWR VPWR booth_b42_m16 sky130_fd_sc_hd__xor2_1
XTAP_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2927 net1109 net523 net1101 net796 VGND VGND VPWR VPWR t$5901 sky130_fd_sc_hd__a22o_1
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_210 net1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_221 net1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2938 t$5906 net1371 VGND VGND VPWR VPWR booth_b42_m27 sky130_fd_sc_hd__xor2_1
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2949 net1002 net521 net994 net794 VGND VGND VPWR VPWR t$5912 sky130_fd_sc_hd__a22o_1
XFILLER_45_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_22_2 pp_row22_8 pp_row22_9 pp_row22_10 VGND VGND VPWR VPWR c$2018 s$2019
+ sky130_fd_sc_hd__fa_1
XANTENNA_232 net1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_243 net1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_254 net1619 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_265 net1723 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_276 c$4206 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_287 sel_1$5038 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_298 net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0790_ clknet_leaf_139_clk booth_b64_m26 VGND VGND VPWR VPWR pp_row90_20 sky130_fd_sc_hd__dfxtp_1
XU$$4477_1859 VGND VGND VPWR VPWR U$$4477_1859/HI net1859 sky130_fd_sc_hd__conb_1
XFILLER_10_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2460_ clknet_leaf_148_clk booth_b30_m38 VGND VGND VPWR VPWR pp_row68_14 sky130_fd_sc_hd__dfxtp_1
XFILLER_5_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1411_ clknet_leaf_41_clk booth_b30_m3 VGND VGND VPWR VPWR pp_row33_15 sky130_fd_sc_hd__dfxtp_1
X_2391_ clknet_leaf_128_clk booth_b58_m53 VGND VGND VPWR VPWR pp_row111_6 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_74_5 s$791 s$793 s$795 VGND VGND VPWR VPWR c$1624 s$1625 sky130_fd_sc_hd__fa_1
X_1342_ clknet_leaf_0_clk booth_b16_m14 VGND VGND VPWR VPWR pp_row30_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_96_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_67_4 s$659 s$661 s$663 VGND VGND VPWR VPWR c$1538 s$1539 sky130_fd_sc_hd__fa_1
XFILLER_69_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1273_ clknet_leaf_10_clk booth_b20_m6 VGND VGND VPWR VPWR pp_row26_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0224_ clknet_leaf_196_clk booth_b22_m49 VGND VGND VPWR VPWR pp_row71_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_0_68_0_1891 VGND VGND VPWR VPWR net1891 dadda_fa_0_68_0_1891/LO sky130_fd_sc_hd__conb_1
XFILLER_149_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4501_1871 VGND VGND VPWR VPWR U$$4501_1871/HI net1871 sky130_fd_sc_hd__conb_1
XFILLER_193_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0988_ clknet_leaf_181_clk net153 VGND VGND VPWR VPWR pp_row121_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_138_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_104_1 s$3315 s$3317 s$3319 VGND VGND VPWR VPWR c$3814 s$3815 sky130_fd_sc_hd__fa_1
XFILLER_106_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1609_ clknet_leaf_240_clk booth_b16_m26 VGND VGND VPWR VPWR pp_row42_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_154_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_62_3 pp_row62_26 pp_row62_27 pp_row62_28 VGND VGND VPWR VPWR c$570 s$571
+ sky130_fd_sc_hd__fa_1
XFILLER_170_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_55_2 pp_row55_11 pp_row55_12 pp_row55_13 VGND VGND VPWR VPWR c$442 s$443
+ sky130_fd_sc_hd__fa_1
Xdadda_fa_4_32_1 c$2090 c$2092 s$2095 VGND VGND VPWR VPWR c$2884 s$2885 sky130_fd_sc_hd__fa_1
XFILLER_27_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_48_1 pp_row48_3 pp_row48_4 pp_row48_5 VGND VGND VPWR VPWR c$318 s$319
+ sky130_fd_sc_hd__fa_1
XFILLER_28_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_25_0 s$1061 c$2030 c$2032 VGND VGND VPWR VPWR c$2840 s$2841 sky130_fd_sc_hd__fa_1
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_77_3 s$1655 s$1657 s$1659 VGND VGND VPWR VPWR c$2460 s$2461 sky130_fd_sc_hd__fa_1
XFILLER_3_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1601 net1602 VGND VGND VPWR VPWR net1601 sky130_fd_sc_hd__buf_2
Xfanout1612 net1614 VGND VGND VPWR VPWR net1612 sky130_fd_sc_hd__buf_4
XFILLER_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1623 net1627 VGND VGND VPWR VPWR net1623 sky130_fd_sc_hd__buf_4
Xfanout1634 net1636 VGND VGND VPWR VPWR net1634 sky130_fd_sc_hd__buf_4
Xfanout1645 net112 VGND VGND VPWR VPWR net1645 sky130_fd_sc_hd__buf_2
Xfanout1656 net110 VGND VGND VPWR VPWR net1656 sky130_fd_sc_hd__clkbuf_8
XFILLER_93_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4104 t$6501 net1285 VGND VGND VPWR VPWR booth_b58_m62 sky130_fd_sc_hd__xor2_1
XFILLER_144_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1667 net11 VGND VGND VPWR VPWR net1667 sky130_fd_sc_hd__buf_6
XU$$4115 net57 net1284 VGND VGND VPWR VPWR sel_1$6508 sky130_fd_sc_hd__xor2_1
Xfanout680 net681 VGND VGND VPWR VPWR net680 sky130_fd_sc_hd__clkbuf_4
XU$$4126 net1677 net438 net1566 net720 VGND VGND VPWR VPWR t$6514 sky130_fd_sc_hd__a22o_1
Xfanout1678 net109 VGND VGND VPWR VPWR net1678 sky130_fd_sc_hd__buf_6
Xfanout1689 net107 VGND VGND VPWR VPWR net1689 sky130_fd_sc_hd__buf_4
XU$$4137 t$6519 net1264 VGND VGND VPWR VPWR booth_b60_m10 sky130_fd_sc_hd__xor2_1
Xfanout691 net692 VGND VGND VPWR VPWR net691 sky130_fd_sc_hd__buf_6
XU$$4148 net1168 net434 net1159 net716 VGND VGND VPWR VPWR t$6525 sky130_fd_sc_hd__a22o_1
Xdadda_ha_3_14_0 pp_row14_0 pp_row14_1 VGND VGND VPWR VPWR c$1974 s$1975 sky130_fd_sc_hd__ha_1
XU$$3403 t$6143 net1345 VGND VGND VPWR VPWR booth_b48_m54 sky130_fd_sc_hd__xor2_1
XU$$4159 t$6530 net1263 VGND VGND VPWR VPWR booth_b60_m21 sky130_fd_sc_hd__xor2_1
XU$$3414 net1583 net499 net1556 net772 VGND VGND VPWR VPWR t$6149 sky130_fd_sc_hd__a22o_1
XU$$3425 net1342 VGND VGND VPWR VPWR notblock$6155\[0\] sky130_fd_sc_hd__inv_1
XU$$3436 t$6161 net1333 VGND VGND VPWR VPWR booth_b50_m2 sky130_fd_sc_hd__xor2_1
XFILLER_19_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2702 t$5785 net1396 VGND VGND VPWR VPWR booth_b38_m46 sky130_fd_sc_hd__xor2_1
XU$$3447 net1514 net487 net1506 net760 VGND VGND VPWR VPWR t$6167 sky130_fd_sc_hd__a22o_1
XTAP_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3458 t$6172 net1329 VGND VGND VPWR VPWR booth_b50_m13 sky130_fd_sc_hd__xor2_1
XU$$2713 net1651 net548 net1643 net821 VGND VGND VPWR VPWR t$5791 sky130_fd_sc_hd__a22o_1
XU$$2724 t$5796 net1400 VGND VGND VPWR VPWR booth_b38_m57 sky130_fd_sc_hd__xor2_1
XU$$3469 net1145 net488 net1137 net761 VGND VGND VPWR VPWR t$6178 sky130_fd_sc_hd__a22o_1
XFILLER_61_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2735 net1542 net547 net1534 net820 VGND VGND VPWR VPWR t$5802 sky130_fd_sc_hd__a22o_1
XTAP_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2746 net1782 net535 net1227 net808 VGND VGND VPWR VPWR t$5809 sky130_fd_sc_hd__a22o_1
XTAP_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2757 t$5814 net1377 VGND VGND VPWR VPWR booth_b40_m5 sky130_fd_sc_hd__xor2_1
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2768 net1225 net539 net1218 net812 VGND VGND VPWR VPWR t$5820 sky130_fd_sc_hd__a22o_1
XU$$2779 t$5825 net1381 VGND VGND VPWR VPWR booth_b40_m16 sky130_fd_sc_hd__xor2_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1960_ clknet_leaf_64_clk booth_b24_m30 VGND VGND VPWR VPWR pp_row54_12 sky130_fd_sc_hd__dfxtp_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0911_ clknet_leaf_104_clk booth_b48_m48 VGND VGND VPWR VPWR pp_row96_9 sky130_fd_sc_hd__dfxtp_1
X_1891_ clknet_leaf_39_clk booth_b14_m38 VGND VGND VPWR VPWR pp_row52_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_187_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0842_ clknet_leaf_106_clk booth_b36_m57 VGND VGND VPWR VPWR pp_row93_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_146_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0773_ clknet_leaf_144_clk booth_b34_m56 VGND VGND VPWR VPWR pp_row90_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2443_ clknet_leaf_97_clk booth_b64_m3 VGND VGND VPWR VPWR pp_row67_32 sky130_fd_sc_hd__dfxtp_1
XFILLER_103_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_72_2 c$736 c$738 c$740 VGND VGND VPWR VPWR c$1594 s$1595 sky130_fd_sc_hd__fa_2
XFILLER_130_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2374_ clknet_leaf_84_clk booth_b8_m58 VGND VGND VPWR VPWR pp_row66_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_65_1 c$604 c$606 c$608 VGND VGND VPWR VPWR c$1508 s$1509 sky130_fd_sc_hd__fa_2
X_1325_ clknet_leaf_1_clk booth_b18_m11 VGND VGND VPWR VPWR pp_row29_9 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$708 final_adder.p_new$732 final_adder.p_new$716 VGND VGND VPWR VPWR
+ final_adder.p_new$836 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$719 final_adder.p_new$726 final_adder.g_new$743 final_adder.g_new$727
+ VGND VGND VPWR VPWR final_adder.g_new$847 sky130_fd_sc_hd__a21o_1
Xdadda_fa_5_42_0 c$2936 c$2938 c$2940 VGND VGND VPWR VPWR c$3564 s$3565 sky130_fd_sc_hd__fa_1
XFILLER_69_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_58_0 s$31 c$474 c$476 VGND VGND VPWR VPWR c$1422 s$1423 sky130_fd_sc_hd__fa_1
XFILLER_151_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1256_ clknet_leaf_11_clk booth_b18_m7 VGND VGND VPWR VPWR pp_row25_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_83_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0207_ clknet_leaf_152_clk booth_b54_m16 VGND VGND VPWR VPWR pp_row70_25 sky130_fd_sc_hd__dfxtp_1
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1187_ clknet_leaf_49_clk booth_b0_m21 VGND VGND VPWR VPWR pp_row21_0 sky130_fd_sc_hd__dfxtp_1
XU$$3970 net1529 net462 net1800 net735 VGND VGND VPWR VPWR t$6433 sky130_fd_sc_hd__a22o_1
XFILLER_80_832 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3981 net1233 net451 net1129 net724 VGND VGND VPWR VPWR t$6440 sky130_fd_sc_hd__a22o_1
XU$$3992 t$6445 net1287 VGND VGND VPWR VPWR booth_b58_m6 sky130_fd_sc_hd__xor2_1
XFILLER_52_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_606 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4499_1870 VGND VGND VPWR VPWR U$$4499_1870/HI net1870 sky130_fd_sc_hd__conb_1
XFILLER_193_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_672 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_87_2 s$2537 s$2539 s$2541 VGND VGND VPWR VPWR c$3216 s$3217 sky130_fd_sc_hd__fa_1
XFILLER_160_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput261 net261 VGND VGND VPWR VPWR o[103] sky130_fd_sc_hd__buf_2
Xdadda_fa_7_57_0 s$3627 c$4008 s$4011 VGND VGND VPWR VPWR c$4266 s$4267 sky130_fd_sc_hd__fa_1
XFILLER_133_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput272 net272 VGND VGND VPWR VPWR o[113] sky130_fd_sc_hd__buf_2
Xoutput283 net283 VGND VGND VPWR VPWR o[123] sky130_fd_sc_hd__buf_2
XFILLER_160_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput294 net294 VGND VGND VPWR VPWR o[18] sky130_fd_sc_hd__buf_2
XFILLER_87_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_60_0 pp_row60_14 pp_row60_15 pp_row60_16 VGND VGND VPWR VPWR c$528 s$529
+ sky130_fd_sc_hd__fa_1
XFILLER_101_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2009 t$5431 net1455 VGND VGND VPWR VPWR booth_b28_m42 sky130_fd_sc_hd__xor2_1
XFILLER_71_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1308 t$5073 net1665 VGND VGND VPWR VPWR booth_b18_m34 sky130_fd_sc_hd__xor2_1
XFILLER_15_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1319 net944 net639 net928 net912 VGND VGND VPWR VPWR t$5079 sky130_fd_sc_hd__a22o_1
XFILLER_70_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_82_1 c$1702 c$1704 c$1706 VGND VGND VPWR VPWR c$2496 s$2497 sky130_fd_sc_hd__fa_1
XFILLER_139_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_75_0 s$815 c$1614 c$1616 VGND VGND VPWR VPWR c$2438 s$2439 sky130_fd_sc_hd__fa_1
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1420 net1422 VGND VGND VPWR VPWR net1420 sky130_fd_sc_hd__buf_6
Xfanout1431 net1438 VGND VGND VPWR VPWR net1431 sky130_fd_sc_hd__buf_8
XFILLER_79_976 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1442 net1443 VGND VGND VPWR VPWR net1442 sky130_fd_sc_hd__buf_8
Xfanout1453 net1454 VGND VGND VPWR VPWR net1453 sky130_fd_sc_hd__buf_6
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1464 net1465 VGND VGND VPWR VPWR net1464 sky130_fd_sc_hd__buf_8
Xfanout1475 net1477 VGND VGND VPWR VPWR net1475 sky130_fd_sc_hd__buf_6
X_1110_ clknet_leaf_13_clk booth_b14_m0 VGND VGND VPWR VPWR pp_row14_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_120_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1486 net1490 VGND VGND VPWR VPWR net1486 sky130_fd_sc_hd__buf_6
XFILLER_94_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3200 t$6040 net1353 VGND VGND VPWR VPWR booth_b46_m21 sky130_fd_sc_hd__xor2_1
X_2090_ clknet_leaf_37_clk booth_b18_m40 VGND VGND VPWR VPWR pp_row58_9 sky130_fd_sc_hd__dfxtp_1
Xfanout1497 net1498 VGND VGND VPWR VPWR net1497 sky130_fd_sc_hd__buf_2
XFILLER_171_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3211 net1065 net501 net1059 net774 VGND VGND VPWR VPWR t$6046 sky130_fd_sc_hd__a22o_1
XU$$3222 t$6051 net1351 VGND VGND VPWR VPWR booth_b46_m32 sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_111_1 c$2720 c$2722 c$2724 VGND VGND VPWR VPWR c$3358 s$3359 sky130_fd_sc_hd__fa_1
X_1041_ clknet_leaf_57_clk booth_b2_m4 VGND VGND VPWR VPWR pp_row6_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_150_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3233 net959 net503 net950 net776 VGND VGND VPWR VPWR t$6057 sky130_fd_sc_hd__a22o_1
XFILLER_24_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3244 t$6062 net1350 VGND VGND VPWR VPWR booth_b46_m43 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$15 c$4180 s$4183 VGND VGND VPWR VPWR final_adder.$signal$32 final_adder.$signal$1105
+ sky130_fd_sc_hd__ha_1
XU$$3255 net1691 net505 net1683 net778 VGND VGND VPWR VPWR t$6068 sky130_fd_sc_hd__a22o_1
XU$$2510 net1144 net554 net1134 net827 VGND VGND VPWR VPWR t$5688 sky130_fd_sc_hd__a22o_1
XFILLER_34_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$26 c$4202 s$4205 VGND VGND VPWR VPWR final_adder.$signal$54 final_adder.$signal$1116
+ sky130_fd_sc_hd__ha_2
Xdadda_fa_4_104_0 s$1961 c$2662 c$2664 VGND VGND VPWR VPWR c$3314 s$3315 sky130_fd_sc_hd__fa_1
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_37_5 c$208 c$210 s$213 VGND VGND VPWR VPWR c$1180 s$1181 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$37 c$4224 s$4227 VGND VGND VPWR VPWR final_adder.$signal$76 final_adder.$signal$1127
+ sky130_fd_sc_hd__ha_1
XU$$3266 t$6073 net1355 VGND VGND VPWR VPWR booth_b46_m54 sky130_fd_sc_hd__xor2_1
XU$$2521 t$5693 net1405 VGND VGND VPWR VPWR booth_b36_m24 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$48 c$4246 s$4249 VGND VGND VPWR VPWR final_adder.$signal$98 final_adder.$signal$1138
+ sky130_fd_sc_hd__ha_1
XU$$2532 net1046 net559 net1030 net832 VGND VGND VPWR VPWR t$5699 sky130_fd_sc_hd__a22o_1
XU$$3277 net1583 net508 net1556 net781 VGND VGND VPWR VPWR t$6079 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$59 c$4268 s$4271 VGND VGND VPWR VPWR final_adder.$signal$120 final_adder.$signal$1149
+ sky130_fd_sc_hd__ha_1
XU$$2543 t$5704 net1409 VGND VGND VPWR VPWR booth_b36_m35 sky130_fd_sc_hd__xor2_1
XU$$3288 net1350 VGND VGND VPWR VPWR notblock$6085\[0\] sky130_fd_sc_hd__inv_1
XFILLER_34_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2554 net927 net555 net1746 net828 VGND VGND VPWR VPWR t$5710 sky130_fd_sc_hd__a22o_1
XU$$3299 t$6091 net1339 VGND VGND VPWR VPWR booth_b48_m2 sky130_fd_sc_hd__xor2_1
XU$$1820 t$5335 net1457 VGND VGND VPWR VPWR booth_b26_m16 sky130_fd_sc_hd__xor2_1
XU$$2565 t$5715 net1408 VGND VGND VPWR VPWR booth_b36_m46 sky130_fd_sc_hd__xor2_1
XFILLER_55_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1831 net1107 net595 net1098 net868 VGND VGND VPWR VPWR t$5341 sky130_fd_sc_hd__a22o_1
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2576 net1648 net556 net1640 net829 VGND VGND VPWR VPWR t$5721 sky130_fd_sc_hd__a22o_1
XU$$2587 t$5726 net1410 VGND VGND VPWR VPWR booth_b36_m57 sky130_fd_sc_hd__xor2_1
XU$$1842 t$5346 net1461 VGND VGND VPWR VPWR booth_b26_m27 sky130_fd_sc_hd__xor2_1
XU$$2598 net1542 net558 net1534 net831 VGND VGND VPWR VPWR t$5732 sky130_fd_sc_hd__a22o_1
XFILLER_21_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1853 net999 net597 net991 net870 VGND VGND VPWR VPWR t$5352 sky130_fd_sc_hd__a22o_1
XU$$1864 t$5357 net1462 VGND VGND VPWR VPWR booth_b26_m38 sky130_fd_sc_hd__xor2_1
XU$$1875 net1733 net600 net1724 net873 VGND VGND VPWR VPWR t$5363 sky130_fd_sc_hd__a22o_1
XU$$1886 t$5368 net1464 VGND VGND VPWR VPWR booth_b26_m49 sky130_fd_sc_hd__xor2_1
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1943_ clknet_leaf_72_clk booth_b50_m3 VGND VGND VPWR VPWR pp_row53_25 sky130_fd_sc_hd__dfxtp_1
XU$$1897 net1622 net599 net1613 net872 VGND VGND VPWR VPWR t$5374 sky130_fd_sc_hd__a22o_1
XFILLER_175_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1874_ clknet_leaf_69_clk booth_b36_m15 VGND VGND VPWR VPWR pp_row51_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_174_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_97_1 s$3273 s$3275 s$3277 VGND VGND VPWR VPWR c$3786 s$3787 sky130_fd_sc_hd__fa_1
X_0825_ clknet_leaf_109_clk booth_b46_m46 VGND VGND VPWR VPWR pp_row92_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_128_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0756_ clknet_leaf_161_clk booth_b44_m45 VGND VGND VPWR VPWR pp_row89_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_143_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0687_ clknet_leaf_168_clk booth_b56_m30 VGND VGND VPWR VPWR pp_row86_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_66_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2426_ clknet_leaf_98_clk booth_b32_m35 VGND VGND VPWR VPWR pp_row67_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_9_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2357_ clknet_leaf_75_clk booth_b44_m21 VGND VGND VPWR VPWR pp_row65_22 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$505 final_adder.p_new$506 final_adder.g_new$383 final_adder.g_new$507
+ VGND VGND VPWR VPWR final_adder.g_new$633 sky130_fd_sc_hd__a21o_4
XFILLER_57_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$516 final_adder.p_new$528 final_adder.p_new$520 VGND VGND VPWR VPWR
+ final_adder.p_new$644 sky130_fd_sc_hd__and2_1
XFILLER_69_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$527 final_adder.p_new$530 final_adder.g_new$539 final_adder.g_new$531
+ VGND VGND VPWR VPWR final_adder.g_new$655 sky130_fd_sc_hd__a21o_1
XTAP_3809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1308_ clknet_leaf_1_clk booth_b20_m8 VGND VGND VPWR VPWR pp_row28_10 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$538 final_adder.p_new$550 final_adder.p_new$542 VGND VGND VPWR VPWR
+ final_adder.p_new$666 sky130_fd_sc_hd__and2_1
XFILLER_38_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2288_ clknet_leaf_210_clk booth_b50_m13 VGND VGND VPWR VPWR pp_row63_25 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$549 final_adder.p_new$552 final_adder.g_new$561 final_adder.g_new$553
+ VGND VGND VPWR VPWR final_adder.g_new$677 sky130_fd_sc_hd__a21o_1
XFILLER_38_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1239_ clknet_leaf_13_clk booth_b16_m8 VGND VGND VPWR VPWR pp_row24_8 sky130_fd_sc_hd__dfxtp_1
XU$$4490 net1685 sel_0$6647 net1659 net697 VGND VGND VPWR VPWR t$6699 sky130_fd_sc_hd__a22o_1
XFILLER_52_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1081 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_92_0 s$1841 c$2566 c$2568 VGND VGND VPWR VPWR c$3242 s$3243 sky130_fd_sc_hd__fa_1
XFILLER_165_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_106_2 pp_row106_11 pp_row106_12 pp_row106_13 VGND VGND VPWR VPWR c$2690
+ s$2691 sky130_fd_sc_hd__fa_2
XFILLER_118_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$900 net973 net394 net964 net660 VGND VGND VPWR VPWR t$4865 sky130_fd_sc_hd__a22o_1
XFILLER_75_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$911 t$4870 net1314 VGND VGND VPWR VPWR booth_b12_m41 sky130_fd_sc_hd__xor2_1
XFILLER_28_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$922 net1705 net395 net1697 net661 VGND VGND VPWR VPWR t$4876 sky130_fd_sc_hd__a22o_1
XFILLER_29_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$933 t$4881 net1318 VGND VGND VPWR VPWR booth_b12_m52 sky130_fd_sc_hd__xor2_1
XU$$944 net1599 net399 net1590 net665 VGND VGND VPWR VPWR t$4887 sky130_fd_sc_hd__a22o_1
XU$$955 t$4892 net1316 VGND VGND VPWR VPWR booth_b12_m63 sky130_fd_sc_hd__xor2_1
XU$$1105 t$4970 net1006 VGND VGND VPWR VPWR booth_b16_m1 sky130_fd_sc_hd__xor2_1
XU$$966 t$4899 net1185 VGND VGND VPWR VPWR booth_b14_m0 sky130_fd_sc_hd__xor2_1
XU$$1116 net1521 net646 net1513 net919 VGND VGND VPWR VPWR t$4976 sky130_fd_sc_hd__a22o_1
XU$$977 net1564 net389 net1523 net655 VGND VGND VPWR VPWR t$4905 sky130_fd_sc_hd__a22o_1
XU$$1127 t$4981 net1006 VGND VGND VPWR VPWR booth_b16_m12 sky130_fd_sc_hd__xor2_1
XU$$988 t$4910 net1184 VGND VGND VPWR VPWR booth_b14_m11 sky130_fd_sc_hd__xor2_1
XU$$999 net1155 net385 net1146 net651 VGND VGND VPWR VPWR t$4916 sky130_fd_sc_hd__a22o_1
XU$$1138 net1149 net646 net1143 net919 VGND VGND VPWR VPWR t$4987 sky130_fd_sc_hd__a22o_1
XU$$1149 t$4992 net1008 VGND VGND VPWR VPWR booth_b16_m23 sky130_fd_sc_hd__xor2_1
XFILLER_71_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1034 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0610_ clknet_leaf_181_clk net147 VGND VGND VPWR VPWR pp_row116_8 sky130_fd_sc_hd__dfxtp_2
X_1590_ clknet_leaf_9_clk booth_b26_m15 VGND VGND VPWR VPWR pp_row41_13 sky130_fd_sc_hd__dfxtp_1
XFILLER_171_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0541_ clknet_leaf_169_clk booth_b34_m47 VGND VGND VPWR VPWR pp_row81_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_113_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0472_ clknet_leaf_193_clk notsign$4964 VGND VGND VPWR VPWR pp_row79_0 sky130_fd_sc_hd__dfxtp_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4116_1805 VGND VGND VPWR VPWR U$$4116_1805/HI net1805 sky130_fd_sc_hd__conb_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2211_ clknet_leaf_212_clk booth_b44_m17 VGND VGND VPWR VPWR pp_row61_22 sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1250 net1252 VGND VGND VPWR VPWR net1250 sky130_fd_sc_hd__buf_6
XFILLER_38_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1261 net1262 VGND VGND VPWR VPWR net1261 sky130_fd_sc_hd__buf_6
Xdadda_ha_2_29_3 pp_row29_9 pp_row29_10 VGND VGND VPWR VPWR c$1088 s$1089 sky130_fd_sc_hd__ha_1
X_2142_ clknet_leaf_219_clk booth_b48_m11 VGND VGND VPWR VPWR pp_row59_24 sky130_fd_sc_hd__dfxtp_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1272 net58 VGND VGND VPWR VPWR net1272 sky130_fd_sc_hd__buf_4
XFILLER_66_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1283 net55 VGND VGND VPWR VPWR net1283 sky130_fd_sc_hd__clkbuf_4
Xfanout1294 net1295 VGND VGND VPWR VPWR net1294 sky130_fd_sc_hd__buf_6
XFILLER_94_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_42_3 pp_row42_23 c$236 c$238 VGND VGND VPWR VPWR c$1236 s$1237 sky130_fd_sc_hd__fa_1
X_2073_ clknet_leaf_32_clk booth_b46_m11 VGND VGND VPWR VPWR pp_row57_23 sky130_fd_sc_hd__dfxtp_1
XU$$3030 net1674 net510 net1563 net783 VGND VGND VPWR VPWR t$5954 sky130_fd_sc_hd__a22o_1
XU$$3041 t$5959 net1362 VGND VGND VPWR VPWR booth_b44_m10 sky130_fd_sc_hd__xor2_1
XU$$3052 net1165 net510 net1156 net783 VGND VGND VPWR VPWR t$5965 sky130_fd_sc_hd__a22o_1
XU$$3063 t$5970 net1362 VGND VGND VPWR VPWR booth_b44_m21 sky130_fd_sc_hd__xor2_1
X_1024_ clknet_leaf_60_clk net1391 VGND VGND VPWR VPWR pp_row2_2 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_35_2 pp_row35_8 pp_row35_9 pp_row35_10 VGND VGND VPWR VPWR c$1150 s$1151
+ sky130_fd_sc_hd__fa_1
XU$$3074 net1068 net511 net1060 net784 VGND VGND VPWR VPWR t$5976 sky130_fd_sc_hd__a22o_1
XU$$2340 t$5601 net1423 VGND VGND VPWR VPWR booth_b34_m2 sky130_fd_sc_hd__xor2_1
XU$$3085 t$5981 net1359 VGND VGND VPWR VPWR booth_b44_m32 sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_12_1 s$2763 s$2765 s$2767 VGND VGND VPWR VPWR c$3446 s$3447 sky130_fd_sc_hd__fa_1
XU$$3096 net959 net512 net950 net785 VGND VGND VPWR VPWR t$5987 sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_28_1 pp_row28_3 pp_row28_4 pp_row28_5 VGND VGND VPWR VPWR c$1076 s$1077
+ sky130_fd_sc_hd__fa_1
XU$$2351 net1512 net560 net1504 net833 VGND VGND VPWR VPWR t$5607 sky130_fd_sc_hd__a22o_1
XU$$2362 t$5612 net1420 VGND VGND VPWR VPWR booth_b34_m13 sky130_fd_sc_hd__xor2_1
XU$$2373 net1144 net563 net1134 net836 VGND VGND VPWR VPWR t$5618 sky130_fd_sc_hd__a22o_1
XFILLER_50_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2384 t$5623 net1421 VGND VGND VPWR VPWR booth_b34_m24 sky130_fd_sc_hd__xor2_1
XU$$1650 net1765 net603 net1228 net876 VGND VGND VPWR VPWR t$5249 sky130_fd_sc_hd__a22o_1
XU$$2395 net1042 net562 net1026 net835 VGND VGND VPWR VPWR t$5629 sky130_fd_sc_hd__a22o_1
XU$$1661 t$5254 net1466 VGND VGND VPWR VPWR booth_b24_m5 sky130_fd_sc_hd__xor2_1
XU$$1672 net1225 net605 net1216 net878 VGND VGND VPWR VPWR t$5260 sky130_fd_sc_hd__a22o_1
XFILLER_22_559 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1683 t$5265 net1467 VGND VGND VPWR VPWR booth_b24_m16 sky130_fd_sc_hd__xor2_1
XU$$1694 net1107 net603 net1098 net876 VGND VGND VPWR VPWR t$5271 sky130_fd_sc_hd__a22o_1
XFILLER_188_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1926_ clknet_leaf_65_clk booth_b20_m33 VGND VGND VPWR VPWR pp_row53_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_187_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1857_ clknet_leaf_79_clk booth_b6_m45 VGND VGND VPWR VPWR pp_row51_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0808_ clknet_leaf_101_clk booth_b56_m35 VGND VGND VPWR VPWR pp_row91_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_146_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1788_ clknet_leaf_220_clk booth_b44_m4 VGND VGND VPWR VPWR pp_row48_22 sky130_fd_sc_hd__dfxtp_1
XFILLER_104_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1052 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0739_ clknet_leaf_163_clk booth_b58_m30 VGND VGND VPWR VPWR pp_row88_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_118_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2409_ clknet_leaf_84_clk notsign$4544 VGND VGND VPWR VPWR pp_row67_1 sky130_fd_sc_hd__dfxtp_1
XTAP_4307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$302 final_adder.p_new$304 final_adder.p_new$302 VGND VGND VPWR VPWR
+ final_adder.p_new$430 sky130_fd_sc_hd__and2_1
XTAP_4329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$313 final_adder.p_new$312 final_adder.g_new$315 final_adder.g_new$313
+ VGND VGND VPWR VPWR final_adder.g_new$441 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$324 final_adder.p_new$326 final_adder.p_new$324 VGND VGND VPWR VPWR
+ final_adder.p_new$452 sky130_fd_sc_hd__and2_1
XTAP_3606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$335 final_adder.p_new$334 final_adder.g_new$337 final_adder.g_new$335
+ VGND VGND VPWR VPWR final_adder.g_new$463 sky130_fd_sc_hd__a21o_1
XTAP_3617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$346 final_adder.p_new$348 final_adder.p_new$346 VGND VGND VPWR VPWR
+ final_adder.p_new$474 sky130_fd_sc_hd__and2_1
XTAP_3628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$357 final_adder.p_new$356 final_adder.g_new$359 final_adder.g_new$357
+ VGND VGND VPWR VPWR final_adder.g_new$485 sky130_fd_sc_hd__a21o_1
XTAP_3639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$207 net1017 net623 net1000 net896 VGND VGND VPWR VPWR t$4511 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$368 final_adder.p_new$370 final_adder.p_new$368 VGND VGND VPWR VPWR
+ final_adder.p_new$496 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$379 final_adder.p_new$378 final_adder.g_new$381 final_adder.g_new$379
+ VGND VGND VPWR VPWR final_adder.g_new$507 sky130_fd_sc_hd__a21o_1
XFILLER_55_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$218 t$4516 net1391 VGND VGND VPWR VPWR booth_b2_m37 sky130_fd_sc_hd__xor2_1
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$229 net1738 net622 net1730 net895 VGND VGND VPWR VPWR t$4522 sky130_fd_sc_hd__a22o_1
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_111_0 pp_row111_0 pp_row111_1 pp_row111_2 VGND VGND VPWR VPWR c$2726 s$2727
+ sky130_fd_sc_hd__fa_1
XFILLER_4_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_52_2 c$1348 s$1351 s$1353 VGND VGND VPWR VPWR c$2258 s$2259 sky130_fd_sc_hd__fa_1
Xdadda_fa_0_68_2 pp_row68_6 pp_row68_7 pp_row68_8 VGND VGND VPWR VPWR c$136 s$137
+ sky130_fd_sc_hd__fa_1
Xdadda_fa_3_45_1 c$1258 c$1260 c$1262 VGND VGND VPWR VPWR c$2200 s$2201 sky130_fd_sc_hd__fa_1
XFILLER_64_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_22_0 c$3480 c$3482 s$3485 VGND VGND VPWR VPWR c$3940 s$3941 sky130_fd_sc_hd__fa_1
Xdadda_fa_3_38_0 s$221 c$1170 c$1172 VGND VGND VPWR VPWR c$2142 s$2143 sky130_fd_sc_hd__fa_1
XFILLER_90_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$891 final_adder.p_new$922 final_adder.g_new$631 final_adder.g_new$923
+ VGND VGND VPWR VPWR final_adder.g_new$1019 sky130_fd_sc_hd__a21o_1
XU$$730 t$4778 net1412 VGND VGND VPWR VPWR booth_b10_m19 sky130_fd_sc_hd__xor2_1
XFILLER_28_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$741 net1084 net404 net1075 net670 VGND VGND VPWR VPWR t$4784 sky130_fd_sc_hd__a22o_1
XFILLER_1_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$752 t$4789 net1412 VGND VGND VPWR VPWR booth_b10_m30 sky130_fd_sc_hd__xor2_1
XU$$763 net973 net401 net964 net667 VGND VGND VPWR VPWR t$4795 sky130_fd_sc_hd__a22o_1
XU$$774 t$4800 net1416 VGND VGND VPWR VPWR booth_b10_m41 sky130_fd_sc_hd__xor2_1
XFILLER_32_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$785 net1706 net405 net1698 net671 VGND VGND VPWR VPWR t$4806 sky130_fd_sc_hd__a22o_1
XU$$796 t$4811 net1418 VGND VGND VPWR VPWR booth_b10_m52 sky130_fd_sc_hd__xor2_1
XFILLER_188_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1711_ clknet_leaf_237_clk booth_b8_m38 VGND VGND VPWR VPWR pp_row46_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_185_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$143_1761 VGND VGND VPWR VPWR U$$143_1761/HI net1761 sky130_fd_sc_hd__conb_1
XANTENNA_2 c$1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1642_ clknet_leaf_240_clk booth_b26_m17 VGND VGND VPWR VPWR pp_row43_13 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_97_4 pp_row97_12 pp_row97_13 pp_row97_14 VGND VGND VPWR VPWR c$1898 s$1899
+ sky130_fd_sc_hd__fa_1
XFILLER_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_110_0_1909 VGND VGND VPWR VPWR net1909 dadda_fa_3_110_0_1909/LO sky130_fd_sc_hd__conb_1
XFILLER_99_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1573_ clknet_leaf_21_clk booth_b40_m0 VGND VGND VPWR VPWR pp_row40_20 sky130_fd_sc_hd__dfxtp_1
XFILLER_141_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0524_ clknet_leaf_167_clk booth_b54_m26 VGND VGND VPWR VPWR pp_row80_20 sky130_fd_sc_hd__dfxtp_1
Xfanout509 sel_0$6017 VGND VGND VPWR VPWR net509 sky130_fd_sc_hd__buf_4
XFILLER_112_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0455_ clknet_leaf_131_clk booth_b54_m61 VGND VGND VPWR VPWR pp_row115_2 sky130_fd_sc_hd__dfxtp_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0386_ clknet_leaf_195_clk booth_b24_m52 VGND VGND VPWR VPWR pp_row76_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1057 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1080 net1081 VGND VGND VPWR VPWR net1080 sky130_fd_sc_hd__buf_4
XFILLER_66_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1091 net1092 VGND VGND VPWR VPWR net1091 sky130_fd_sc_hd__clkbuf_8
XFILLER_55_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2125_ clknet_leaf_217_clk booth_b18_m41 VGND VGND VPWR VPWR pp_row59_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_82_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_40_0 pp_row40_11 pp_row40_12 pp_row40_13 VGND VGND VPWR VPWR c$1206 s$1207
+ sky130_fd_sc_hd__fa_1
XFILLER_187_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2056_ clknet_leaf_38_clk booth_b18_m39 VGND VGND VPWR VPWR pp_row57_9 sky130_fd_sc_hd__dfxtp_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1007_ clknet_leaf_119_clk booth_b54_m47 VGND VGND VPWR VPWR pp_row101_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_35_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2170 t$5513 net1444 VGND VGND VPWR VPWR booth_b30_m54 sky130_fd_sc_hd__xor2_1
XU$$2181 net1580 net579 net1554 net852 VGND VGND VPWR VPWR t$5519 sky130_fd_sc_hd__a22o_1
XU$$2192 net1444 VGND VGND VPWR VPWR notblock$5525\[0\] sky130_fd_sc_hd__inv_1
XFILLER_22_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1480 net1646 net632 net1640 net905 VGND VGND VPWR VPWR t$5161 sky130_fd_sc_hd__a22o_1
XU$$1491 t$5166 net1492 VGND VGND VPWR VPWR booth_b20_m57 sky130_fd_sc_hd__xor2_1
XFILLER_50_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1909_ clknet_leaf_70_clk booth_b46_m6 VGND VGND VPWR VPWR pp_row52_23 sky130_fd_sc_hd__dfxtp_1
XFILLER_108_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_85_2 pp_row85_6 pp_row85_7 pp_row85_8 VGND VGND VPWR VPWR c$970 s$971
+ sky130_fd_sc_hd__fa_2
XFILLER_132_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_62_1 c$2330 c$2332 s$2335 VGND VGND VPWR VPWR c$3064 s$3065 sky130_fd_sc_hd__fa_1
Xdadda_fa_1_78_1 pp_row78_5 pp_row78_6 pp_row78_7 VGND VGND VPWR VPWR c$854 s$855
+ sky130_fd_sc_hd__fa_1
XFILLER_77_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_55_0 s$1397 c$2270 c$2272 VGND VGND VPWR VPWR c$3020 s$3021 sky130_fd_sc_hd__fa_1
XTAP_4104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$110 c$4370 s$4373 VGND VGND VPWR VPWR final_adder.$signal$222 final_adder.$signal$1200
+ sky130_fd_sc_hd__ha_1
XTAP_4137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$121 c$4392 s$4395 VGND VGND VPWR VPWR final_adder.$signal$244 final_adder.$signal$1211
+ sky130_fd_sc_hd__ha_2
XTAP_4148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$132 final_adder.$signal$1212 final_adder.$signal$1213 VGND VGND VPWR
+ VPWR final_adder.p_new$260 sky130_fd_sc_hd__and2_1
XTAP_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$143 final_adder.$signal$1203 final_adder.$signal$226 final_adder.$signal$228
+ VGND VGND VPWR VPWR final_adder.g_new$271 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$154 final_adder.$signal$1190 final_adder.$signal$1191 VGND VGND VPWR
+ VPWR final_adder.p_new$282 sky130_fd_sc_hd__and2_1
XTAP_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$165 final_adder.$signal$1181 final_adder.$signal$182 final_adder.$signal$184
+ VGND VGND VPWR VPWR final_adder.g_new$293 sky130_fd_sc_hd__a21o_1
XTAP_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_990 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$176 final_adder.$signal$1168 final_adder.$signal$1169 VGND VGND VPWR
+ VPWR final_adder.p_new$304 sky130_fd_sc_hd__and2_1
XTAP_3458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_403 net1667 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$187 final_adder.$signal$1159 final_adder.$signal$138 final_adder.$signal$140
+ VGND VGND VPWR VPWR final_adder.g_new$315 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$198 final_adder.$signal$1146 final_adder.$signal$1147 VGND VGND VPWR
+ VPWR final_adder.p_new$326 sky130_fd_sc_hd__and2_1
XTAP_3469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_414 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_425 net601 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_436 net854 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_447 net1502 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_458 net1640 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_0_74_2 pp_row74_6 pp_row74_7 VGND VGND VPWR VPWR c$190 s$191 sky130_fd_sc_hd__ha_1
XFILLER_154_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_73_0 pp_row73_0 pp_row73_1 pp_row73_2 VGND VGND VPWR VPWR c$180 s$181
+ sky130_fd_sc_hd__fa_1
XFILLER_49_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0240_ clknet_leaf_150_clk booth_b52_m19 VGND VGND VPWR VPWR pp_row71_23 sky130_fd_sc_hd__dfxtp_1
Xinput150 c[119] VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_1
Xinput161 c[13] VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_1
Xinput172 c[23] VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0171_ clknet_leaf_97_clk booth_b50_m19 VGND VGND VPWR VPWR pp_row69_23 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_196_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_196_clk
+ sky130_fd_sc_hd__clkbuf_16
Xinput183 c[33] VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_1
Xinput194 c[43] VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_1
XTAP_3970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$560 net1036 net414 net936 net680 VGND VGND VPWR VPWR t$4692 sky130_fd_sc_hd__a22o_1
XFILLER_17_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$571 t$4697 net1236 VGND VGND VPWR VPWR booth_b8_m8 sky130_fd_sc_hd__xor2_1
XU$$582 net1198 net413 net1179 net679 VGND VGND VPWR VPWR t$4703 sky130_fd_sc_hd__a22o_1
XU$$593 t$4708 net1235 VGND VGND VPWR VPWR booth_b8_m19 sky130_fd_sc_hd__xor2_1
XFILLER_147_1051 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_120_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_120_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_172_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_95_1 pp_row95_6 pp_row95_7 pp_row95_8 VGND VGND VPWR VPWR c$1868 s$1869
+ sky130_fd_sc_hd__fa_1
XFILLER_133_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1625_ clknet_leaf_239_clk net1367 VGND VGND VPWR VPWR pp_row42_22 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_72_0 c$3116 c$3118 c$3120 VGND VGND VPWR VPWR c$3684 s$3685 sky130_fd_sc_hd__fa_1
Xdadda_fa_2_88_0 pp_row88_14 pp_row88_15 pp_row88_16 VGND VGND VPWR VPWR c$1782 s$1783
+ sky130_fd_sc_hd__fa_1
XFILLER_141_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1556_ clknet_leaf_9_clk booth_b10_m30 VGND VGND VPWR VPWR pp_row40_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_141_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_71_8 s$165 s$167 s$169 VGND VGND VPWR VPWR c$742 s$743 sky130_fd_sc_hd__fa_2
X_0507_ clknet_leaf_172_clk booth_b24_m56 VGND VGND VPWR VPWR pp_row80_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_113_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1487_ clknet_leaf_34_clk booth_b12_m25 VGND VGND VPWR VPWR pp_row37_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_64_7 c$82 s$85 s$87 VGND VGND VPWR VPWR c$614 s$615 sky130_fd_sc_hd__fa_1
X_0438_ clknet_leaf_160_clk booth_b60_m17 VGND VGND VPWR VPWR pp_row77_24 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_57_6 pp_row57_26 pp_row57_27 pp_row57_28 VGND VGND VPWR VPWR c$486 s$487
+ sky130_fd_sc_hd__fa_1
Xclkbuf_leaf_187_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_187_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_28_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0369_ clknet_leaf_205_clk booth_b48_m27 VGND VGND VPWR VPWR pp_row75_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_39_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_746 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2108_ clknet_leaf_33_clk booth_b50_m8 VGND VGND VPWR VPWR pp_row58_25 sky130_fd_sc_hd__dfxtp_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_9_0 s$3435 c$3912 s$3915 VGND VGND VPWR VPWR c$4170 s$4171 sky130_fd_sc_hd__fa_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2039_ clknet_leaf_81_clk booth_b48_m8 VGND VGND VPWR VPWR pp_row56_24 sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_87_0 s$3747 c$4068 s$4071 VGND VGND VPWR VPWR c$4326 s$4327 sky130_fd_sc_hd__fa_2
XFILLER_182_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_111_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_111_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_184_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_90_0 net1901 pp_row90_1 pp_row90_2 VGND VGND VPWR VPWR c$1018 s$1019 sky130_fd_sc_hd__fa_1
XFILLER_2_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout840 net841 VGND VGND VPWR VPWR net840 sky130_fd_sc_hd__clkbuf_8
Xfanout851 net852 VGND VGND VPWR VPWR net851 sky130_fd_sc_hd__buf_4
Xfanout862 net865 VGND VGND VPWR VPWR net862 sky130_fd_sc_hd__clkbuf_8
XU$$4308 t$6606 net1258 VGND VGND VPWR VPWR booth_b62_m27 sky130_fd_sc_hd__xor2_1
Xfanout873 net874 VGND VGND VPWR VPWR net873 sky130_fd_sc_hd__buf_6
XFILLER_120_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4319 net1004 net425 net996 net707 VGND VGND VPWR VPWR t$6612 sky130_fd_sc_hd__a22o_1
Xfanout884 net885 VGND VGND VPWR VPWR net884 sky130_fd_sc_hd__buf_2
XFILLER_133_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout895 sel_1$4478 VGND VGND VPWR VPWR net895 sky130_fd_sc_hd__clkbuf_8
XTAP_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3607 t$6248 net1320 VGND VGND VPWR VPWR booth_b52_m19 sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_178_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_178_clk
+ sky130_fd_sc_hd__clkbuf_16
XU$$3618 net1085 net478 net1076 net751 VGND VGND VPWR VPWR t$6254 sky130_fd_sc_hd__a22o_1
XTAP_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3629 t$6259 net1323 VGND VGND VPWR VPWR booth_b52_m30 sky130_fd_sc_hd__xor2_1
XTAP_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_102_0 c$3800 c$3802 s$3805 VGND VGND VPWR VPWR c$4100 s$4101 sky130_fd_sc_hd__fa_1
XFILLER_18_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2906 t$5890 net1372 VGND VGND VPWR VPWR booth_b42_m11 sky130_fd_sc_hd__xor2_1
XFILLER_46_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_200 net1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2917 net1158 net520 net1148 net793 VGND VGND VPWR VPWR t$5896 sky130_fd_sc_hd__a22o_1
XTAP_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2928 t$5901 net1372 VGND VGND VPWR VPWR booth_b42_m22 sky130_fd_sc_hd__xor2_1
XANTENNA_211 net1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_222 net1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2939 net1060 net522 net1051 net795 VGND VGND VPWR VPWR t$5907 sky130_fd_sc_hd__a22o_1
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_233 net1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdadda_fa_3_22_3 pp_row22_11 pp_row22_12 pp_row22_13 VGND VGND VPWR VPWR c$2020 s$2021
+ sky130_fd_sc_hd__fa_1
XTAP_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_244 net1559 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_255 net1619 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_266 net1728 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_277 c$4210 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_288 sel_1$5248 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_299 net356 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_102_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_102_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_10_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1410_ clknet_leaf_58_clk booth_b28_m5 VGND VGND VPWR VPWR pp_row33_14 sky130_fd_sc_hd__dfxtp_1
X_2390_ clknet_leaf_96_clk booth_b38_m28 VGND VGND VPWR VPWR pp_row66_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_111_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1341_ clknet_leaf_0_clk booth_b14_m16 VGND VGND VPWR VPWR pp_row30_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_122_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_67_5 s$665 s$667 s$669 VGND VGND VPWR VPWR c$1540 s$1541 sky130_fd_sc_hd__fa_1
XFILLER_3_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1272_ clknet_leaf_10_clk booth_b18_m8 VGND VGND VPWR VPWR pp_row26_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0223_ clknet_leaf_196_clk booth_b20_m51 VGND VGND VPWR VPWR pp_row71_7 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_169_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_169_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_92_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$390 net1620 net530 net1612 net803 VGND VGND VPWR VPWR t$4604 sky130_fd_sc_hd__a22o_1
XFILLER_189_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0987_ clknet_leaf_115_clk booth_b50_m50 VGND VGND VPWR VPWR pp_row100_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_164_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1608_ clknet_leaf_240_clk booth_b14_m28 VGND VGND VPWR VPWR pp_row42_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_113_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_28__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_5_28__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_1539_ clknet_leaf_121_clk booth_b48_m57 VGND VGND VPWR VPWR pp_row105_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_86_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_62_4 pp_row62_29 pp_row62_30 pp_row62_31 VGND VGND VPWR VPWR c$572 s$573
+ sky130_fd_sc_hd__fa_1
Xdadda_fa_1_55_3 pp_row55_14 pp_row55_15 pp_row55_16 VGND VGND VPWR VPWR c$444 s$445
+ sky130_fd_sc_hd__fa_1
XFILLER_80_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_32_2 s$2097 s$2099 s$2101 VGND VGND VPWR VPWR c$2886 s$2887 sky130_fd_sc_hd__fa_1
Xdadda_fa_1_48_2 pp_row48_6 pp_row48_7 pp_row48_8 VGND VGND VPWR VPWR c$320 s$321
+ sky130_fd_sc_hd__fa_1
XFILLER_83_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_874 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_25_1 c$2034 c$2036 s$2039 VGND VGND VPWR VPWR c$2842 s$2843 sky130_fd_sc_hd__fa_1
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_18_0 pp_row18_8 pp_row18_9 pp_row18_10 VGND VGND VPWR VPWR c$2798 s$2799
+ sky130_fd_sc_hd__fa_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1602 net1603 VGND VGND VPWR VPWR net1602 sky130_fd_sc_hd__buf_4
XFILLER_137_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1613 net1614 VGND VGND VPWR VPWR net1613 sky130_fd_sc_hd__clkbuf_8
Xfanout1624 net1626 VGND VGND VPWR VPWR net1624 sky130_fd_sc_hd__buf_4
Xfanout1635 net1636 VGND VGND VPWR VPWR net1635 sky130_fd_sc_hd__buf_4
Xfanout1646 net1648 VGND VGND VPWR VPWR net1646 sky130_fd_sc_hd__clkbuf_8
XU$$4105 net1541 net454 net1533 net727 VGND VGND VPWR VPWR t$6502 sky130_fd_sc_hd__a22o_1
Xfanout1657 net110 VGND VGND VPWR VPWR net1657 sky130_fd_sc_hd__buf_4
Xfanout1668 net1669 VGND VGND VPWR VPWR net1668 sky130_fd_sc_hd__buf_6
XU$$4116 net1805 net434 net1229 net716 VGND VGND VPWR VPWR t$6509 sky130_fd_sc_hd__a22o_1
Xfanout670 net673 VGND VGND VPWR VPWR net670 sky130_fd_sc_hd__buf_4
XU$$4127 t$6514 net1269 VGND VGND VPWR VPWR booth_b60_m5 sky130_fd_sc_hd__xor2_1
Xfanout1679 net1681 VGND VGND VPWR VPWR net1679 sky130_fd_sc_hd__buf_4
Xfanout681 net683 VGND VGND VPWR VPWR net681 sky130_fd_sc_hd__buf_4
Xfanout692 sel_1 VGND VGND VPWR VPWR net692 sky130_fd_sc_hd__buf_6
XU$$4138 net1223 net434 net1215 net716 VGND VGND VPWR VPWR t$6520 sky130_fd_sc_hd__a22o_1
XU$$4149 t$6525 net1263 VGND VGND VPWR VPWR booth_b60_m16 sky130_fd_sc_hd__xor2_1
XU$$3404 net1624 net495 net1616 net768 VGND VGND VPWR VPWR t$6144 sky130_fd_sc_hd__a22o_1
XU$$3415 t$6149 net1345 VGND VGND VPWR VPWR booth_b48_m60 sky130_fd_sc_hd__xor2_1
XFILLER_18_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3426 net46 VGND VGND VPWR VPWR notblock$6155\[1\] sky130_fd_sc_hd__inv_1
XU$$3437 net1037 net488 net938 net761 VGND VGND VPWR VPWR t$6162 sky130_fd_sc_hd__a22o_1
XTAP_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2703 net1704 net545 net1696 net818 VGND VGND VPWR VPWR t$5786 sky130_fd_sc_hd__a22o_1
XFILLER_92_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3448 t$6167 net1332 VGND VGND VPWR VPWR booth_b50_m8 sky130_fd_sc_hd__xor2_1
XTAP_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2714 t$5791 net1401 VGND VGND VPWR VPWR booth_b38_m52 sky130_fd_sc_hd__xor2_1
XTAP_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3459 net1200 net488 net1181 net761 VGND VGND VPWR VPWR t$6173 sky130_fd_sc_hd__a22o_1
XFILLER_34_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2725 net1603 net547 net1593 net820 VGND VGND VPWR VPWR t$5797 sky130_fd_sc_hd__a22o_1
XFILLER_74_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2736 t$5802 net1401 VGND VGND VPWR VPWR booth_b38_m63 sky130_fd_sc_hd__xor2_1
XFILLER_61_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2747 t$5809 net1376 VGND VGND VPWR VPWR booth_b40_m0 sky130_fd_sc_hd__xor2_1
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2758 net1562 net536 net1521 net809 VGND VGND VPWR VPWR t$5815 sky130_fd_sc_hd__a22o_1
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_20_0 pp_row20_0 pp_row20_1 pp_row20_2 VGND VGND VPWR VPWR c$1998 s$1999
+ sky130_fd_sc_hd__fa_1
XTAP_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2769 t$5820 net1381 VGND VGND VPWR VPWR booth_b40_m11 sky130_fd_sc_hd__xor2_1
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0910_ clknet_leaf_133_clk booth_b64_m56 VGND VGND VPWR VPWR pp_row120_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_109_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1890_ clknet_leaf_39_clk booth_b12_m40 VGND VGND VPWR VPWR pp_row52_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_186_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0841_ clknet_leaf_102_clk booth_b34_m59 VGND VGND VPWR VPWR pp_row93_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_128_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0772_ clknet_leaf_144_clk booth_b32_m58 VGND VGND VPWR VPWR pp_row90_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_127_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2442_ clknet_leaf_98_clk booth_b62_m5 VGND VGND VPWR VPWR pp_row67_31 sky130_fd_sc_hd__dfxtp_1
XFILLER_5_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_72_3 c$742 s$745 s$747 VGND VGND VPWR VPWR c$1596 s$1597 sky130_fd_sc_hd__fa_1
X_2373_ clknet_leaf_84_clk booth_b6_m60 VGND VGND VPWR VPWR pp_row66_3 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_65_2 c$610 c$612 c$614 VGND VGND VPWR VPWR c$1510 s$1511 sky130_fd_sc_hd__fa_2
XFILLER_190_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1324_ clknet_leaf_250_clk booth_b16_m13 VGND VGND VPWR VPWR pp_row29_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_97_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$709 final_adder.p_new$716 final_adder.g_new$733 final_adder.g_new$717
+ VGND VGND VPWR VPWR final_adder.g_new$837 sky130_fd_sc_hd__a21o_1
Xdadda_fa_5_42_1 s$2943 s$2945 s$2947 VGND VGND VPWR VPWR c$3566 s$3567 sky130_fd_sc_hd__fa_2
XFILLER_112_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_58_1 c$478 c$480 c$482 VGND VGND VPWR VPWR c$1424 s$1425 sky130_fd_sc_hd__fa_1
XFILLER_56_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1255_ clknet_leaf_11_clk booth_b16_m9 VGND VGND VPWR VPWR pp_row25_8 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_35_0 c$2894 c$2896 c$2898 VGND VGND VPWR VPWR c$3536 s$3537 sky130_fd_sc_hd__fa_1
X_0206_ clknet_leaf_152_clk booth_b52_m18 VGND VGND VPWR VPWR pp_row70_24 sky130_fd_sc_hd__dfxtp_1
X_1186_ clknet_leaf_244_clk net169 VGND VGND VPWR VPWR pp_row20_12 sky130_fd_sc_hd__dfxtp_2
XU$$3960 net1591 net462 net1583 net735 VGND VGND VPWR VPWR t$6428 sky130_fd_sc_hd__a22o_1
XU$$3971 t$6433 net1293 VGND VGND VPWR VPWR booth_b56_m64 sky130_fd_sc_hd__xor2_1
XU$$3982 t$6440 net1282 VGND VGND VPWR VPWR booth_b58_m1 sky130_fd_sc_hd__xor2_1
XU$$3993 net1525 net455 net1517 net728 VGND VGND VPWR VPWR t$6446 sky130_fd_sc_hd__a22o_1
XFILLER_80_844 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_900 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput262 net262 VGND VGND VPWR VPWR o[104] sky130_fd_sc_hd__buf_2
XFILLER_160_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput273 net273 VGND VGND VPWR VPWR o[114] sky130_fd_sc_hd__buf_2
XFILLER_114_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput284 net284 VGND VGND VPWR VPWR o[124] sky130_fd_sc_hd__buf_2
XFILLER_160_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput295 net295 VGND VGND VPWR VPWR o[19] sky130_fd_sc_hd__buf_2
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3705_1797 VGND VGND VPWR VPWR U$$3705_1797/HI net1797 sky130_fd_sc_hd__conb_1
XFILLER_59_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_60_1 pp_row60_17 pp_row60_18 pp_row60_19 VGND VGND VPWR VPWR c$530 s$531
+ sky130_fd_sc_hd__fa_1
XFILLER_87_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_988 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_53_0 pp_row53_2 pp_row53_3 pp_row53_4 VGND VGND VPWR VPWR c$402 s$403
+ sky130_fd_sc_hd__fa_1
XFILLER_74_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1309 net987 net639 net978 net912 VGND VGND VPWR VPWR t$5074 sky130_fd_sc_hd__a22o_1
XFILLER_15_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_82_2 c$1708 s$1711 s$1713 VGND VGND VPWR VPWR c$2498 s$2499 sky130_fd_sc_hd__fa_1
XFILLER_125_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_75_1 c$1618 c$1620 c$1622 VGND VGND VPWR VPWR c$2440 s$2441 sky130_fd_sc_hd__fa_1
XFILLER_135_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_52_0 c$3600 c$3602 s$3605 VGND VGND VPWR VPWR c$4000 s$4001 sky130_fd_sc_hd__fa_2
Xfanout1410 net1411 VGND VGND VPWR VPWR net1410 sky130_fd_sc_hd__buf_6
Xdadda_fa_3_68_0 s$689 c$1530 c$1532 VGND VGND VPWR VPWR c$2382 s$2383 sky130_fd_sc_hd__fa_1
Xfanout1421 net1422 VGND VGND VPWR VPWR net1421 sky130_fd_sc_hd__buf_4
Xfanout1432 net1433 VGND VGND VPWR VPWR net1432 sky130_fd_sc_hd__buf_6
Xclkbuf_5_11__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_5_11__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xfanout1443 net1447 VGND VGND VPWR VPWR net1443 sky130_fd_sc_hd__buf_6
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1454 net1456 VGND VGND VPWR VPWR net1454 sky130_fd_sc_hd__buf_6
Xfanout1465 net20 VGND VGND VPWR VPWR net1465 sky130_fd_sc_hd__buf_8
Xfanout1476 net1477 VGND VGND VPWR VPWR net1476 sky130_fd_sc_hd__clkbuf_4
XFILLER_65_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1487 net1489 VGND VGND VPWR VPWR net1487 sky130_fd_sc_hd__buf_6
XU$$3201 net1113 net506 net1104 net779 VGND VGND VPWR VPWR t$6041 sky130_fd_sc_hd__a22o_1
Xfanout1498 net1502 VGND VGND VPWR VPWR net1498 sky130_fd_sc_hd__buf_6
XU$$3212 t$6046 net1348 VGND VGND VPWR VPWR booth_b46_m27 sky130_fd_sc_hd__xor2_1
XFILLER_4_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3223 net1002 net504 net994 net777 VGND VGND VPWR VPWR t$6052 sky130_fd_sc_hd__a22o_1
XFILLER_93_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_111_2 s$2727 s$2729 s$2731 VGND VGND VPWR VPWR c$3360 s$3361 sky130_fd_sc_hd__fa_1
XFILLER_171_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1040_ clknet_leaf_57_clk booth_b0_m6 VGND VGND VPWR VPWR pp_row6_0 sky130_fd_sc_hd__dfxtp_1
XU$$3234 t$6057 net1351 VGND VGND VPWR VPWR booth_b46_m38 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$16 c$4182 s$4185 VGND VGND VPWR VPWR final_adder.$signal$34 final_adder.$signal$1106
+ sky130_fd_sc_hd__ha_1
XU$$2500 net1198 net554 net1180 net827 VGND VGND VPWR VPWR t$5683 sky130_fd_sc_hd__a22o_1
Xdadda_fa_1_94_0_1903 VGND VGND VPWR VPWR net1903 dadda_fa_1_94_0_1903/LO sky130_fd_sc_hd__conb_1
XU$$3245 net1735 net508 net1727 net781 VGND VGND VPWR VPWR t$6063 sky130_fd_sc_hd__a22o_1
XFILLER_185_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3256 t$6068 net1354 VGND VGND VPWR VPWR booth_b46_m49 sky130_fd_sc_hd__xor2_1
XU$$2511 t$5688 net1406 VGND VGND VPWR VPWR booth_b36_m19 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$27 c$4204 s$4207 VGND VGND VPWR VPWR final_adder.$signal$56 final_adder.$signal$1117
+ sky130_fd_sc_hd__ha_2
XU$$3267 net1626 net508 net1618 net781 VGND VGND VPWR VPWR t$6074 sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_104_1 c$2666 c$2668 s$2671 VGND VGND VPWR VPWR c$3316 s$3317 sky130_fd_sc_hd__fa_1
XU$$2522 net1082 net553 net1079 net826 VGND VGND VPWR VPWR t$5694 sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$38 c$4226 s$4229 VGND VGND VPWR VPWR final_adder.$signal$78 final_adder.$signal$1128
+ sky130_fd_sc_hd__ha_1
XU$$2533 t$5699 net1407 VGND VGND VPWR VPWR booth_b36_m30 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$49 c$4248 s$4251 VGND VGND VPWR VPWR final_adder.$signal$100 final_adder.$signal$101
+ sky130_fd_sc_hd__ha_1
XU$$3278 t$6079 net1356 VGND VGND VPWR VPWR booth_b46_m60 sky130_fd_sc_hd__xor2_1
XU$$2544 net976 net556 net967 net829 VGND VGND VPWR VPWR t$5705 sky130_fd_sc_hd__a22o_1
XU$$3289 net43 VGND VGND VPWR VPWR notblock$6085\[1\] sky130_fd_sc_hd__inv_1
XFILLER_185_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2555 t$5710 net1409 VGND VGND VPWR VPWR booth_b36_m41 sky130_fd_sc_hd__xor2_1
XU$$1810 t$5330 net1460 VGND VGND VPWR VPWR booth_b26_m11 sky130_fd_sc_hd__xor2_1
XFILLER_34_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2566 net1704 net555 net1696 net828 VGND VGND VPWR VPWR t$5716 sky130_fd_sc_hd__a22o_1
XU$$1821 net1156 net593 net1147 net866 VGND VGND VPWR VPWR t$5336 sky130_fd_sc_hd__a22o_1
XU$$1832 t$5341 net1459 VGND VGND VPWR VPWR booth_b26_m22 sky130_fd_sc_hd__xor2_1
XFILLER_62_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2577 t$5721 net1411 VGND VGND VPWR VPWR booth_b36_m52 sky130_fd_sc_hd__xor2_1
XU$$2588 net1599 net557 net1593 net830 VGND VGND VPWR VPWR t$5727 sky130_fd_sc_hd__a22o_1
XU$$1843 net1057 net597 net1049 net870 VGND VGND VPWR VPWR t$5347 sky130_fd_sc_hd__a22o_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1854 t$5352 net1462 VGND VGND VPWR VPWR booth_b26_m33 sky130_fd_sc_hd__xor2_1
XU$$2599 t$5732 net1411 VGND VGND VPWR VPWR booth_b36_m63 sky130_fd_sc_hd__xor2_1
XU$$1865 net955 net601 net944 net874 VGND VGND VPWR VPWR t$5358 sky130_fd_sc_hd__a22o_1
XU$$1876 t$5363 net1465 VGND VGND VPWR VPWR booth_b26_m44 sky130_fd_sc_hd__xor2_1
X_1942_ clknet_leaf_72_clk booth_b48_m5 VGND VGND VPWR VPWR pp_row53_24 sky130_fd_sc_hd__dfxtp_1
XU$$1887 net1679 net598 net1654 net871 VGND VGND VPWR VPWR t$5369 sky130_fd_sc_hd__a22o_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1898 t$5374 net1464 VGND VGND VPWR VPWR booth_b26_m55 sky130_fd_sc_hd__xor2_1
Xdadda_fa_7_125_0 s$3897 c$4144 s$4147 VGND VGND VPWR VPWR c$4402 s$4403 sky130_fd_sc_hd__fa_2
XFILLER_159_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1873_ clknet_leaf_71_clk booth_b34_m17 VGND VGND VPWR VPWR pp_row51_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_174_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0824_ clknet_leaf_109_clk booth_b44_m48 VGND VGND VPWR VPWR pp_row92_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_960 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0755_ clknet_leaf_132_clk booth_b62_m56 VGND VGND VPWR VPWR pp_row118_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_171_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0686_ clknet_leaf_168_clk booth_b54_m32 VGND VGND VPWR VPWR pp_row86_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_103_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2425_ clknet_leaf_124_clk booth_b64_m47 VGND VGND VPWR VPWR pp_row111_9 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_70_0 s$163 c$690 c$692 VGND VGND VPWR VPWR c$1566 s$1567 sky130_fd_sc_hd__fa_1
XFILLER_9_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2356_ clknet_leaf_98_clk booth_b42_m23 VGND VGND VPWR VPWR pp_row65_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_9_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$517 final_adder.p_new$520 final_adder.g_new$529 final_adder.g_new$521
+ VGND VGND VPWR VPWR final_adder.g_new$645 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$528 final_adder.p_new$540 final_adder.p_new$532 VGND VGND VPWR VPWR
+ final_adder.p_new$656 sky130_fd_sc_hd__and2_1
X_1307_ clknet_leaf_1_clk booth_b18_m10 VGND VGND VPWR VPWR pp_row28_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_29_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$539 final_adder.p_new$542 final_adder.g_new$551 final_adder.g_new$543
+ VGND VGND VPWR VPWR final_adder.g_new$667 sky130_fd_sc_hd__a21o_1
X_2287_ clknet_leaf_210_clk booth_b48_m15 VGND VGND VPWR VPWR pp_row63_24 sky130_fd_sc_hd__dfxtp_1
XFILLER_56_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1238_ clknet_leaf_109_clk booth_b50_m53 VGND VGND VPWR VPWR pp_row103_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_65_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4480 net1727 sel_0$6647 net1719 net696 VGND VGND VPWR VPWR t$6694 sky130_fd_sc_hd__a22o_1
XU$$4491 t$6699 net1866 VGND VGND VPWR VPWR booth_b64_m50 sky130_fd_sc_hd__xor2_1
X_1169_ clknet_leaf_47_clk booth_b18_m1 VGND VGND VPWR VPWR pp_row19_9 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_91_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_91_clk sky130_fd_sc_hd__clkbuf_16
XU$$3790 t$6341 net1307 VGND VGND VPWR VPWR booth_b54_m42 sky130_fd_sc_hd__xor2_1
XFILLER_52_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_92_1 c$2570 c$2572 s$2575 VGND VGND VPWR VPWR c$3244 s$3245 sky130_fd_sc_hd__fa_1
XU$$4393_1817 VGND VGND VPWR VPWR U$$4393_1817/HI net1817 sky130_fd_sc_hd__conb_1
XFILLER_10_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_85_0 s$1757 c$2510 c$2512 VGND VGND VPWR VPWR c$3200 s$3201 sky130_fd_sc_hd__fa_1
Xdadda_fa_3_106_3 c$1962 c$1964 s$1967 VGND VGND VPWR VPWR c$2692 s$2693 sky130_fd_sc_hd__fa_1
XFILLER_192_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$901 t$4865 net1311 VGND VGND VPWR VPWR booth_b12_m36 sky130_fd_sc_hd__xor2_1
XU$$912 net1752 net398 net1744 net664 VGND VGND VPWR VPWR t$4871 sky130_fd_sc_hd__a22o_1
XU$$923 t$4876 net1317 VGND VGND VPWR VPWR booth_b12_m47 sky130_fd_sc_hd__xor2_1
XU$$934 net1641 net399 net1633 net665 VGND VGND VPWR VPWR t$4882 sky130_fd_sc_hd__a22o_1
XFILLER_28_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$945 t$4887 net1318 VGND VGND VPWR VPWR booth_b12_m58 sky130_fd_sc_hd__xor2_1
XU$$956 net1530 net395 net1888 net661 VGND VGND VPWR VPWR t$4893 sky130_fd_sc_hd__a22o_1
XFILLER_141_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1106 net1123 net646 net1032 net919 VGND VGND VPWR VPWR t$4971 sky130_fd_sc_hd__a22o_1
XU$$967 net1230 net387 net1123 net653 VGND VGND VPWR VPWR t$4900 sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_82_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_82_clk sky130_fd_sc_hd__clkbuf_16
XU$$1117 t$4976 net1009 VGND VGND VPWR VPWR booth_b16_m7 sky130_fd_sc_hd__xor2_1
XU$$978 t$4905 net1187 VGND VGND VPWR VPWR booth_b14_m6 sky130_fd_sc_hd__xor2_1
XU$$1128 net1201 net643 net1192 net916 VGND VGND VPWR VPWR t$4982 sky130_fd_sc_hd__a22o_1
XU$$989 net1210 net385 net1201 net651 VGND VGND VPWR VPWR t$4911 sky130_fd_sc_hd__a22o_1
XU$$1139 t$4987 net1010 VGND VGND VPWR VPWR booth_b16_m18 sky130_fd_sc_hd__xor2_1
XFILLER_70_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1046 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0540_ clknet_leaf_165_clk booth_b32_m49 VGND VGND VPWR VPWR pp_row81_8 sky130_fd_sc_hd__dfxtp_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0471_ clknet_leaf_197_clk net232 VGND VGND VPWR VPWR pp_row78_27 sky130_fd_sc_hd__dfxtp_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ clknet_leaf_212_clk booth_b42_m19 VGND VGND VPWR VPWR pp_row61_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_79_752 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1240 net1243 VGND VGND VPWR VPWR net1240 sky130_fd_sc_hd__buf_2
XFILLER_26_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1251 net1252 VGND VGND VPWR VPWR net1251 sky130_fd_sc_hd__buf_6
X_2141_ clknet_leaf_219_clk booth_b46_m13 VGND VGND VPWR VPWR pp_row59_23 sky130_fd_sc_hd__dfxtp_1
Xfanout1262 net60 VGND VGND VPWR VPWR net1262 sky130_fd_sc_hd__buf_6
Xfanout1273 net1274 VGND VGND VPWR VPWR net1273 sky130_fd_sc_hd__buf_6
XFILLER_94_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_906 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1284 net1285 VGND VGND VPWR VPWR net1284 sky130_fd_sc_hd__clkbuf_4
XFILLER_66_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1295 net53 VGND VGND VPWR VPWR net1295 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_42_4 c$240 c$242 s$245 VGND VGND VPWR VPWR c$1238 s$1239 sky130_fd_sc_hd__fa_1
XU$$3020 net1787 net510 net1229 net783 VGND VGND VPWR VPWR t$5949 sky130_fd_sc_hd__a22o_1
X_2072_ clknet_leaf_143_clk notsign$6014 VGND VGND VPWR VPWR pp_row109_0 sky130_fd_sc_hd__dfxtp_1
XU$$3031 t$5954 net1357 VGND VGND VPWR VPWR booth_b44_m5 sky130_fd_sc_hd__xor2_1
XU$$3042 net1226 net514 net1217 net787 VGND VGND VPWR VPWR t$5960 sky130_fd_sc_hd__a22o_1
XFILLER_47_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1023_ clknet_leaf_60_clk booth_b2_m0 VGND VGND VPWR VPWR pp_row2_1 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_35_3 pp_row35_11 pp_row35_12 pp_row35_13 VGND VGND VPWR VPWR c$1152 s$1153
+ sky130_fd_sc_hd__fa_1
XU$$3053 t$5965 net1357 VGND VGND VPWR VPWR booth_b44_m16 sky130_fd_sc_hd__xor2_1
XU$$3064 net1113 net517 net1104 net790 VGND VGND VPWR VPWR t$5971 sky130_fd_sc_hd__a22o_1
XFILLER_81_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_73_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_73_clk sky130_fd_sc_hd__clkbuf_16
XU$$2330 net28 VGND VGND VPWR VPWR notblock$5595\[1\] sky130_fd_sc_hd__inv_1
XFILLER_62_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3075 t$5976 net1358 VGND VGND VPWR VPWR booth_b44_m27 sky130_fd_sc_hd__xor2_1
XU$$3086 net1002 net510 net994 net783 VGND VGND VPWR VPWR t$5982 sky130_fd_sc_hd__a22o_1
XU$$2341 net1036 net563 net936 net836 VGND VGND VPWR VPWR t$5602 sky130_fd_sc_hd__a22o_1
XU$$2352 t$5607 net1420 VGND VGND VPWR VPWR booth_b34_m8 sky130_fd_sc_hd__xor2_1
XU$$3097 t$5987 net1359 VGND VGND VPWR VPWR booth_b44_m38 sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_28_2 pp_row28_6 pp_row28_7 pp_row28_8 VGND VGND VPWR VPWR c$1078 s$1079
+ sky130_fd_sc_hd__fa_1
XU$$2363 net1193 net560 net1174 net833 VGND VGND VPWR VPWR t$5613 sky130_fd_sc_hd__a22o_1
XFILLER_179_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2374 t$5618 net1423 VGND VGND VPWR VPWR booth_b34_m19 sky130_fd_sc_hd__xor2_1
XFILLER_34_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1640 t$5242 net1481 VGND VGND VPWR VPWR booth_b22_m63 sky130_fd_sc_hd__xor2_1
XU$$2385 net1082 net561 net1073 net834 VGND VGND VPWR VPWR t$5624 sky130_fd_sc_hd__a22o_1
XU$$1651 t$5249 net1466 VGND VGND VPWR VPWR booth_b24_m0 sky130_fd_sc_hd__xor2_1
XU$$2396 t$5629 net1422 VGND VGND VPWR VPWR booth_b34_m30 sky130_fd_sc_hd__xor2_1
XU$$1662 net1560 net602 net1519 net875 VGND VGND VPWR VPWR t$5255 sky130_fd_sc_hd__a22o_1
XU$$1673 t$5260 net1469 VGND VGND VPWR VPWR booth_b24_m11 sky130_fd_sc_hd__xor2_1
XFILLER_50_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1684 net1155 net602 net1146 net875 VGND VGND VPWR VPWR t$5266 sky130_fd_sc_hd__a22o_1
XU$$1695 t$5271 net1467 VGND VGND VPWR VPWR booth_b24_m22 sky130_fd_sc_hd__xor2_1
XFILLER_188_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1925_ clknet_leaf_65_clk booth_b18_m35 VGND VGND VPWR VPWR pp_row53_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1856_ clknet_leaf_67_clk booth_b4_m47 VGND VGND VPWR VPWR pp_row51_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0807_ clknet_leaf_94_clk booth_b54_m37 VGND VGND VPWR VPWR pp_row91_14 sky130_fd_sc_hd__dfxtp_1
X_1787_ clknet_leaf_220_clk booth_b42_m6 VGND VGND VPWR VPWR pp_row48_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_760 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0738_ clknet_leaf_163_clk booth_b56_m32 VGND VGND VPWR VPWR pp_row88_17 sky130_fd_sc_hd__dfxtp_1
XFILLER_1_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0669_ clknet_leaf_180_clk booth_b22_m64 VGND VGND VPWR VPWR pp_row86_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_103_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2408_ clknet_leaf_84_clk notsign VGND VGND VPWR VPWR pp_row67_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_162_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$303 final_adder.p_new$302 final_adder.g_new$305 final_adder.g_new$303
+ VGND VGND VPWR VPWR final_adder.g_new$431 sky130_fd_sc_hd__a21o_1
XTAP_4319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2339_ clknet_leaf_89_clk booth_b10_m55 VGND VGND VPWR VPWR pp_row65_5 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$314 final_adder.p_new$316 final_adder.p_new$314 VGND VGND VPWR VPWR
+ final_adder.p_new$442 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$325 final_adder.p_new$324 final_adder.g_new$327 final_adder.g_new$325
+ VGND VGND VPWR VPWR final_adder.g_new$453 sky130_fd_sc_hd__a21o_1
XTAP_3607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$336 final_adder.p_new$338 final_adder.p_new$336 VGND VGND VPWR VPWR
+ final_adder.p_new$464 sky130_fd_sc_hd__and2_1
XTAP_3618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$347 final_adder.p_new$346 final_adder.g_new$349 final_adder.g_new$347
+ VGND VGND VPWR VPWR final_adder.g_new$475 sky130_fd_sc_hd__a21o_1
XTAP_3629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$358 final_adder.p_new$360 final_adder.p_new$358 VGND VGND VPWR VPWR
+ final_adder.p_new$486 sky130_fd_sc_hd__and2_1
XU$$208 t$4511 net1389 VGND VGND VPWR VPWR booth_b2_m32 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$369 final_adder.p_new$368 final_adder.g_new$371 final_adder.g_new$369
+ VGND VGND VPWR VPWR final_adder.g_new$497 sky130_fd_sc_hd__a21o_1
XFILLER_26_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$219 net956 net619 net948 net892 VGND VGND VPWR VPWR t$4517 sky130_fd_sc_hd__a22o_1
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_64_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_64_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_37_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_111_1 pp_row111_3 pp_row111_4 pp_row111_5 VGND VGND VPWR VPWR c$2728 s$2729
+ sky130_fd_sc_hd__fa_1
XFILLER_14_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_579 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_104_0 pp_row104_8 pp_row104_9 pp_row104_10 VGND VGND VPWR VPWR c$2670
+ s$2671 sky130_fd_sc_hd__fa_1
XFILLER_122_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_52_3 s$1355 s$1357 s$1359 VGND VGND VPWR VPWR c$2260 s$2261 sky130_fd_sc_hd__fa_1
XFILLER_0_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_0_68_3 pp_row68_9 pp_row68_10 pp_row68_11 VGND VGND VPWR VPWR c$138 s$139
+ sky130_fd_sc_hd__fa_1
XFILLER_49_969 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_45_2 c$1264 s$1267 s$1269 VGND VGND VPWR VPWR c$2202 s$2203 sky130_fd_sc_hd__fa_1
XFILLER_29_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$881 final_adder.p_new$912 final_adder.g_new$865 final_adder.g_new$913
+ VGND VGND VPWR VPWR final_adder.g_new$1009 sky130_fd_sc_hd__a21o_1
XFILLER_21_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$720 t$4773 net1415 VGND VGND VPWR VPWR booth_b10_m14 sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_38_1 c$1174 c$1176 c$1178 VGND VGND VPWR VPWR c$2144 s$2145 sky130_fd_sc_hd__fa_1
XU$$731 net1130 net401 net1114 net667 VGND VGND VPWR VPWR t$4779 sky130_fd_sc_hd__a22o_1
XU$$742 t$4784 net1414 VGND VGND VPWR VPWR booth_b10_m25 sky130_fd_sc_hd__xor2_1
Xdadda_fa_6_15_0 c$3452 c$3454 s$3457 VGND VGND VPWR VPWR c$3926 s$3927 sky130_fd_sc_hd__fa_2
Xclkbuf_leaf_55_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_55_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_28_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$753 net1023 net401 net1015 net667 VGND VGND VPWR VPWR t$4790 sky130_fd_sc_hd__a22o_1
XU$$764 t$4795 net1413 VGND VGND VPWR VPWR booth_b10_m36 sky130_fd_sc_hd__xor2_1
XU$$775 net1749 net405 net1741 net671 VGND VGND VPWR VPWR t$4801 sky130_fd_sc_hd__a22o_1
XU$$786 t$4806 net1416 VGND VGND VPWR VPWR booth_b10_m47 sky130_fd_sc_hd__xor2_1
XFILLER_32_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$797 net1638 net403 net1629 net669 VGND VGND VPWR VPWR t$4812 sky130_fd_sc_hd__a22o_1
XFILLER_43_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_3_110_3 pp_row110_9 pp_row110_10 VGND VGND VPWR VPWR c$2724 s$2725 sky130_fd_sc_hd__ha_1
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1710_ clknet_leaf_236_clk booth_b6_m40 VGND VGND VPWR VPWR pp_row46_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_145_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1641_ clknet_leaf_240_clk booth_b24_m19 VGND VGND VPWR VPWR pp_row43_12 sky130_fd_sc_hd__dfxtp_1
XANTENNA_3 c$4184 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_790 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_97_5 pp_row97_15 pp_row97_16 pp_row97_17 VGND VGND VPWR VPWR c$1900 s$1901
+ sky130_fd_sc_hd__fa_2
XFILLER_6_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1572_ clknet_leaf_108_clk booth_b54_m51 VGND VGND VPWR VPWR pp_row105_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_99_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_5_9__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_5_9__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_4_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0523_ clknet_leaf_163_clk booth_b52_m28 VGND VGND VPWR VPWR pp_row80_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_112_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0454_ clknet_leaf_158_clk booth_b36_m42 VGND VGND VPWR VPWR pp_row78_12 sky130_fd_sc_hd__dfxtp_1
XFILLER_100_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0385_ clknet_leaf_195_clk booth_b22_m54 VGND VGND VPWR VPWR pp_row76_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_66_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1070 net83 VGND VGND VPWR VPWR net1070 sky130_fd_sc_hd__buf_6
XFILLER_6_1069 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1081 net1082 VGND VGND VPWR VPWR net1081 sky130_fd_sc_hd__buf_4
Xfanout1092 net1093 VGND VGND VPWR VPWR net1092 sky130_fd_sc_hd__clkbuf_8
X_2124_ clknet_leaf_218_clk booth_b16_m43 VGND VGND VPWR VPWR pp_row59_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_67_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_40_1 pp_row40_14 pp_row40_15 pp_row40_16 VGND VGND VPWR VPWR c$1208 s$1209
+ sky130_fd_sc_hd__fa_1
XFILLER_187_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2055_ clknet_leaf_38_clk booth_b16_m41 VGND VGND VPWR VPWR pp_row57_8 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_46_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_46_clk sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_2_33_0 pp_row33_0 pp_row33_1 pp_row33_2 VGND VGND VPWR VPWR c$1122 s$1123
+ sky130_fd_sc_hd__fa_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1006_ clknet_leaf_117_clk booth_b52_m49 VGND VGND VPWR VPWR pp_row101_8 sky130_fd_sc_hd__dfxtp_1
XU$$2160 t$5508 net1445 VGND VGND VPWR VPWR booth_b30_m49 sky130_fd_sc_hd__xor2_1
XFILLER_35_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2171 net1622 net578 net1613 net851 VGND VGND VPWR VPWR t$5514 sky130_fd_sc_hd__a22o_1
XU$$2182 t$5519 net1446 VGND VGND VPWR VPWR booth_b30_m60 sky130_fd_sc_hd__xor2_1
XFILLER_168_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2193 net26 VGND VGND VPWR VPWR notblock$5525\[1\] sky130_fd_sc_hd__inv_1
XFILLER_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1470 net1710 net634 net1702 net907 VGND VGND VPWR VPWR t$5156 sky130_fd_sc_hd__a22o_1
XU$$1481 t$5161 net1492 VGND VGND VPWR VPWR booth_b20_m52 sky130_fd_sc_hd__xor2_1
XU$$1492 net1596 net632 net1587 net905 VGND VGND VPWR VPWR t$5167 sky130_fd_sc_hd__a22o_1
XFILLER_50_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1908_ clknet_leaf_70_clk booth_b44_m8 VGND VGND VPWR VPWR pp_row52_22 sky130_fd_sc_hd__dfxtp_1
Xdadda_ha_1_86_5 pp_row86_15 pp_row86_16 VGND VGND VPWR VPWR c$988 s$989 sky130_fd_sc_hd__ha_1
XFILLER_148_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1839_ clknet_leaf_181_clk net155 VGND VGND VPWR VPWR pp_row123_4 sky130_fd_sc_hd__dfxtp_2
XFILLER_135_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_85_3 pp_row85_9 pp_row85_10 pp_row85_11 VGND VGND VPWR VPWR c$972 s$973
+ sky130_fd_sc_hd__fa_1
XFILLER_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_62_2 s$2337 s$2339 s$2341 VGND VGND VPWR VPWR c$3066 s$3067 sky130_fd_sc_hd__fa_1
XFILLER_132_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_1020 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_78_2 pp_row78_8 pp_row78_9 pp_row78_10 VGND VGND VPWR VPWR c$856 s$857
+ sky130_fd_sc_hd__fa_1
Xdadda_fa_4_55_1 c$2274 c$2276 s$2279 VGND VGND VPWR VPWR c$3022 s$3023 sky130_fd_sc_hd__fa_1
XFILLER_83_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$100 c$4350 s$4353 VGND VGND VPWR VPWR final_adder.$signal$202 final_adder.$signal$1190
+ sky130_fd_sc_hd__ha_1
XTAP_4116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_32_0 s$3527 c$3958 s$3961 VGND VGND VPWR VPWR c$4216 s$4217 sky130_fd_sc_hd__fa_2
XFILLER_97_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$111 c$4372 s$4375 VGND VGND VPWR VPWR final_adder.$signal$224 final_adder.$signal$1201
+ sky130_fd_sc_hd__ha_1
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$122 c$4394 s$4397 VGND VGND VPWR VPWR final_adder.$signal$246 final_adder.$signal$1212
+ sky130_fd_sc_hd__ha_2
XTAP_4138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_48_0 s$1313 c$2214 c$2216 VGND VGND VPWR VPWR c$2978 s$2979 sky130_fd_sc_hd__fa_1
XTAP_4149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$133 final_adder.$signal$1213 final_adder.$signal$246 final_adder.$signal$248
+ VGND VGND VPWR VPWR final_adder.g_new$261 sky130_fd_sc_hd__a21o_1
XFILLER_131_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$144 final_adder.$signal$1200 final_adder.$signal$1201 VGND VGND VPWR
+ VPWR final_adder.p_new$272 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$155 final_adder.$signal$1191 final_adder.$signal$202 final_adder.$signal$204
+ VGND VGND VPWR VPWR final_adder.g_new$283 sky130_fd_sc_hd__a21o_1
XTAP_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$166 final_adder.$signal$1178 final_adder.$signal$1179 VGND VGND VPWR
+ VPWR final_adder.p_new$294 sky130_fd_sc_hd__and2_1
XTAP_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$177 final_adder.$signal$1169 final_adder.$signal$158 final_adder.$signal$160
+ VGND VGND VPWR VPWR final_adder.g_new$305 sky130_fd_sc_hd__a21o_1
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_404 net1683 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$188 final_adder.$signal$1156 final_adder.$signal$1157 VGND VGND VPWR
+ VPWR final_adder.p_new$316 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$199 final_adder.$signal$1147 final_adder.$signal$114 final_adder.$signal$116
+ VGND VGND VPWR VPWR final_adder.g_new$327 sky130_fd_sc_hd__a21o_1
XFILLER_38_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_415 net125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_426 net658 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_37_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_16
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_437 net865 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_448 net1502 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_459 net1640 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_963 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_760 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_0_73_1 pp_row73_3 pp_row73_4 pp_row73_5 VGND VGND VPWR VPWR c$182 s$183
+ sky130_fd_sc_hd__fa_1
XFILLER_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput140 c[10] VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_3_50_0 s$365 c$1314 c$1316 VGND VGND VPWR VPWR c$2238 s$2239 sky130_fd_sc_hd__fa_1
Xdadda_fa_0_66_0 pp_row0_1 pp_row66_1 pp_row66_2 VGND VGND VPWR VPWR c$108 s$109 sky130_fd_sc_hd__fa_1
Xinput151 c[11] VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_1
Xinput162 c[14] VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_1
Xinput173 c[24] VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_1
X_0170_ clknet_leaf_97_clk booth_b48_m21 VGND VGND VPWR VPWR pp_row69_22 sky130_fd_sc_hd__dfxtp_1
Xinput184 c[34] VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_1
Xinput195 c[44] VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_28_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_16
XTAP_3971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$550 net1237 VGND VGND VPWR VPWR notblock$4685\[2\] sky130_fd_sc_hd__inv_1
XTAP_3993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$561 t$4692 net1239 VGND VGND VPWR VPWR booth_b8_m3 sky130_fd_sc_hd__xor2_1
XFILLER_32_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$572 net1505 net410 net1496 net676 VGND VGND VPWR VPWR t$4698 sky130_fd_sc_hd__a22o_1
XU$$583 t$4703 net1239 VGND VGND VPWR VPWR booth_b8_m14 sky130_fd_sc_hd__xor2_1
XU$$594 net1130 net409 net1114 net675 VGND VGND VPWR VPWR t$4709 sky130_fd_sc_hd__a22o_1
XFILLER_16_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_95_2 pp_row95_9 pp_row95_10 pp_row95_11 VGND VGND VPWR VPWR c$1870 s$1871
+ sky130_fd_sc_hd__fa_1
XFILLER_172_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_579 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1624_ clknet_leaf_239_clk booth_b42_m0 VGND VGND VPWR VPWR pp_row42_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_114_900 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1031 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_72_1 s$3123 s$3125 s$3127 VGND VGND VPWR VPWR c$3686 s$3687 sky130_fd_sc_hd__fa_2
Xdadda_fa_2_88_1 pp_row88_17 pp_row88_18 pp_row88_19 VGND VGND VPWR VPWR c$1784 s$1785
+ sky130_fd_sc_hd__fa_1
XFILLER_28_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1555_ clknet_leaf_7_clk booth_b8_m32 VGND VGND VPWR VPWR pp_row40_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_65_0 c$3074 c$3076 c$3078 VGND VGND VPWR VPWR c$3656 s$3657 sky130_fd_sc_hd__fa_1
XFILLER_113_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3842_1799 VGND VGND VPWR VPWR U$$3842_1799/HI net1799 sky130_fd_sc_hd__conb_1
X_0506_ clknet_leaf_172_clk booth_b22_m58 VGND VGND VPWR VPWR pp_row80_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_87_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1486_ clknet_leaf_43_clk booth_b10_m27 VGND VGND VPWR VPWR pp_row37_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_141_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0437_ clknet_leaf_153_clk booth_b58_m19 VGND VGND VPWR VPWR pp_row77_23 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_64_8 s$89 s$91 s$93 VGND VGND VPWR VPWR c$616 s$617 sky130_fd_sc_hd__fa_1
XFILLER_189_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_57_7 pp_row57_29 c$12 c$14 VGND VGND VPWR VPWR c$488 s$489 sky130_fd_sc_hd__fa_1
X_0368_ clknet_leaf_205_clk booth_b46_m29 VGND VGND VPWR VPWR pp_row75_18 sky130_fd_sc_hd__dfxtp_1
XFILLER_55_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2107_ clknet_leaf_33_clk booth_b48_m10 VGND VGND VPWR VPWR pp_row58_24 sky130_fd_sc_hd__dfxtp_1
XFILLER_27_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_19_clk clknet_5_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_16
X_0299_ clknet_leaf_226_clk booth_b38_m35 VGND VGND VPWR VPWR pp_row73_15 sky130_fd_sc_hd__dfxtp_1
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2038_ clknet_leaf_135_clk booth_b62_m46 VGND VGND VPWR VPWR pp_row108_10 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_6_4_0 pp_row4_2 pp_row4_3 pp_row4_4 VGND VGND VPWR VPWR c$3904 s$3905 sky130_fd_sc_hd__fa_1
XFILLER_39_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_90_1 pp_row90_3 pp_row90_4 pp_row90_5 VGND VGND VPWR VPWR c$1020 s$1021
+ sky130_fd_sc_hd__fa_1
XFILLER_117_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_83_0 pp_row83_0 pp_row83_1 pp_row83_2 VGND VGND VPWR VPWR c$938 s$939
+ sky130_fd_sc_hd__fa_1
XFILLER_116_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout830 net831 VGND VGND VPWR VPWR net830 sky130_fd_sc_hd__buf_4
Xfanout841 sel_1$5598 VGND VGND VPWR VPWR net841 sky130_fd_sc_hd__buf_8
Xfanout852 net856 VGND VGND VPWR VPWR net852 sky130_fd_sc_hd__buf_6
Xfanout863 net865 VGND VGND VPWR VPWR net863 sky130_fd_sc_hd__clkbuf_4
XFILLER_58_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4309 net1062 net422 net1053 net704 VGND VGND VPWR VPWR t$6607 sky130_fd_sc_hd__a22o_1
Xfanout874 sel_1$5318 VGND VGND VPWR VPWR net874 sky130_fd_sc_hd__buf_6
Xfanout885 sel_1$5178 VGND VGND VPWR VPWR net885 sky130_fd_sc_hd__buf_6
Xfanout896 net898 VGND VGND VPWR VPWR net896 sky130_fd_sc_hd__clkbuf_4
XFILLER_133_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3608 net1136 net476 net1120 net749 VGND VGND VPWR VPWR t$6249 sky130_fd_sc_hd__a22o_1
XFILLER_133_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3619 t$6254 net1322 VGND VGND VPWR VPWR booth_b52_m25 sky130_fd_sc_hd__xor2_1
XTAP_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2907 net1217 net523 net1207 net796 VGND VGND VPWR VPWR t$5891 sky130_fd_sc_hd__a22o_1
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2918 t$5896 net1368 VGND VGND VPWR VPWR booth_b42_m17 sky130_fd_sc_hd__xor2_1
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_201 net1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2929 net1104 net523 net1092 net796 VGND VGND VPWR VPWR t$5902 sky130_fd_sc_hd__a22o_1
XANTENNA_212 net1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_223 net1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_234 net1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_245 net1559 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_256 net1619 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_267 net1728 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_278 c$4212 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_289 sel_1$6228 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_997 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_82_0 c$3720 c$3722 s$3725 VGND VGND VPWR VPWR c$4060 s$4061 sky130_fd_sc_hd__fa_1
Xdadda_fa_3_98_0 pp_row98_17 c$1890 c$1892 VGND VGND VPWR VPWR c$2622 s$2623 sky130_fd_sc_hd__fa_1
XFILLER_170_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1340_ clknet_leaf_0_clk booth_b12_m18 VGND VGND VPWR VPWR pp_row30_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_69_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1271_ clknet_leaf_120_clk booth_b56_m47 VGND VGND VPWR VPWR pp_row103_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_3_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0222_ clknet_leaf_126_clk notsign$6154 VGND VGND VPWR VPWR pp_row113_0 sky130_fd_sc_hd__dfxtp_1
XFILLER_37_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_1013 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$380 net1683 net534 net1658 net807 VGND VGND VPWR VPWR t$4599 sky130_fd_sc_hd__a22o_1
XU$$391 t$4604 net1276 VGND VGND VPWR VPWR booth_b4_m55 sky130_fd_sc_hd__xor2_1
XFILLER_189_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0986_ clknet_leaf_115_clk booth_b48_m52 VGND VGND VPWR VPWR pp_row100_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_118_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_8_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_191_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1607_ clknet_leaf_240_clk booth_b12_m30 VGND VGND VPWR VPWR pp_row42_6 sky130_fd_sc_hd__dfxtp_1
XFILLER_172_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1538_ clknet_leaf_8_clk booth_b20_m19 VGND VGND VPWR VPWR pp_row39_10 sky130_fd_sc_hd__dfxtp_1
XFILLER_114_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_62_5 pp_row62_32 pp_row62_33 c$50 VGND VGND VPWR VPWR c$574 s$575 sky130_fd_sc_hd__fa_1
X_1469_ clknet_leaf_39_clk booth_b22_m14 VGND VGND VPWR VPWR pp_row36_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_80_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_55_4 pp_row55_17 pp_row55_18 pp_row55_19 VGND VGND VPWR VPWR c$446 s$447
+ sky130_fd_sc_hd__fa_1
XFILLER_67_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_48_3 pp_row48_9 pp_row48_10 pp_row48_11 VGND VGND VPWR VPWR c$322 s$323
+ sky130_fd_sc_hd__fa_1
XFILLER_43_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_25_2 s$2041 s$2043 s$2045 VGND VGND VPWR VPWR c$2844 s$2845 sky130_fd_sc_hd__fa_1
XFILLER_83_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_18_1 pp_row18_11 c$1982 c$1984 VGND VGND VPWR VPWR c$2800 s$2801 sky130_fd_sc_hd__fa_1
XFILLER_179_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_761 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4253_1808 VGND VGND VPWR VPWR U$$4253_1808/HI net1808 sky130_fd_sc_hd__conb_1
XFILLER_151_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1603 net117 VGND VGND VPWR VPWR net1603 sky130_fd_sc_hd__clkbuf_4
XFILLER_105_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1614 net115 VGND VGND VPWR VPWR net1614 sky130_fd_sc_hd__buf_4
Xfanout1625 net1626 VGND VGND VPWR VPWR net1625 sky130_fd_sc_hd__buf_2
Xfanout1636 net1637 VGND VGND VPWR VPWR net1636 sky130_fd_sc_hd__clkbuf_4
XFILLER_144_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1647 net1648 VGND VGND VPWR VPWR net1647 sky130_fd_sc_hd__buf_6
XFILLER_120_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1658 net110 VGND VGND VPWR VPWR net1658 sky130_fd_sc_hd__buf_2
Xfanout660 net666 VGND VGND VPWR VPWR net660 sky130_fd_sc_hd__buf_6
XU$$4106 t$6502 net1285 VGND VGND VPWR VPWR booth_b58_m63 sky130_fd_sc_hd__xor2_1
Xfanout671 net672 VGND VGND VPWR VPWR net671 sky130_fd_sc_hd__buf_2
Xdadda_ha_3_21_3 pp_row21_9 pp_row21_10 VGND VGND VPWR VPWR c$2012 s$2013 sky130_fd_sc_hd__ha_1
Xfanout1669 net1670 VGND VGND VPWR VPWR net1669 sky130_fd_sc_hd__buf_8
XFILLER_19_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4117 t$6509 net1263 VGND VGND VPWR VPWR booth_b60_m0 sky130_fd_sc_hd__xor2_1
XFILLER_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_777 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4128 net1567 net438 net1525 net720 VGND VGND VPWR VPWR t$6515 sky130_fd_sc_hd__a22o_1
Xfanout682 net683 VGND VGND VPWR VPWR net682 sky130_fd_sc_hd__buf_4
Xfanout693 net694 VGND VGND VPWR VPWR net693 sky130_fd_sc_hd__clkbuf_4
XU$$4139 t$6520 net1264 VGND VGND VPWR VPWR booth_b60_m11 sky130_fd_sc_hd__xor2_1
XFILLER_59_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3405 t$6144 net1340 VGND VGND VPWR VPWR booth_b48_m55 sky130_fd_sc_hd__xor2_1
XU$$3416 net1556 net499 net1548 net772 VGND VGND VPWR VPWR t$6150 sky130_fd_sc_hd__a22o_1
XFILLER_46_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3427 net1330 VGND VGND VPWR VPWR notblock$6155\[2\] sky130_fd_sc_hd__inv_1
XTAP_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3438 t$6162 net1333 VGND VGND VPWR VPWR booth_b50_m3 sky130_fd_sc_hd__xor2_1
XTAP_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2704 t$5786 net1396 VGND VGND VPWR VPWR booth_b38_m47 sky130_fd_sc_hd__xor2_1
XU$$3449 net1507 net484 net1498 net757 VGND VGND VPWR VPWR t$6168 sky130_fd_sc_hd__a22o_1
XTAP_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2715 net1643 net548 net1634 net821 VGND VGND VPWR VPWR t$5792 sky130_fd_sc_hd__a22o_1
XU$$2726 t$5797 net1400 VGND VGND VPWR VPWR booth_b38_m58 sky130_fd_sc_hd__xor2_1
XTAP_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2737 net1534 net548 net1781 net821 VGND VGND VPWR VPWR t$5803 sky130_fd_sc_hd__a22o_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2748 net1227 net535 net1122 net808 VGND VGND VPWR VPWR t$5810 sky130_fd_sc_hd__a22o_1
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_20_1 pp_row20_3 pp_row20_4 pp_row20_5 VGND VGND VPWR VPWR c$2000 s$2001
+ sky130_fd_sc_hd__fa_1
XU$$2759 t$5815 net1377 VGND VGND VPWR VPWR booth_b40_m6 sky130_fd_sc_hd__xor2_1
XTAP_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0840_ clknet_leaf_105_clk booth_b32_m61 VGND VGND VPWR VPWR pp_row93_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_169_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0771_ clknet_leaf_144_clk booth_b30_m60 VGND VGND VPWR VPWR pp_row90_3 sky130_fd_sc_hd__dfxtp_1
XFILLER_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2441_ clknet_leaf_98_clk booth_b60_m7 VGND VGND VPWR VPWR pp_row67_30 sky130_fd_sc_hd__dfxtp_1
XFILLER_29_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_72_4 s$749 s$751 s$753 VGND VGND VPWR VPWR c$1598 s$1599 sky130_fd_sc_hd__fa_1
XFILLER_97_923 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2372_ clknet_leaf_85_clk booth_b4_m62 VGND VGND VPWR VPWR pp_row66_2 sky130_fd_sc_hd__dfxtp_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1323_ clknet_leaf_1_clk booth_b14_m15 VGND VGND VPWR VPWR pp_row29_7 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_65_3 c$616 s$619 s$621 VGND VGND VPWR VPWR c$1512 s$1513 sky130_fd_sc_hd__fa_1
XFILLER_151_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_58_2 c$484 c$486 c$488 VGND VGND VPWR VPWR c$1426 s$1427 sky130_fd_sc_hd__fa_1
X_1254_ clknet_leaf_10_clk booth_b14_m11 VGND VGND VPWR VPWR pp_row25_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_84_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_35_1 s$2901 s$2903 s$2905 VGND VGND VPWR VPWR c$3538 s$3539 sky130_fd_sc_hd__fa_1
XFILLER_49_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0205_ clknet_leaf_152_clk booth_b50_m20 VGND VGND VPWR VPWR pp_row70_23 sky130_fd_sc_hd__dfxtp_1
X_1185_ clknet_leaf_46_clk net1487 VGND VGND VPWR VPWR pp_row20_11 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_28_0 c$2852 c$2854 c$2856 VGND VGND VPWR VPWR c$3508 s$3509 sky130_fd_sc_hd__fa_1
XU$$3950 net1634 net465 net1624 net738 VGND VGND VPWR VPWR t$6423 sky130_fd_sc_hd__a22o_1
XU$$3961 t$6428 net1292 VGND VGND VPWR VPWR booth_b56_m59 sky130_fd_sc_hd__xor2_1
XFILLER_65_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3972 net1293 VGND VGND VPWR VPWR notsign$6434 sky130_fd_sc_hd__inv_1
XU$$3983 net1125 net451 net1034 net724 VGND VGND VPWR VPWR t$6441 sky130_fd_sc_hd__a22o_1
XU$$3994 t$6446 net1287 VGND VGND VPWR VPWR booth_b58_m7 sky130_fd_sc_hd__xor2_1
XFILLER_80_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0969_ clknet_leaf_116_clk booth_b48_m51 VGND VGND VPWR VPWR pp_row99_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_146_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$819_1886 VGND VGND VPWR VPWR U$$819_1886/HI net1886 sky130_fd_sc_hd__conb_1
XFILLER_174_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_102_0 c$3296 c$3298 c$3300 VGND VGND VPWR VPWR c$3804 s$3805 sky130_fd_sc_hd__fa_1
XFILLER_106_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput263 net263 VGND VGND VPWR VPWR o[105] sky130_fd_sc_hd__buf_2
XFILLER_88_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput274 net274 VGND VGND VPWR VPWR o[115] sky130_fd_sc_hd__buf_2
Xoutput285 net285 VGND VGND VPWR VPWR o[125] sky130_fd_sc_hd__buf_2
XFILLER_114_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput296 net296 VGND VGND VPWR VPWR o[1] sky130_fd_sc_hd__buf_2
XFILLER_59_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_250_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_250_clk
+ sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_1_60_2 pp_row60_20 pp_row60_21 pp_row60_22 VGND VGND VPWR VPWR c$532 s$533
+ sky130_fd_sc_hd__fa_1
XFILLER_87_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_53_1 pp_row53_5 pp_row53_6 pp_row53_7 VGND VGND VPWR VPWR c$404 s$405
+ sky130_fd_sc_hd__fa_1
XFILLER_74_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_30_0 s$1099 c$2070 c$2072 VGND VGND VPWR VPWR c$2870 s$2871 sky130_fd_sc_hd__fa_1
Xdadda_fa_1_46_0 pp_row46_0 pp_row46_1 pp_row46_2 VGND VGND VPWR VPWR c$288 s$289
+ sky130_fd_sc_hd__fa_2
XFILLER_28_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_82_3 s$1715 s$1717 s$1719 VGND VGND VPWR VPWR c$2500 s$2501 sky130_fd_sc_hd__fa_1
XFILLER_174_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_75_2 c$1624 s$1627 s$1629 VGND VGND VPWR VPWR c$2442 s$2443 sky130_fd_sc_hd__fa_1
XFILLER_97_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_839 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1400 net1401 VGND VGND VPWR VPWR net1400 sky130_fd_sc_hd__buf_6
Xfanout1411 net31 VGND VGND VPWR VPWR net1411 sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_3_68_1 c$1534 c$1536 c$1538 VGND VGND VPWR VPWR c$2384 s$2385 sky130_fd_sc_hd__fa_1
XFILLER_2_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1422 net1429 VGND VGND VPWR VPWR net1422 sky130_fd_sc_hd__buf_6
XU$$4411_1826 VGND VGND VPWR VPWR U$$4411_1826/HI net1826 sky130_fd_sc_hd__conb_1
Xdadda_fa_6_45_0 c$3572 c$3574 s$3577 VGND VGND VPWR VPWR c$3986 s$3987 sky130_fd_sc_hd__fa_2
Xfanout1433 net1438 VGND VGND VPWR VPWR net1433 sky130_fd_sc_hd__buf_8
Xclkbuf_leaf_241_clk clknet_5_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_241_clk
+ sky130_fd_sc_hd__clkbuf_16
Xfanout1444 net1445 VGND VGND VPWR VPWR net1444 sky130_fd_sc_hd__buf_6
Xfanout1455 net1456 VGND VGND VPWR VPWR net1455 sky130_fd_sc_hd__buf_6
Xfanout1466 net1468 VGND VGND VPWR VPWR net1466 sky130_fd_sc_hd__buf_6
XFILLER_4_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1477 net16 VGND VGND VPWR VPWR net1477 sky130_fd_sc_hd__buf_6
XFILLER_78_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout490 net491 VGND VGND VPWR VPWR net490 sky130_fd_sc_hd__buf_4
Xfanout1488 net1489 VGND VGND VPWR VPWR net1488 sky130_fd_sc_hd__clkbuf_4
XU$$3202 t$6041 net1354 VGND VGND VPWR VPWR booth_b46_m22 sky130_fd_sc_hd__xor2_1
XFILLER_65_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1499 net1501 VGND VGND VPWR VPWR net1499 sky130_fd_sc_hd__buf_4
XU$$3213 net1059 net501 net1054 net774 VGND VGND VPWR VPWR t$6047 sky130_fd_sc_hd__a22o_1
XU$$3224 t$6052 net1350 VGND VGND VPWR VPWR booth_b46_m33 sky130_fd_sc_hd__xor2_1
XU$$3235 net950 net503 net942 net776 VGND VGND VPWR VPWR t$6058 sky130_fd_sc_hd__a22o_1
XU$$2501 t$5683 net1406 VGND VGND VPWR VPWR booth_b36_m14 sky130_fd_sc_hd__xor2_1
XFILLER_0_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$17 c$4184 s$4187 VGND VGND VPWR VPWR final_adder.$signal$36 final_adder.$signal$1107
+ sky130_fd_sc_hd__ha_1
XFILLER_0_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3246 t$6063 net1356 VGND VGND VPWR VPWR booth_b46_m44 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$28 c$4206 s$4209 VGND VGND VPWR VPWR final_adder.$signal$58 final_adder.$signal$1118
+ sky130_fd_sc_hd__ha_1
XU$$3257 net1684 net507 net1660 net780 VGND VGND VPWR VPWR t$6069 sky130_fd_sc_hd__a22o_1
XU$$2512 net1134 net554 net1118 net827 VGND VGND VPWR VPWR t$5689 sky130_fd_sc_hd__a22o_1
XFILLER_185_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3268 t$6074 net1355 VGND VGND VPWR VPWR booth_b46_m55 sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_104_2 s$2673 s$2675 s$2677 VGND VGND VPWR VPWR c$3318 s$3319 sky130_fd_sc_hd__fa_1
XU$$2523 t$5694 net1405 VGND VGND VPWR VPWR booth_b36_m25 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$39 c$4228 s$4231 VGND VGND VPWR VPWR final_adder.$signal$80 final_adder.$signal$1129
+ sky130_fd_sc_hd__ha_1
XU$$2534 net1029 net559 net1021 net832 VGND VGND VPWR VPWR t$5700 sky130_fd_sc_hd__a22o_1
XFILLER_34_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3279 net1555 net508 net1547 net781 VGND VGND VPWR VPWR t$6080 sky130_fd_sc_hd__a22o_1
XU$$2545 t$5705 net1409 VGND VGND VPWR VPWR booth_b36_m36 sky130_fd_sc_hd__xor2_1
XU$$1800 t$5325 net1460 VGND VGND VPWR VPWR booth_b26_m6 sky130_fd_sc_hd__xor2_1
XU$$2556 net1748 net556 net1739 net829 VGND VGND VPWR VPWR t$5711 sky130_fd_sc_hd__a22o_1
XU$$1811 net1211 net596 net1203 net869 VGND VGND VPWR VPWR t$5331 sky130_fd_sc_hd__a22o_1
XU$$1822 t$5336 net1457 VGND VGND VPWR VPWR booth_b26_m17 sky130_fd_sc_hd__xor2_1
XFILLER_62_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2567 t$5716 net1409 VGND VGND VPWR VPWR booth_b36_m47 sky130_fd_sc_hd__xor2_1
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2578 net1640 net555 net1632 net828 VGND VGND VPWR VPWR t$5722 sky130_fd_sc_hd__a22o_1
XU$$1833 net1098 net593 net1090 net866 VGND VGND VPWR VPWR t$5342 sky130_fd_sc_hd__a22o_1
XU$$2589 t$5727 net1410 VGND VGND VPWR VPWR booth_b36_m58 sky130_fd_sc_hd__xor2_1
XU$$1844 t$5347 net1461 VGND VGND VPWR VPWR booth_b26_m28 sky130_fd_sc_hd__xor2_1
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1855 net991 net597 net983 net870 VGND VGND VPWR VPWR t$5353 sky130_fd_sc_hd__a22o_1
XU$$1866 t$5358 net1462 VGND VGND VPWR VPWR booth_b26_m39 sky130_fd_sc_hd__xor2_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1877 net1721 net598 net1712 net871 VGND VGND VPWR VPWR t$5364 sky130_fd_sc_hd__a22o_1
XFILLER_187_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1941_ clknet_leaf_72_clk booth_b46_m7 VGND VGND VPWR VPWR pp_row53_23 sky130_fd_sc_hd__dfxtp_1
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1888 t$5369 net1464 VGND VGND VPWR VPWR booth_b26_m50 sky130_fd_sc_hd__xor2_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1899 net1613 net599 net1605 net872 VGND VGND VPWR VPWR t$5375 sky130_fd_sc_hd__a22o_1
XFILLER_14_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1872_ clknet_leaf_134_clk booth_b56_m51 VGND VGND VPWR VPWR pp_row107_7 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_7_118_0 s$3871 c$4130 s$4133 VGND VGND VPWR VPWR c$4388 s$4389 sky130_fd_sc_hd__fa_1
X_0823_ clknet_leaf_108_clk booth_b42_m50 VGND VGND VPWR VPWR pp_row92_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_162_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0754_ clknet_leaf_160_clk booth_b42_m47 VGND VGND VPWR VPWR pp_row89_9 sky130_fd_sc_hd__dfxtp_1
XFILLER_171_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0685_ clknet_leaf_174_clk booth_b52_m34 VGND VGND VPWR VPWR pp_row86_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_142_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2424_ clknet_leaf_98_clk booth_b30_m37 VGND VGND VPWR VPWR pp_row67_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_9_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_70_1 c$694 c$696 c$698 VGND VGND VPWR VPWR c$1568 s$1569 sky130_fd_sc_hd__fa_2
XFILLER_9_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2355_ clknet_leaf_75_clk booth_b40_m25 VGND VGND VPWR VPWR pp_row65_20 sky130_fd_sc_hd__dfxtp_1
XFILLER_96_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_63_0 s$83 c$564 c$566 VGND VGND VPWR VPWR c$1482 s$1483 sky130_fd_sc_hd__fa_1
Xclkbuf_leaf_232_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_232_clk
+ sky130_fd_sc_hd__clkbuf_16
X_1306_ clknet_leaf_1_clk booth_b16_m12 VGND VGND VPWR VPWR pp_row28_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_9_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$518 final_adder.p_new$530 final_adder.p_new$522 VGND VGND VPWR VPWR
+ final_adder.p_new$646 sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$529 final_adder.p_new$532 final_adder.g_new$541 final_adder.g_new$533
+ VGND VGND VPWR VPWR final_adder.g_new$657 sky130_fd_sc_hd__a21o_1
XFILLER_42_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2286_ clknet_leaf_216_clk booth_b46_m17 VGND VGND VPWR VPWR pp_row63_23 sky130_fd_sc_hd__dfxtp_1
XFILLER_111_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1237_ clknet_leaf_13_clk booth_b14_m10 VGND VGND VPWR VPWR pp_row24_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_84_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4470 net946 sel_0$6647 net930 net697 VGND VGND VPWR VPWR t$6689 sky130_fd_sc_hd__a22o_1
XU$$4481 t$6694 net1861 VGND VGND VPWR VPWR booth_b64_m45 sky130_fd_sc_hd__xor2_1
XU$$4492 net1661 sel_0$6647 net1653 net697 VGND VGND VPWR VPWR t$6700 sky130_fd_sc_hd__a22o_1
XFILLER_65_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1168_ clknet_leaf_46_clk booth_b16_m3 VGND VGND VPWR VPWR pp_row19_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_53_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3780 t$6336 net1304 VGND VGND VPWR VPWR booth_b54_m37 sky130_fd_sc_hd__xor2_1
XU$$3791 net1742 net474 net1734 net747 VGND VGND VPWR VPWR t$6342 sky130_fd_sc_hd__a22o_1
X_1099_ clknet_leaf_52_clk booth_b10_m3 VGND VGND VPWR VPWR pp_row13_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_193_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_92_2 s$2577 s$2579 s$2581 VGND VGND VPWR VPWR c$3246 s$3247 sky130_fd_sc_hd__fa_1
XFILLER_193_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_85_1 c$2514 c$2516 s$2519 VGND VGND VPWR VPWR c$3202 s$3203 sky130_fd_sc_hd__fa_1
XFILLER_109_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_62_0 s$3647 c$4018 s$4021 VGND VGND VPWR VPWR c$4276 s$4277 sky130_fd_sc_hd__fa_1
XFILLER_192_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_78_0 s$1673 c$2454 c$2456 VGND VGND VPWR VPWR c$3158 s$3159 sky130_fd_sc_hd__fa_1
XFILLER_0_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1084 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_223_clk clknet_5_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_223_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_75_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$902 net964 net395 net956 net661 VGND VGND VPWR VPWR t$4866 sky130_fd_sc_hd__a22o_1
XFILLER_84_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$913 t$4871 net1314 VGND VGND VPWR VPWR booth_b12_m42 sky130_fd_sc_hd__xor2_1
XFILLER_18_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$924 net1697 net400 net1689 net666 VGND VGND VPWR VPWR t$4877 sky130_fd_sc_hd__a22o_1
XFILLER_29_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$935 t$4882 net1318 VGND VGND VPWR VPWR booth_b12_m53 sky130_fd_sc_hd__xor2_1
XU$$946 net1586 net395 net1578 net661 VGND VGND VPWR VPWR t$4888 sky130_fd_sc_hd__a22o_1
XFILLER_16_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$957 t$4893 net1316 VGND VGND VPWR VPWR booth_b12_m64 sky130_fd_sc_hd__xor2_1
XFILLER_28_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1107 t$4971 net1009 VGND VGND VPWR VPWR booth_b16_m2 sky130_fd_sc_hd__xor2_1
XU$$968 t$4900 net1185 VGND VGND VPWR VPWR booth_b14_m1 sky130_fd_sc_hd__xor2_1
XU$$1118 net1513 net643 net1505 net916 VGND VGND VPWR VPWR t$4977 sky130_fd_sc_hd__a22o_1
XU$$979 net1523 net387 net1515 net653 VGND VGND VPWR VPWR t$4906 sky130_fd_sc_hd__a22o_1
XFILLER_189_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1129 t$4982 net1006 VGND VGND VPWR VPWR booth_b16_m13 sky130_fd_sc_hd__xor2_1
XFILLER_16_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_1022 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_80_0 s$905 c$1674 c$1676 VGND VGND VPWR VPWR c$2478 s$2479 sky130_fd_sc_hd__fa_1
XFILLER_3_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0470_ clknet_leaf_192_clk booth_b64_m14 VGND VGND VPWR VPWR pp_row78_26 sky130_fd_sc_hd__dfxtp_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_214_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_214_clk
+ sky130_fd_sc_hd__clkbuf_16
Xfanout1230 net1232 VGND VGND VPWR VPWR net1230 sky130_fd_sc_hd__clkbuf_4
XFILLER_39_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1241 net1243 VGND VGND VPWR VPWR net1241 sky130_fd_sc_hd__buf_8
XFILLER_152_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2140_ clknet_leaf_33_clk booth_b44_m15 VGND VGND VPWR VPWR pp_row59_22 sky130_fd_sc_hd__dfxtp_1
XFILLER_94_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1252 net1253 VGND VGND VPWR VPWR net1252 sky130_fd_sc_hd__clkbuf_8
Xfanout1263 net58 VGND VGND VPWR VPWR net1263 sky130_fd_sc_hd__buf_6
Xfanout1274 net1276 VGND VGND VPWR VPWR net1274 sky130_fd_sc_hd__buf_6
Xfanout1285 net1286 VGND VGND VPWR VPWR net1285 sky130_fd_sc_hd__buf_4
XFILLER_93_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1296 net1299 VGND VGND VPWR VPWR net1296 sky130_fd_sc_hd__buf_6
XU$$3010 t$5942 net1374 VGND VGND VPWR VPWR booth_b42_m63 sky130_fd_sc_hd__xor2_1
XFILLER_66_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2071_ clknet_leaf_35_clk booth_b44_m13 VGND VGND VPWR VPWR pp_row57_22 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_42_5 s$247 s$249 s$251 VGND VGND VPWR VPWR c$1240 s$1241 sky130_fd_sc_hd__fa_2
XFILLER_35_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3021 t$5949 net1357 VGND VGND VPWR VPWR booth_b44_m0 sky130_fd_sc_hd__xor2_1
XU$$3032 net1565 net514 net1524 net787 VGND VGND VPWR VPWR t$5955 sky130_fd_sc_hd__a22o_1
XU$$3043 t$5960 net1362 VGND VGND VPWR VPWR booth_b44_m11 sky130_fd_sc_hd__xor2_1
X_1022_ clknet_leaf_60_clk booth_b0_m2 VGND VGND VPWR VPWR pp_row2_0 sky130_fd_sc_hd__dfxtp_1
XU$$3054 net1159 net510 net1151 net783 VGND VGND VPWR VPWR t$5966 sky130_fd_sc_hd__a22o_1
XFILLER_81_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2320 net1555 net575 net1547 net848 VGND VGND VPWR VPWR t$5590 sky130_fd_sc_hd__a22o_1
XU$$3065 t$5971 net1362 VGND VGND VPWR VPWR booth_b44_m22 sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_35_4 pp_row35_14 pp_row35_15 pp_row35_16 VGND VGND VPWR VPWR c$1154 s$1155
+ sky130_fd_sc_hd__fa_1
XU$$2331 net1426 VGND VGND VPWR VPWR notblock$5595\[2\] sky130_fd_sc_hd__inv_1
XU$$3076 net1059 net510 net1048 net783 VGND VGND VPWR VPWR t$5977 sky130_fd_sc_hd__a22o_1
XFILLER_179_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3087 t$5982 net1357 VGND VGND VPWR VPWR booth_b44_m33 sky130_fd_sc_hd__xor2_1
XU$$2342 t$5602 net1423 VGND VGND VPWR VPWR booth_b34_m3 sky130_fd_sc_hd__xor2_1
XU$$3098 net950 net512 net942 net785 VGND VGND VPWR VPWR t$5988 sky130_fd_sc_hd__a22o_1
XU$$2353 net1504 net560 net1495 net833 VGND VGND VPWR VPWR t$5608 sky130_fd_sc_hd__a22o_1
XU$$2364 t$5613 net1420 VGND VGND VPWR VPWR booth_b34_m14 sky130_fd_sc_hd__xor2_1
XU$$2375 net1134 net564 net1118 net837 VGND VGND VPWR VPWR t$5619 sky130_fd_sc_hd__a22o_1
XU$$1630 t$5237 net1482 VGND VGND VPWR VPWR booth_b22_m58 sky130_fd_sc_hd__xor2_1
XFILLER_34_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1641 net1528 net617 net1764 net890 VGND VGND VPWR VPWR t$5243 sky130_fd_sc_hd__a22o_1
XU$$2386 t$5624 net1421 VGND VGND VPWR VPWR booth_b34_m25 sky130_fd_sc_hd__xor2_1
XU$$2397 net1026 net564 net1018 net837 VGND VGND VPWR VPWR t$5630 sky130_fd_sc_hd__a22o_1
XU$$1652 net1228 net602 net1122 net875 VGND VGND VPWR VPWR t$5250 sky130_fd_sc_hd__a22o_1
XU$$1663 t$5255 net1466 VGND VGND VPWR VPWR booth_b24_m6 sky130_fd_sc_hd__xor2_1
XFILLER_50_848 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1674 net1216 net606 net1206 net879 VGND VGND VPWR VPWR t$5261 sky130_fd_sc_hd__a22o_1
XU$$1685 t$5266 net1466 VGND VGND VPWR VPWR booth_b24_m17 sky130_fd_sc_hd__xor2_1
XU$$1696 net1098 net604 net1090 net877 VGND VGND VPWR VPWR t$5272 sky130_fd_sc_hd__a22o_1
XFILLER_91_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1924_ clknet_leaf_65_clk booth_b16_m37 VGND VGND VPWR VPWR pp_row53_8 sky130_fd_sc_hd__dfxtp_1
XFILLER_187_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1855_ clknet_leaf_68_clk booth_b2_m49 VGND VGND VPWR VPWR pp_row51_1 sky130_fd_sc_hd__dfxtp_1
XFILLER_163_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_95_0 c$3254 c$3256 c$3258 VGND VGND VPWR VPWR c$3776 s$3777 sky130_fd_sc_hd__fa_1
XFILLER_135_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0806_ clknet_leaf_106_clk booth_b52_m39 VGND VGND VPWR VPWR pp_row91_13 sky130_fd_sc_hd__dfxtp_1
X_1786_ clknet_leaf_222_clk booth_b40_m8 VGND VGND VPWR VPWR pp_row48_20 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0737_ clknet_leaf_134_clk booth_b54_m34 VGND VGND VPWR VPWR pp_row88_16 sky130_fd_sc_hd__dfxtp_1
XFILLER_171_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0668_ clknet_leaf_184_clk net240 VGND VGND VPWR VPWR pp_row85_23 sky130_fd_sc_hd__dfxtp_1
X_2407_ clknet_leaf_198_clk net219 VGND VGND VPWR VPWR pp_row66_33 sky130_fd_sc_hd__dfxtp_2
XFILLER_97_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0599_ clknet_leaf_126_clk booth_b64_m52 VGND VGND VPWR VPWR pp_row116_7 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_205_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_205_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$304 final_adder.p_new$306 final_adder.p_new$304 VGND VGND VPWR VPWR
+ final_adder.p_new$432 sky130_fd_sc_hd__and2_1
X_2338_ clknet_leaf_91_clk booth_b8_m57 VGND VGND VPWR VPWR pp_row65_4 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$315 final_adder.p_new$314 final_adder.g_new$317 final_adder.g_new$315
+ VGND VGND VPWR VPWR final_adder.g_new$443 sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$326 final_adder.p_new$328 final_adder.p_new$326 VGND VGND VPWR VPWR
+ final_adder.p_new$454 sky130_fd_sc_hd__and2_1
XFILLER_58_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$337 final_adder.p_new$336 final_adder.g_new$339 final_adder.g_new$337
+ VGND VGND VPWR VPWR final_adder.g_new$465 sky130_fd_sc_hd__a21o_1
XTAP_3619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$348 final_adder.p_new$350 final_adder.p_new$348 VGND VGND VPWR VPWR
+ final_adder.p_new$476 sky130_fd_sc_hd__and2_1
XFILLER_55_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2269_ clknet_leaf_210_clk booth_b18_m45 VGND VGND VPWR VPWR pp_row63_9 sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$359 final_adder.p_new$358 final_adder.g_new$361 final_adder.g_new$359
+ VGND VGND VPWR VPWR final_adder.g_new$487 sky130_fd_sc_hd__a21o_1
XU$$209 net1000 net623 net992 net896 VGND VGND VPWR VPWR t$4512 sky130_fd_sc_hd__a22o_1
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_758 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_111_2 pp_row111_6 pp_row111_7 pp_row111_8 VGND VGND VPWR VPWR c$2730 s$2731
+ sky130_fd_sc_hd__fa_1
XFILLER_107_633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_104_1 pp_row104_11 pp_row104_12 pp_row104_13 VGND VGND VPWR VPWR c$2672
+ s$2673 sky130_fd_sc_hd__fa_1
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_125_0 pp_row125_3 c$3892 c$3894 VGND VGND VPWR VPWR c$4146 s$4147 sky130_fd_sc_hd__fa_2
Xdadda_fa_0_68_4 pp_row68_12 pp_row68_13 pp_row68_14 VGND VGND VPWR VPWR c$140 s$141
+ sky130_fd_sc_hd__fa_1
XFILLER_48_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_45_3 s$1271 s$1273 s$1275 VGND VGND VPWR VPWR c$2204 s$2205 sky130_fd_sc_hd__fa_1
XFILLER_91_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$710 t$4768 net1414 VGND VGND VPWR VPWR booth_b10_m9 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$871 final_adder.p_new$902 final_adder.g_new$855 final_adder.g_new$903
+ VGND VGND VPWR VPWR final_adder.g_new$999 sky130_fd_sc_hd__a21o_1
XFILLER_57_992 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_38_2 c$1180 s$1183 s$1185 VGND VGND VPWR VPWR c$2146 s$2147 sky130_fd_sc_hd__fa_1
XU$$721 net1174 net402 net1164 net668 VGND VGND VPWR VPWR t$4774 sky130_fd_sc_hd__a22o_1
XU$$732 t$4779 net1412 VGND VGND VPWR VPWR booth_b10_m20 sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$893 final_adder.p_new$924 final_adder.g_new$633 final_adder.g_new$925
+ VGND VGND VPWR VPWR final_adder.g_new$1021 sky130_fd_sc_hd__a21o_1
XU$$743 net1074 net405 net1066 net671 VGND VGND VPWR VPWR t$4785 sky130_fd_sc_hd__a22o_1
XU$$754 t$4790 net1413 VGND VGND VPWR VPWR booth_b10_m31 sky130_fd_sc_hd__xor2_1
XFILLER_17_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$765 net964 net401 net956 net667 VGND VGND VPWR VPWR t$4796 sky130_fd_sc_hd__a22o_1
XU$$776 t$4801 net1416 VGND VGND VPWR VPWR booth_b10_m42 sky130_fd_sc_hd__xor2_1
XU$$787 net1698 net407 net1690 net673 VGND VGND VPWR VPWR t$4807 sky130_fd_sc_hd__a22o_1
XU$$798 t$4812 net1418 VGND VGND VPWR VPWR booth_b10_m53 sky130_fd_sc_hd__xor2_1
XFILLER_182_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1640_ clknet_leaf_240_clk booth_b22_m21 VGND VGND VPWR VPWR pp_row43_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_184_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_4 c$4188 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1571_ clknet_leaf_20_clk booth_b38_m2 VGND VGND VPWR VPWR pp_row40_19 sky130_fd_sc_hd__dfxtp_1
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0522_ clknet_leaf_181_clk net146 VGND VGND VPWR VPWR pp_row115_8 sky130_fd_sc_hd__dfxtp_2
XFILLER_99_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0453_ clknet_leaf_158_clk booth_b34_m44 VGND VGND VPWR VPWR pp_row78_11 sky130_fd_sc_hd__dfxtp_1
XFILLER_112_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0384_ clknet_leaf_193_clk booth_b20_m56 VGND VGND VPWR VPWR pp_row76_5 sky130_fd_sc_hd__dfxtp_1
Xfanout1060 net1062 VGND VGND VPWR VPWR net1060 sky130_fd_sc_hd__buf_4
Xdadda_ha_2_27_2 pp_row27_6 pp_row27_7 VGND VGND VPWR VPWR c$1072 s$1073 sky130_fd_sc_hd__ha_1
Xfanout1071 net1072 VGND VGND VPWR VPWR net1071 sky130_fd_sc_hd__buf_4
X_2123_ clknet_leaf_219_clk booth_b14_m45 VGND VGND VPWR VPWR pp_row59_7 sky130_fd_sc_hd__dfxtp_1
Xfanout1082 net81 VGND VGND VPWR VPWR net1082 sky130_fd_sc_hd__buf_6
Xfanout1093 net80 VGND VGND VPWR VPWR net1093 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_40_2 pp_row40_17 pp_row40_18 pp_row40_19 VGND VGND VPWR VPWR c$1210 s$1211
+ sky130_fd_sc_hd__fa_1
X_2054_ clknet_leaf_38_clk booth_b14_m43 VGND VGND VPWR VPWR pp_row57_7 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_2_33_1 pp_row33_3 pp_row33_4 pp_row33_5 VGND VGND VPWR VPWR c$1124 s$1125
+ sky130_fd_sc_hd__fa_1
X_1005_ clknet_leaf_118_clk booth_b50_m51 VGND VGND VPWR VPWR pp_row101_7 sky130_fd_sc_hd__dfxtp_1
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2150 t$5503 net1443 VGND VGND VPWR VPWR booth_b30_m44 sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_10_0 pp_row10_5 pp_row10_6 pp_row10_7 VGND VGND VPWR VPWR c$3436 s$3437
+ sky130_fd_sc_hd__fa_1
XFILLER_179_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4463_1852 VGND VGND VPWR VPWR U$$4463_1852/HI net1852 sky130_fd_sc_hd__conb_1
Xdadda_fa_2_26_0 pp_row26_0 pp_row26_1 pp_row26_2 VGND VGND VPWR VPWR c$1062 s$1063
+ sky130_fd_sc_hd__fa_1
XFILLER_50_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2161 net1680 net578 net1655 net851 VGND VGND VPWR VPWR t$5509 sky130_fd_sc_hd__a22o_1
XU$$2172 t$5514 net1444 VGND VGND VPWR VPWR booth_b30_m55 sky130_fd_sc_hd__xor2_1
XU$$2183 net1555 net582 net1547 net855 VGND VGND VPWR VPWR t$5520 sky130_fd_sc_hd__a22o_1
XFILLER_22_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2194 net1435 VGND VGND VPWR VPWR notblock$5525\[2\] sky130_fd_sc_hd__inv_1
XFILLER_50_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1460 net1745 net631 net1737 net904 VGND VGND VPWR VPWR t$5151 sky130_fd_sc_hd__a22o_1
XU$$1471 t$5156 net1493 VGND VGND VPWR VPWR booth_b20_m47 sky130_fd_sc_hd__xor2_1
XU$$1482 net1638 net632 net1629 net905 VGND VGND VPWR VPWR t$5162 sky130_fd_sc_hd__a22o_1
XU$$1493 t$5167 net1492 VGND VGND VPWR VPWR booth_b20_m58 sky130_fd_sc_hd__xor2_1
XFILLER_148_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1907_ clknet_leaf_70_clk booth_b42_m10 VGND VGND VPWR VPWR pp_row52_21 sky130_fd_sc_hd__dfxtp_1
XFILLER_175_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1838_ clknet_leaf_135_clk booth_b50_m57 VGND VGND VPWR VPWR pp_row107_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1769_ clknet_leaf_237_clk booth_b10_m38 VGND VGND VPWR VPWR pp_row48_5 sky130_fd_sc_hd__dfxtp_1
XFILLER_190_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_85_4 pp_row85_12 pp_row85_13 pp_row85_14 VGND VGND VPWR VPWR c$974 s$975
+ sky130_fd_sc_hd__fa_1
XFILLER_103_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_78_3 pp_row78_11 pp_row78_12 pp_row78_13 VGND VGND VPWR VPWR c$858 s$859
+ sky130_fd_sc_hd__fa_1
XFILLER_44_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_55_2 s$2281 s$2283 s$2285 VGND VGND VPWR VPWR c$3024 s$3025 sky130_fd_sc_hd__fa_1
XTAP_4106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$101 c$4352 s$4355 VGND VGND VPWR VPWR final_adder.$signal$204 final_adder.$signal$1191
+ sky130_fd_sc_hd__ha_1
XFILLER_170_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$112 c$4374 s$4377 VGND VGND VPWR VPWR final_adder.$signal$226 final_adder.$signal$1202
+ sky130_fd_sc_hd__ha_1
XTAP_4139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_48_1 c$2218 c$2220 s$2223 VGND VGND VPWR VPWR c$2980 s$2981 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$123 c$4396 s$4399 VGND VGND VPWR VPWR final_adder.$signal$248 final_adder.$signal$1213
+ sky130_fd_sc_hd__ha_2
XFILLER_111_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$134 final_adder.$signal$1210 final_adder.$signal$1211 VGND VGND VPWR
+ VPWR final_adder.p_new$262 sky130_fd_sc_hd__and2_1
XTAP_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$145 final_adder.$signal$1201 final_adder.$signal$222 final_adder.$signal$224
+ VGND VGND VPWR VPWR final_adder.g_new$273 sky130_fd_sc_hd__a21o_1
Xdadda_fa_7_25_0 s$3499 c$3944 s$3947 VGND VGND VPWR VPWR c$4202 s$4203 sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$156 final_adder.$signal$1188 final_adder.$signal$1189 VGND VGND VPWR
+ VPWR final_adder.p_new$284 sky130_fd_sc_hd__and2_1
XTAP_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$167 final_adder.$signal$1179 final_adder.$signal$178 final_adder.$signal$180
+ VGND VGND VPWR VPWR final_adder.g_new$295 sky130_fd_sc_hd__a21o_1
XTAP_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$178 final_adder.$signal$1166 final_adder.$signal$1167 VGND VGND VPWR
+ VPWR final_adder.p_new$306 sky130_fd_sc_hd__and2_1
XFILLER_26_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$189 final_adder.$signal$1157 final_adder.$signal$134 final_adder.$signal$136
+ VGND VGND VPWR VPWR final_adder.g_new$317 sky130_fd_sc_hd__a21o_1
XANTENNA_405 net1714 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_416 net400 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_427 net678 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_438 net931 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_449 net1506 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_0_73_2 pp_row73_6 pp_row73_7 pp_row73_8 VGND VGND VPWR VPWR c$184 s$185
+ sky130_fd_sc_hd__fa_1
XFILLER_1_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput130 c[100] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_1
XFILLER_163_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput141 c[110] VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_50_1 c$1318 c$1320 c$1322 VGND VGND VPWR VPWR c$2240 s$2241 sky130_fd_sc_hd__fa_1
Xinput152 c[120] VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_0_66_1 pp_row66_3 pp_row66_4 pp_row66_5 VGND VGND VPWR VPWR c$110 s$111
+ sky130_fd_sc_hd__fa_1
Xinput163 c[15] VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_1
Xinput174 c[25] VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_3_43_0 s$263 c$1230 c$1232 VGND VGND VPWR VPWR c$2182 s$2183 sky130_fd_sc_hd__fa_1
Xinput185 c[35] VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_1
Xinput196 c[45] VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_0_59_0 pp_row59_0 pp_row59_1 pp_row59_2 VGND VGND VPWR VPWR c$32 s$33 sky130_fd_sc_hd__fa_1
XFILLER_76_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$690 final_adder.p_new$714 final_adder.p_new$698 VGND VGND VPWR VPWR
+ final_adder.p_new$818 sky130_fd_sc_hd__and2_1
XTAP_3972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$540 t$4680 net1252 VGND VGND VPWR VPWR booth_b6_m61 sky130_fd_sc_hd__xor2_1
XTAP_3983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$551 net1237 notblock$4685\[1\] VGND VGND VPWR VPWR t$4686 sky130_fd_sc_hd__and2_1
XTAP_3994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$562 net937 net414 net1675 net680 VGND VGND VPWR VPWR t$4693 sky130_fd_sc_hd__a22o_1
XFILLER_44_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$573 t$4698 net1236 VGND VGND VPWR VPWR booth_b8_m9 sky130_fd_sc_hd__xor2_1
XU$$584 net1179 net415 net1170 net681 VGND VGND VPWR VPWR t$4704 sky130_fd_sc_hd__a22o_1
XFILLER_17_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$595 t$4709 net1235 VGND VGND VPWR VPWR booth_b8_m20 sky130_fd_sc_hd__xor2_1
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$956_1888 VGND VGND VPWR VPWR U$$956_1888/HI net1888 sky130_fd_sc_hd__conb_1
XFILLER_145_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_100_0 s$3799 c$4094 s$4097 VGND VGND VPWR VPWR c$4352 s$4353 sky130_fd_sc_hd__fa_1
XFILLER_68_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_95_3 pp_row95_12 pp_row95_13 pp_row95_14 VGND VGND VPWR VPWR c$1872 s$1873
+ sky130_fd_sc_hd__fa_1
X_1623_ clknet_leaf_240_clk booth_b40_m2 VGND VGND VPWR VPWR pp_row42_20 sky130_fd_sc_hd__dfxtp_1
XU$$4493_1867 VGND VGND VPWR VPWR U$$4493_1867/HI net1867 sky130_fd_sc_hd__conb_1
XFILLER_114_912 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_88_2 pp_row88_20 pp_row88_21 pp_row88_22 VGND VGND VPWR VPWR c$1786 s$1787
+ sky130_fd_sc_hd__fa_1
X_1554_ clknet_leaf_6_clk booth_b6_m34 VGND VGND VPWR VPWR pp_row40_3 sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_5_65_1 s$3081 s$3083 s$3085 VGND VGND VPWR VPWR c$3658 s$3659 sky130_fd_sc_hd__fa_1
X_0505_ clknet_leaf_172_clk booth_b20_m60 VGND VGND VPWR VPWR pp_row80_3 sky130_fd_sc_hd__dfxtp_1
X_1485_ clknet_leaf_45_clk booth_b8_m29 VGND VGND VPWR VPWR pp_row37_4 sky130_fd_sc_hd__dfxtp_1
XFILLER_154_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_58_0 c$3032 c$3034 c$3036 VGND VGND VPWR VPWR c$3628 s$3629 sky130_fd_sc_hd__fa_1
XFILLER_140_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0436_ clknet_leaf_154_clk booth_b56_m21 VGND VGND VPWR VPWR pp_row77_22 sky130_fd_sc_hd__dfxtp_1
.ends

