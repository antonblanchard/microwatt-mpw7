* NGSPICE file created from Microwatt_FP_DFFRFile.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

.subckt Microwatt_FP_DFFRFile CLK D1[0] D1[10] D1[11] D1[12] D1[13] D1[14] D1[15]
+ D1[16] D1[17] D1[18] D1[19] D1[1] D1[20] D1[21] D1[22] D1[23] D1[24] D1[25] D1[26]
+ D1[27] D1[28] D1[29] D1[2] D1[30] D1[31] D1[32] D1[33] D1[34] D1[35] D1[36] D1[37]
+ D1[38] D1[39] D1[3] D1[40] D1[41] D1[42] D1[43] D1[44] D1[45] D1[46] D1[47] D1[48]
+ D1[49] D1[4] D1[50] D1[51] D1[52] D1[53] D1[54] D1[55] D1[56] D1[57] D1[58] D1[59]
+ D1[5] D1[60] D1[61] D1[62] D1[63] D1[6] D1[7] D1[8] D1[9] D2[0] D2[10] D2[11] D2[12]
+ D2[13] D2[14] D2[15] D2[16] D2[17] D2[18] D2[19] D2[1] D2[20] D2[21] D2[22] D2[23]
+ D2[24] D2[25] D2[26] D2[27] D2[28] D2[29] D2[2] D2[30] D2[31] D2[32] D2[33] D2[34]
+ D2[35] D2[36] D2[37] D2[38] D2[39] D2[3] D2[40] D2[41] D2[42] D2[43] D2[44] D2[45]
+ D2[46] D2[47] D2[48] D2[49] D2[4] D2[50] D2[51] D2[52] D2[53] D2[54] D2[55] D2[56]
+ D2[57] D2[58] D2[59] D2[5] D2[60] D2[61] D2[62] D2[63] D2[6] D2[7] D2[8] D2[9] D3[0]
+ D3[10] D3[11] D3[12] D3[13] D3[14] D3[15] D3[16] D3[17] D3[18] D3[19] D3[1] D3[20]
+ D3[21] D3[22] D3[23] D3[24] D3[25] D3[26] D3[27] D3[28] D3[29] D3[2] D3[30] D3[31]
+ D3[32] D3[33] D3[34] D3[35] D3[36] D3[37] D3[38] D3[39] D3[3] D3[40] D3[41] D3[42]
+ D3[43] D3[44] D3[45] D3[46] D3[47] D3[48] D3[49] D3[4] D3[50] D3[51] D3[52] D3[53]
+ D3[54] D3[55] D3[56] D3[57] D3[58] D3[59] D3[5] D3[60] D3[61] D3[62] D3[63] D3[6]
+ D3[7] D3[8] D3[9] DW[0] DW[10] DW[11] DW[12] DW[13] DW[14] DW[15] DW[16] DW[17]
+ DW[18] DW[19] DW[1] DW[20] DW[21] DW[22] DW[23] DW[24] DW[25] DW[26] DW[27] DW[28]
+ DW[29] DW[2] DW[30] DW[31] DW[32] DW[33] DW[34] DW[35] DW[36] DW[37] DW[38] DW[39]
+ DW[3] DW[40] DW[41] DW[42] DW[43] DW[44] DW[45] DW[46] DW[47] DW[48] DW[49] DW[4]
+ DW[50] DW[51] DW[52] DW[53] DW[54] DW[55] DW[56] DW[57] DW[58] DW[59] DW[5] DW[60]
+ DW[61] DW[62] DW[63] DW[6] DW[7] DW[8] DW[9] R1[0] R1[1] R1[2] R1[3] R1[4] R1[5]
+ R2[0] R2[1] R2[2] R2[3] R2[4] R2[5] R3[0] R3[1] R3[2] R3[3] R3[4] R3[5] RW[0] RW[1]
+ RW[2] RW[3] RW[4] RW[5] VGND VPWR WE
X_34984_ _35624_/CLK _34984_/D VGND VGND VPWR VPWR _34984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_223_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33935_ _36113_/CLK _33935_/D VGND VGND VPWR VPWR _33935_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18869_ _18865_/X _18868_/X _18726_/X VGND VGND VPWR VPWR _18895_/A sky130_fd_sc_hd__o21ba_1
XFILLER_55_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_884 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20900_ _22469_/A VGND VGND VPWR VPWR _20900_/X sky130_fd_sc_hd__buf_4
XFILLER_243_816 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21880_ _22586_/A VGND VGND VPWR VPWR _21880_/X sky130_fd_sc_hd__buf_6
X_33866_ _36105_/CLK _33866_/D VGND VGND VPWR VPWR _33866_/Q sky130_fd_sc_hd__dfxtp_1
X_35605_ _35733_/CLK _35605_/D VGND VGND VPWR VPWR _35605_/Q sky130_fd_sc_hd__dfxtp_1
X_20831_ _20660_/X _20829_/X _20830_/X _20672_/X VGND VGND VPWR VPWR _20831_/X sky130_fd_sc_hd__a22o_1
XFILLER_36_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32817_ _35953_/CLK _32817_/D VGND VGND VPWR VPWR _32817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33797_ _36159_/CLK _33797_/D VGND VGND VPWR VPWR _33797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20762_ _20648_/X _20760_/X _20761_/X _20658_/X VGND VGND VPWR VPWR _20762_/X sky130_fd_sc_hd__a22o_1
X_23550_ _23550_/A VGND VGND VPWR VPWR _32269_/D sky130_fd_sc_hd__clkbuf_1
X_35536_ _35731_/CLK _35536_/D VGND VGND VPWR VPWR _35536_/Q sky130_fd_sc_hd__dfxtp_1
X_32748_ _32875_/CLK _32748_/D VGND VGND VPWR VPWR _32748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_243_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22501_ _22464_/X _22499_/X _22500_/X _22469_/X VGND VGND VPWR VPWR _22501_/X sky130_fd_sc_hd__a22o_1
XFILLER_17_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23481_ input54/X VGND VGND VPWR VPWR _23481_/X sky130_fd_sc_hd__buf_4
XFILLER_50_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35467_ _35723_/CLK _35467_/D VGND VGND VPWR VPWR _35467_/Q sky130_fd_sc_hd__dfxtp_1
X_20693_ _22366_/A VGND VGND VPWR VPWR _21477_/A sky130_fd_sc_hd__buf_8
X_32679_ _32871_/CLK _32679_/D VGND VGND VPWR VPWR _32679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_818 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22432_ _22152_/X _22430_/X _22431_/X _22157_/X VGND VGND VPWR VPWR _22432_/X sky130_fd_sc_hd__a22o_1
X_25220_ _33086_/Q _23420_/X _25238_/S VGND VGND VPWR VPWR _25221_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34418_ _34611_/CLK _34418_/D VGND VGND VPWR VPWR _34418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35398_ _35525_/CLK _35398_/D VGND VGND VPWR VPWR _35398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22363_ _22159_/X _22361_/X _22362_/X _22162_/X VGND VGND VPWR VPWR _22363_/X sky130_fd_sc_hd__a22o_1
XFILLER_149_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25151_ _25151_/A VGND VGND VPWR VPWR _33053_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34349_ _35630_/CLK _34349_/D VGND VGND VPWR VPWR _34349_/Q sky130_fd_sc_hd__dfxtp_1
X_24102_ _24102_/A VGND VGND VPWR VPWR _32591_/D sky130_fd_sc_hd__clkbuf_1
X_21314_ _22512_/A VGND VGND VPWR VPWR _21314_/X sky130_fd_sc_hd__clkbuf_4
X_25082_ _25130_/S VGND VGND VPWR VPWR _25101_/S sky130_fd_sc_hd__buf_6
XFILLER_108_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22294_ _22290_/X _22293_/X _22085_/X VGND VGND VPWR VPWR _22324_/A sky130_fd_sc_hd__o21ba_1
XFILLER_124_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28910_ _28910_/A VGND VGND VPWR VPWR _34767_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24033_ _24033_/A VGND VGND VPWR VPWR _32558_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21245_ _22459_/A VGND VGND VPWR VPWR _21245_/X sky130_fd_sc_hd__clkbuf_4
X_36019_ _36019_/CLK _36019_/D VGND VGND VPWR VPWR _36019_/Q sky130_fd_sc_hd__dfxtp_1
X_29890_ _29890_/A VGND VGND VPWR VPWR _35201_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28841_ _28841_/A VGND VGND VPWR VPWR _34734_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21176_ _32868_/Q _32804_/Q _32740_/Q _32676_/Q _20887_/X _20888_/X VGND VGND VPWR
+ VPWR _21176_/X sky130_fd_sc_hd__mux4_1
XFILLER_89_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20127_ _20123_/X _20126_/X _19818_/X VGND VGND VPWR VPWR _20128_/D sky130_fd_sc_hd__o21ba_1
X_28772_ _34703_/Q _27211_/X _28776_/S VGND VGND VPWR VPWR _28773_/A sky130_fd_sc_hd__mux2_1
X_25984_ _24852_/X _33447_/Q _25988_/S VGND VGND VPWR VPWR _25985_/A sky130_fd_sc_hd__mux2_1
XFILLER_246_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27723_ input19/X VGND VGND VPWR VPWR _27723_/X sky130_fd_sc_hd__buf_2
XFILLER_86_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20058_ _33670_/Q _33606_/Q _33542_/Q _33478_/Q _19853_/X _19854_/X VGND VGND VPWR
+ VPWR _20058_/X sky130_fd_sc_hd__mux4_1
X_24935_ _24935_/A VGND VGND VPWR VPWR _32961_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27654_ _27654_/A VGND VGND VPWR VPWR _34201_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24866_ _24865_/X _32939_/Q _24890_/S VGND VGND VPWR VPWR _24867_/A sky130_fd_sc_hd__mux2_1
XTAP_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26605_ _26605_/A VGND VGND VPWR VPWR _33740_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23817_ _23817_/A VGND VGND VPWR VPWR _32393_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27585_ _34172_/Q _27152_/X _27587_/S VGND VGND VPWR VPWR _27586_/A sky130_fd_sc_hd__mux2_1
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24797_ _27232_/B _25132_/A input83/X input89/X VGND VGND VPWR VPWR _24798_/A sky130_fd_sc_hd__and4b_1
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29324_ _34964_/Q _27226_/X _29326_/S VGND VGND VPWR VPWR _29325_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26536_ _26536_/A VGND VGND VPWR VPWR _33707_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23748_ _22946_/X _32361_/Q _23748_/S VGND VGND VPWR VPWR _23749_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29255_ _34931_/Q _27124_/X _29255_/S VGND VGND VPWR VPWR _29256_/A sky130_fd_sc_hd__mux2_1
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26467_ _26467_/A VGND VGND VPWR VPWR _33675_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23679_ _23679_/A VGND VGND VPWR VPWR _32329_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28206_ _27782_/X _34435_/Q _28214_/S VGND VGND VPWR VPWR _28207_/A sky130_fd_sc_hd__mux2_1
X_16220_ _16018_/X _16218_/X _16219_/X _16027_/X VGND VGND VPWR VPWR _16220_/X sky130_fd_sc_hd__a22o_1
XFILLER_9_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25418_ _25418_/A VGND VGND VPWR VPWR _33178_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29186_ _29186_/A VGND VGND VPWR VPWR _34898_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26398_ _26398_/A VGND VGND VPWR VPWR _33642_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16151_ _16147_/X _16148_/X _16149_/X _16150_/X VGND VGND VPWR VPWR _16151_/X sky130_fd_sc_hd__a22o_1
XFILLER_154_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28137_ _27680_/X _34402_/Q _28151_/S VGND VGND VPWR VPWR _28138_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25349_ _33147_/Q _23411_/X _25353_/S VGND VGND VPWR VPWR _25350_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28068_ _28068_/A VGND VGND VPWR VPWR _34369_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16082_ _17982_/A VGND VGND VPWR VPWR _17716_/A sky130_fd_sc_hd__buf_12
X_27019_ _33935_/Q _23478_/X _27023_/S VGND VGND VPWR VPWR _27020_/A sky130_fd_sc_hd__mux2_1
X_19910_ _33089_/Q _32065_/Q _35841_/Q _35777_/Q _19731_/X _19732_/X VGND VGND VPWR
+ VPWR _19910_/X sky130_fd_sc_hd__mux4_1
XFILLER_154_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30030_ _35268_/Q _29472_/X _30036_/S VGND VGND VPWR VPWR _30031_/A sky130_fd_sc_hd__mux2_1
X_19841_ _19656_/X _19839_/X _19840_/X _19659_/X VGND VGND VPWR VPWR _19841_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_218_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16984_ _16846_/X _16982_/X _16983_/X _16851_/X VGND VGND VPWR VPWR _16984_/X sky130_fd_sc_hd__a22o_1
XFILLER_7_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19772_ _34941_/Q _34877_/Q _34813_/Q _34749_/Q _19460_/X _19461_/X VGND VGND VPWR
+ VPWR _19772_/X sky130_fd_sc_hd__mux4_1
XFILLER_110_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18723_ _33376_/Q _33312_/Q _33248_/Q _33184_/Q _18721_/X _18722_/X VGND VGND VPWR
+ VPWR _18723_/X sky130_fd_sc_hd__mux4_1
XTAP_5160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31981_ _34790_/CLK _31981_/D VGND VGND VPWR VPWR _31981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30932_ _30932_/A VGND VGND VPWR VPWR _35695_/D sky130_fd_sc_hd__clkbuf_1
X_33720_ _35704_/CLK _33720_/D VGND VGND VPWR VPWR _33720_/Q sky130_fd_sc_hd__dfxtp_1
X_18654_ _20066_/A VGND VGND VPWR VPWR _18654_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_236_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_6_CLK clkbuf_leaf_9_CLK/A VGND VGND VPWR VPWR _34914_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_91_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17605_ _35649_/Q _35009_/Q _34369_/Q _33729_/Q _17497_/X _17498_/X VGND VGND VPWR
+ VPWR _17605_/X sky130_fd_sc_hd__mux4_1
XFILLER_236_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30863_ _35663_/Q input53/X _30867_/S VGND VGND VPWR VPWR _30864_/A sky130_fd_sc_hd__mux2_1
X_18585_ _18318_/X _18583_/X _18584_/X _18327_/X VGND VGND VPWR VPWR _18585_/X sky130_fd_sc_hd__a22o_1
X_33651_ _36082_/CLK _33651_/D VGND VGND VPWR VPWR _33651_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32602_ _36055_/CLK _32602_/D VGND VGND VPWR VPWR _32602_/Q sky130_fd_sc_hd__dfxtp_1
X_17536_ _35711_/Q _32221_/Q _35583_/Q _35519_/Q _17317_/X _17318_/X VGND VGND VPWR
+ VPWR _17536_/X sky130_fd_sc_hd__mux4_1
X_33582_ _33902_/CLK _33582_/D VGND VGND VPWR VPWR _33582_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_1304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30794_ _35630_/Q input17/X _30804_/S VGND VGND VPWR VPWR _30795_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_225_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32533_ _36053_/CLK _32533_/D VGND VGND VPWR VPWR _32533_/Q sky130_fd_sc_hd__dfxtp_1
X_35321_ _35448_/CLK _35321_/D VGND VGND VPWR VPWR _35321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17467_ _17463_/X _17466_/X _17151_/X VGND VGND VPWR VPWR _17475_/C sky130_fd_sc_hd__o21ba_1
XFILLER_177_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16418_ _33632_/Q _33568_/Q _33504_/Q _33440_/Q _16141_/X _16142_/X VGND VGND VPWR
+ VPWR _16418_/X sky130_fd_sc_hd__mux4_1
X_19206_ _19200_/X _19205_/X _19098_/X VGND VGND VPWR VPWR _19214_/C sky130_fd_sc_hd__o21ba_1
X_32464_ _36079_/CLK _32464_/D VGND VGND VPWR VPWR _32464_/Q sky130_fd_sc_hd__dfxtp_1
X_35252_ _35698_/CLK _35252_/D VGND VGND VPWR VPWR _35252_/Q sky130_fd_sc_hd__dfxtp_1
X_17398_ _17153_/X _17396_/X _17397_/X _17156_/X VGND VGND VPWR VPWR _17398_/X sky130_fd_sc_hd__a22o_1
XFILLER_192_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34203_ _36121_/CLK _34203_/D VGND VGND VPWR VPWR _34203_/Q sky130_fd_sc_hd__dfxtp_1
X_31415_ _31415_/A VGND VGND VPWR VPWR _35924_/D sky130_fd_sc_hd__clkbuf_1
X_19137_ _34667_/Q _34603_/Q _34539_/Q _34475_/Q _18886_/X _18887_/X VGND VGND VPWR
+ VPWR _19137_/X sky130_fd_sc_hd__mux4_1
XFILLER_158_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16349_ _33374_/Q _33310_/Q _33246_/Q _33182_/Q _16002_/X _16003_/X VGND VGND VPWR
+ VPWR _16349_/X sky130_fd_sc_hd__mux4_1
XFILLER_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35183_ _35183_/CLK _35183_/D VGND VGND VPWR VPWR _35183_/Q sky130_fd_sc_hd__dfxtp_1
X_32395_ _32907_/CLK _32395_/D VGND VGND VPWR VPWR _32395_/Q sky130_fd_sc_hd__dfxtp_1
X_34134_ _35994_/CLK _34134_/D VGND VGND VPWR VPWR _34134_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19068_ _19064_/X _19067_/X _18759_/X VGND VGND VPWR VPWR _19069_/D sky130_fd_sc_hd__o21ba_1
X_31346_ _31346_/A VGND VGND VPWR VPWR _35891_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18019_ _32141_/Q _32333_/Q _32397_/Q _35917_/Q _17986_/X _17774_/X VGND VGND VPWR
+ VPWR _18019_/X sky130_fd_sc_hd__mux4_1
XFILLER_86_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34065_ _34193_/CLK _34065_/D VGND VGND VPWR VPWR _34065_/Q sky130_fd_sc_hd__dfxtp_1
X_31277_ _27831_/X _35859_/Q _31281_/S VGND VGND VPWR VPWR _31278_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21030_ _20953_/X _21028_/X _21029_/X _20959_/X VGND VGND VPWR VPWR _21030_/X sky130_fd_sc_hd__a22o_1
X_33016_ _36024_/CLK _33016_/D VGND VGND VPWR VPWR _33016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30228_ _30228_/A VGND VGND VPWR VPWR _35361_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30159_ _35329_/Q _29463_/X _30171_/S VGND VGND VPWR VPWR _30160_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34967_ _35673_/CLK _34967_/D VGND VGND VPWR VPWR _34967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22981_ _23083_/S VGND VGND VPWR VPWR _23009_/S sky130_fd_sc_hd__buf_6
XFILLER_95_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24720_ _24720_/A VGND VGND VPWR VPWR _32881_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_216_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33918_ _35711_/CLK _33918_/D VGND VGND VPWR VPWR _33918_/Q sky130_fd_sc_hd__dfxtp_1
X_21932_ _21928_/X _21931_/X _21765_/X VGND VGND VPWR VPWR _21933_/D sky130_fd_sc_hd__o21ba_1
X_34898_ _34964_/CLK _34898_/D VGND VGND VPWR VPWR _34898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24651_ _23070_/X _32849_/Q _24651_/S VGND VGND VPWR VPWR _24652_/A sky130_fd_sc_hd__mux2_1
X_33849_ _33850_/CLK _33849_/D VGND VGND VPWR VPWR _33849_/Q sky130_fd_sc_hd__dfxtp_1
X_21863_ _34423_/Q _36151_/Q _34295_/Q _34231_/Q _21829_/X _21830_/X VGND VGND VPWR
+ VPWR _21863_/X sky130_fd_sc_hd__mux4_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23602_ _22934_/X _32293_/Q _23610_/S VGND VGND VPWR VPWR _23603_/A sky130_fd_sc_hd__mux2_1
X_20814_ _33882_/Q _33818_/Q _33754_/Q _36058_/Q _20712_/X _20713_/X VGND VGND VPWR
+ VPWR _20814_/X sky130_fd_sc_hd__mux4_1
X_27370_ _27502_/S VGND VGND VPWR VPWR _27389_/S sky130_fd_sc_hd__buf_8
XFILLER_242_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24582_ _22968_/X _32816_/Q _24588_/S VGND VGND VPWR VPWR _24583_/A sky130_fd_sc_hd__mux2_1
X_21794_ _34933_/Q _34869_/Q _34805_/Q _34741_/Q _21760_/X _21761_/X VGND VGND VPWR
+ VPWR _21794_/X sky130_fd_sc_hd__mux4_1
XFILLER_196_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26321_ _24951_/X _33607_/Q _26321_/S VGND VGND VPWR VPWR _26322_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23533_ _23533_/A VGND VGND VPWR VPWR _32261_/D sky130_fd_sc_hd__clkbuf_1
X_35519_ _35711_/CLK _35519_/D VGND VGND VPWR VPWR _35519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20745_ _22462_/A VGND VGND VPWR VPWR _20745_/X sky130_fd_sc_hd__buf_4
XFILLER_180_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29040_ _34829_/Q _27205_/X _29048_/S VGND VGND VPWR VPWR _29041_/A sky130_fd_sc_hd__mux2_1
X_26252_ _24849_/X _33574_/Q _26258_/S VGND VGND VPWR VPWR _26253_/A sky130_fd_sc_hd__mux2_1
X_20676_ _20659_/X _20673_/X _20675_/X VGND VGND VPWR VPWR _20706_/C sky130_fd_sc_hd__o21ba_1
X_23464_ _32233_/Q _23463_/X _23485_/S VGND VGND VPWR VPWR _23465_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25203_ _33078_/Q _23396_/X _25217_/S VGND VGND VPWR VPWR _25204_/A sky130_fd_sc_hd__mux2_1
X_22415_ _35655_/Q _35015_/Q _34375_/Q _33735_/Q _22097_/X _22098_/X VGND VGND VPWR
+ VPWR _22415_/X sky130_fd_sc_hd__mux4_1
X_26183_ _26183_/A VGND VGND VPWR VPWR _33541_/D sky130_fd_sc_hd__clkbuf_1
X_23395_ _23395_/A VGND VGND VPWR VPWR _32210_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25134_ _31147_/A _30337_/A VGND VGND VPWR VPWR _25267_/S sky130_fd_sc_hd__nor2_8
X_22346_ _33093_/Q _32069_/Q _35845_/Q _35781_/Q _22031_/X _22032_/X VGND VGND VPWR
+ VPWR _22346_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29942_ _35226_/Q _29342_/X _29952_/S VGND VGND VPWR VPWR _29943_/A sky130_fd_sc_hd__mux2_1
X_22277_ _21956_/X _22275_/X _22276_/X _21959_/X VGND VGND VPWR VPWR _22277_/X sky130_fd_sc_hd__a22o_1
XFILLER_151_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25065_ _25065_/A VGND VGND VPWR VPWR _33013_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21228_ _21228_/A VGND VGND VPWR VPWR _36197_/D sky130_fd_sc_hd__clkbuf_1
X_24016_ _24016_/A VGND VGND VPWR VPWR _32550_/D sky130_fd_sc_hd__clkbuf_1
X_29873_ _29873_/A VGND VGND VPWR VPWR _35193_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28824_ _28824_/A VGND VGND VPWR VPWR _34726_/D sky130_fd_sc_hd__clkbuf_1
X_21159_ _21052_/X _21157_/X _21158_/X _21057_/X VGND VGND VPWR VPWR _21159_/X sky130_fd_sc_hd__a22o_1
XFILLER_24_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28755_ _34695_/Q _27186_/X _28755_/S VGND VGND VPWR VPWR _28756_/A sky130_fd_sc_hd__mux2_1
X_25967_ _24827_/X _33439_/Q _25967_/S VGND VGND VPWR VPWR _25968_/A sky130_fd_sc_hd__mux2_1
XFILLER_246_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27706_ _27704_/X _34218_/Q _27733_/S VGND VGND VPWR VPWR _27707_/A sky130_fd_sc_hd__mux2_1
XTAP_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24918_ _24917_/X _32956_/Q _24921_/S VGND VGND VPWR VPWR _24919_/A sky130_fd_sc_hd__mux2_1
X_28686_ _34662_/Q _27084_/X _28692_/S VGND VGND VPWR VPWR _28687_/A sky130_fd_sc_hd__mux2_1
XTAP_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25898_ _24923_/X _33406_/Q _25916_/S VGND VGND VPWR VPWR _25899_/A sky130_fd_sc_hd__mux2_1
XTAP_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27637_ _34197_/Q _27229_/X _27637_/S VGND VGND VPWR VPWR _27638_/A sky130_fd_sc_hd__mux2_1
XFILLER_218_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24849_ input8/X VGND VGND VPWR VPWR _24849_/X sky130_fd_sc_hd__buf_4
XTAP_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18370_ _33046_/Q _32022_/Q _35798_/Q _35734_/Q _18367_/X _18369_/X VGND VGND VPWR
+ VPWR _18370_/X sky130_fd_sc_hd__mux4_1
XFILLER_215_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27568_ _27637_/S VGND VGND VPWR VPWR _27587_/S sky130_fd_sc_hd__buf_4
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29307_ _29307_/A VGND VGND VPWR VPWR _34955_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_199_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17321_ _16998_/X _17319_/X _17320_/X _17001_/X VGND VGND VPWR VPWR _17321_/X sky130_fd_sc_hd__a22o_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26519_ _26519_/A VGND VGND VPWR VPWR _33699_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27499_ _27499_/A VGND VGND VPWR VPWR _34131_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17252_ _35639_/Q _34999_/Q _34359_/Q _33719_/Q _17144_/X _17145_/X VGND VGND VPWR
+ VPWR _17252_/X sky130_fd_sc_hd__mux4_1
X_29238_ _29238_/A VGND VGND VPWR VPWR _34922_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16203_ _16078_/X _16201_/X _16202_/X _16088_/X VGND VGND VPWR VPWR _16203_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29169_ _34890_/Q _27196_/X _29183_/S VGND VGND VPWR VPWR _29170_/A sky130_fd_sc_hd__mux2_1
XFILLER_179_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17183_ _35701_/Q _32210_/Q _35573_/Q _35509_/Q _16964_/X _16965_/X VGND VGND VPWR
+ VPWR _17183_/X sky130_fd_sc_hd__mux4_1
XFILLER_196_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31200_ _27717_/X _35822_/Q _31210_/S VGND VGND VPWR VPWR _31201_/A sky130_fd_sc_hd__mux2_1
X_16134_ _34391_/Q _36119_/Q _34263_/Q _34199_/Q _16092_/X _16094_/X VGND VGND VPWR
+ VPWR _16134_/X sky130_fd_sc_hd__mux4_1
XFILLER_128_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32180_ _35673_/CLK _32180_/D VGND VGND VPWR VPWR _32180_/Q sky130_fd_sc_hd__dfxtp_1
X_31131_ _35790_/Q input52/X _31137_/S VGND VGND VPWR VPWR _31132_/A sky130_fd_sc_hd__mux2_1
X_16065_ _35414_/Q _35350_/Q _35286_/Q _35222_/Q _16062_/X _16064_/X VGND VGND VPWR
+ VPWR _16065_/X sky130_fd_sc_hd__mux4_1
XFILLER_5_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31062_ _35757_/Q input16/X _31074_/S VGND VGND VPWR VPWR _31063_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30013_ _35260_/Q _29447_/X _30015_/S VGND VGND VPWR VPWR _30014_/A sky130_fd_sc_hd__mux2_1
X_19824_ _19499_/X _19822_/X _19823_/X _19504_/X VGND VGND VPWR VPWR _19824_/X sky130_fd_sc_hd__a22o_1
X_35870_ _35870_/CLK _35870_/D VGND VGND VPWR VPWR _35870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34821_ _36165_/CLK _34821_/D VGND VGND VPWR VPWR _34821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19755_ _33149_/Q _36029_/Q _33021_/Q _32957_/Q _19715_/X _19716_/X VGND VGND VPWR
+ VPWR _19755_/X sky130_fd_sc_hd__mux4_1
X_16967_ _35631_/Q _34991_/Q _34351_/Q _33711_/Q _16791_/X _16792_/X VGND VGND VPWR
+ VPWR _16967_/X sky130_fd_sc_hd__mux4_1
X_18706_ _33055_/Q _32031_/Q _35807_/Q _35743_/Q _18672_/X _18673_/X VGND VGND VPWR
+ VPWR _18706_/X sky130_fd_sc_hd__mux4_1
XFILLER_49_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34752_ _34945_/CLK _34752_/D VGND VGND VPWR VPWR _34752_/Q sky130_fd_sc_hd__dfxtp_1
X_31964_ _34148_/CLK _31964_/D VGND VGND VPWR VPWR _31964_/Q sky130_fd_sc_hd__dfxtp_1
X_16898_ _35693_/Q _32201_/Q _35565_/Q _35501_/Q _16611_/X _16612_/X VGND VGND VPWR
+ VPWR _16898_/X sky130_fd_sc_hd__mux4_1
X_19686_ _32891_/Q _32827_/Q _32763_/Q _32699_/Q _19646_/X _19647_/X VGND VGND VPWR
+ VPWR _19686_/X sky130_fd_sc_hd__mux4_1
XFILLER_65_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33703_ _35559_/CLK _33703_/D VGND VGND VPWR VPWR _33703_/Q sky130_fd_sc_hd__dfxtp_1
X_18637_ _34653_/Q _34589_/Q _34525_/Q _34461_/Q _18533_/X _18534_/X VGND VGND VPWR
+ VPWR _18637_/X sky130_fd_sc_hd__mux4_1
X_30915_ _30915_/A VGND VGND VPWR VPWR _35687_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31895_ _31895_/A VGND VGND VPWR VPWR _36151_/D sky130_fd_sc_hd__clkbuf_1
X_34683_ _34685_/CLK _34683_/D VGND VGND VPWR VPWR _34683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30846_ _35655_/Q input44/X _30846_/S VGND VGND VPWR VPWR _30847_/A sky130_fd_sc_hd__mux2_1
X_33634_ _33827_/CLK _33634_/D VGND VGND VPWR VPWR _33634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18568_ _35163_/Q _35099_/Q _35035_/Q _32155_/Q _18383_/X _18385_/X VGND VGND VPWR
+ VPWR _18568_/X sky130_fd_sc_hd__mux4_1
XFILLER_127_1210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17519_ _17510_/X _17517_/X _17518_/X VGND VGND VPWR VPWR _17520_/D sky130_fd_sc_hd__o21ba_1
XFILLER_36_1126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18499_ _18360_/X _18497_/X _18498_/X _18372_/X VGND VGND VPWR VPWR _18499_/X sky130_fd_sc_hd__a22o_1
X_33565_ _36205_/CLK _33565_/D VGND VGND VPWR VPWR _33565_/Q sky130_fd_sc_hd__dfxtp_1
X_30777_ _35622_/Q input8/X _30783_/S VGND VGND VPWR VPWR _30778_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20530_ _32916_/Q _32852_/Q _32788_/Q _32724_/Q _18284_/X _18287_/X VGND VGND VPWR
+ VPWR _20530_/X sky130_fd_sc_hd__mux4_1
X_35304_ _35685_/CLK _35304_/D VGND VGND VPWR VPWR _35304_/Q sky130_fd_sc_hd__dfxtp_1
X_32516_ _35973_/CLK _32516_/D VGND VGND VPWR VPWR _32516_/Q sky130_fd_sc_hd__dfxtp_1
X_33496_ _36057_/CLK _33496_/D VGND VGND VPWR VPWR _33496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20461_ _20205_/X _20459_/X _20460_/X _20210_/X VGND VGND VPWR VPWR _20461_/X sky130_fd_sc_hd__a22o_1
X_32447_ _36075_/CLK _32447_/D VGND VGND VPWR VPWR _32447_/Q sky130_fd_sc_hd__dfxtp_1
X_35235_ _35814_/CLK _35235_/D VGND VGND VPWR VPWR _35235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22200_ _32129_/Q _32321_/Q _32385_/Q _35905_/Q _21880_/X _22021_/X VGND VGND VPWR
+ VPWR _22200_/X sky130_fd_sc_hd__mux4_1
XFILLER_174_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23180_ _23018_/X _32128_/Q _23194_/S VGND VGND VPWR VPWR _23181_/A sky130_fd_sc_hd__mux2_1
XFILLER_238_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20392_ _20159_/X _20390_/X _20391_/X _20162_/X VGND VGND VPWR VPWR _20392_/X sky130_fd_sc_hd__a22o_1
X_35166_ _35609_/CLK _35166_/D VGND VGND VPWR VPWR _35166_/Q sky130_fd_sc_hd__dfxtp_1
X_32378_ _32890_/CLK _32378_/D VGND VGND VPWR VPWR _32378_/Q sky130_fd_sc_hd__dfxtp_1
X_22131_ _22012_/X _22129_/X _22130_/X _22018_/X VGND VGND VPWR VPWR _22131_/X sky130_fd_sc_hd__a22o_1
X_34117_ _34945_/CLK _34117_/D VGND VGND VPWR VPWR _34117_/Q sky130_fd_sc_hd__dfxtp_1
X_31329_ _27708_/X _35883_/Q _31345_/S VGND VGND VPWR VPWR _31330_/A sky130_fd_sc_hd__mux2_1
XFILLER_238_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35097_ _35799_/CLK _35097_/D VGND VGND VPWR VPWR _35097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput220 _32417_/Q VGND VGND VPWR VPWR D3[11] sky130_fd_sc_hd__buf_2
Xoutput231 _32427_/Q VGND VGND VPWR VPWR D3[21] sky130_fd_sc_hd__buf_2
Xoutput242 _32437_/Q VGND VGND VPWR VPWR D3[31] sky130_fd_sc_hd__buf_2
XTAP_6608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput253 _32447_/Q VGND VGND VPWR VPWR D3[41] sky130_fd_sc_hd__buf_2
X_22062_ _35645_/Q _35005_/Q _34365_/Q _33725_/Q _21744_/X _21745_/X VGND VGND VPWR
+ VPWR _22062_/X sky130_fd_sc_hd__mux4_1
XTAP_6619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34048_ _34942_/CLK _34048_/D VGND VGND VPWR VPWR _34048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput264 _32457_/Q VGND VGND VPWR VPWR D3[51] sky130_fd_sc_hd__buf_2
XFILLER_102_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput275 _32467_/Q VGND VGND VPWR VPWR D3[61] sky130_fd_sc_hd__buf_2
Xclkbuf_6_3__f_CLK clkbuf_5_1_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_3__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_82_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21013_ _34911_/Q _34847_/Q _34783_/Q _34719_/Q _20696_/X _20698_/X VGND VGND VPWR
+ VPWR _21013_/X sky130_fd_sc_hd__mux4_1
XFILLER_87_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26870_ _33864_/Q _23453_/X _26888_/S VGND VGND VPWR VPWR _26871_/A sky130_fd_sc_hd__mux2_1
XTAP_5918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25821_ _25821_/A VGND VGND VPWR VPWR _33369_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35999_ _35999_/CLK _35999_/D VGND VGND VPWR VPWR _35999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28540_ _27677_/X _34593_/Q _28556_/S VGND VGND VPWR VPWR _28541_/A sky130_fd_sc_hd__mux2_1
X_25752_ _24908_/X _33337_/Q _25760_/S VGND VGND VPWR VPWR _25753_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22964_ _22964_/A VGND VGND VPWR VPWR _32046_/D sky130_fd_sc_hd__clkbuf_1
X_24703_ _24703_/A VGND VGND VPWR VPWR _32873_/D sky130_fd_sc_hd__clkbuf_1
X_28471_ _28471_/A VGND VGND VPWR VPWR _34560_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21915_ _21667_/X _21913_/X _21914_/X _21671_/X VGND VGND VPWR VPWR _21915_/X sky130_fd_sc_hd__a22o_1
XFILLER_243_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25683_ _24806_/X _33304_/Q _25697_/S VGND VGND VPWR VPWR _25684_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22895_ _22894_/X _32024_/Q _22916_/S VGND VGND VPWR VPWR _22896_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27422_ _27422_/A VGND VGND VPWR VPWR _34094_/D sky130_fd_sc_hd__clkbuf_1
X_24634_ _24634_/A VGND VGND VPWR VPWR _32840_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21846_ _21659_/X _21844_/X _21845_/X _21665_/X VGND VGND VPWR VPWR _21846_/X sky130_fd_sc_hd__a22o_1
XFILLER_24_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27353_ _34062_/Q _27208_/X _27359_/S VGND VGND VPWR VPWR _27354_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24565_ _22943_/X _32808_/Q _24567_/S VGND VGND VPWR VPWR _24566_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21777_ _33141_/Q _36021_/Q _33013_/Q _32949_/Q _21662_/X _21663_/X VGND VGND VPWR
+ VPWR _21777_/X sky130_fd_sc_hd__mux4_1
X_26304_ _26304_/A VGND VGND VPWR VPWR _33598_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23516_ _23516_/A VGND VGND VPWR VPWR _32253_/D sky130_fd_sc_hd__clkbuf_1
X_20728_ _33047_/Q _32023_/Q _35799_/Q _35735_/Q _20667_/X _20669_/X VGND VGND VPWR
+ VPWR _20728_/X sky130_fd_sc_hd__mux4_1
X_27284_ _34029_/Q _27106_/X _27296_/S VGND VGND VPWR VPWR _27285_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_929 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24496_ _24496_/A VGND VGND VPWR VPWR _32775_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29023_ _34821_/Q _27180_/X _29027_/S VGND VGND VPWR VPWR _29024_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26235_ _24824_/X _33566_/Q _26237_/S VGND VGND VPWR VPWR _26236_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23447_ input43/X VGND VGND VPWR VPWR _23447_/X sky130_fd_sc_hd__buf_6
X_20659_ _20648_/X _20651_/X _20656_/X _20658_/X VGND VGND VPWR VPWR _20659_/X sky130_fd_sc_hd__a22o_1
XFILLER_221_1275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_804 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26166_ _26166_/A VGND VGND VPWR VPWR _33533_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23378_ _23378_/A VGND VGND VPWR VPWR _32204_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25117_ _25117_/A VGND VGND VPWR VPWR _33038_/D sky130_fd_sc_hd__clkbuf_1
X_22329_ _33413_/Q _33349_/Q _33285_/Q _33221_/Q _22080_/X _22081_/X VGND VGND VPWR
+ VPWR _22329_/X sky130_fd_sc_hd__mux4_1
XFILLER_152_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26097_ _26097_/A VGND VGND VPWR VPWR _33500_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29925_ _29925_/A VGND VGND VPWR VPWR _35218_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25048_ _25048_/A VGND VGND VPWR VPWR _33005_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_870 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17870_ _17864_/X _17865_/X _17868_/X _17869_/X VGND VGND VPWR VPWR _17870_/X sky130_fd_sc_hd__a22o_1
X_29856_ _29856_/A VGND VGND VPWR VPWR _35185_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_238_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28807_ _28807_/A VGND VGND VPWR VPWR _34718_/D sky130_fd_sc_hd__clkbuf_1
X_16821_ _16500_/X _16819_/X _16820_/X _16503_/X VGND VGND VPWR VPWR _16821_/X sky130_fd_sc_hd__a22o_1
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29787_ _35153_/Q _29512_/X _29787_/S VGND VGND VPWR VPWR _29788_/A sky130_fd_sc_hd__mux2_1
X_26999_ _26999_/A VGND VGND VPWR VPWR _33925_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19540_ _33399_/Q _33335_/Q _33271_/Q _33207_/Q _19427_/X _19428_/X VGND VGND VPWR
+ VPWR _19540_/X sky130_fd_sc_hd__mux4_1
X_16752_ _32873_/Q _32809_/Q _32745_/Q _32681_/Q _16640_/X _16641_/X VGND VGND VPWR
+ VPWR _16752_/X sky130_fd_sc_hd__mux4_1
X_28738_ _28738_/A VGND VGND VPWR VPWR _34686_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28669_ _34654_/Q _27059_/X _28671_/S VGND VGND VPWR VPWR _28670_/A sky130_fd_sc_hd__mux2_1
X_19471_ _19146_/X _19469_/X _19470_/X _19151_/X VGND VGND VPWR VPWR _19471_/X sky130_fd_sc_hd__a22o_1
X_16683_ _35687_/Q _32194_/Q _35559_/Q _35495_/Q _16611_/X _16612_/X VGND VGND VPWR
+ VPWR _16683_/X sky130_fd_sc_hd__mux4_1
XFILLER_34_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_1006 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30700_ _30700_/A VGND VGND VPWR VPWR _35585_/D sky130_fd_sc_hd__clkbuf_1
X_18422_ _18330_/X _18420_/X _18421_/X _18341_/X VGND VGND VPWR VPWR _18422_/X sky130_fd_sc_hd__a22o_1
XFILLER_46_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31680_ _27828_/X _36050_/Q _31686_/S VGND VGND VPWR VPWR _31681_/A sky130_fd_sc_hd__mux2_1
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18353_ _20298_/A VGND VGND VPWR VPWR _18353_/X sky130_fd_sc_hd__buf_6
XFILLER_61_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30631_ _30631_/A VGND VGND VPWR VPWR _35552_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_203_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_863 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_230_CLK clkbuf_6_55__f_CLK/X VGND VGND VPWR VPWR _34187_/CLK sky130_fd_sc_hd__clkbuf_16
X_17304_ _34169_/Q _34105_/Q _34041_/Q _33977_/Q _17093_/X _17094_/X VGND VGND VPWR
+ VPWR _17304_/X sky130_fd_sc_hd__mux4_1
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33350_ _33415_/CLK _33350_/D VGND VGND VPWR VPWR _33350_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30562_ _35520_/Q _29460_/X _30576_/S VGND VGND VPWR VPWR _30563_/A sky130_fd_sc_hd__mux2_1
X_18284_ _20206_/A VGND VGND VPWR VPWR _18284_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_187_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32301_ _35951_/CLK _32301_/D VGND VGND VPWR VPWR _32301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17235_ _17235_/A _17235_/B _17235_/C _17235_/D VGND VGND VPWR VPWR _17236_/A sky130_fd_sc_hd__or4_4
XFILLER_204_1462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33281_ _33924_/CLK _33281_/D VGND VGND VPWR VPWR _33281_/Q sky130_fd_sc_hd__dfxtp_1
X_30493_ _30493_/A VGND VGND VPWR VPWR _35487_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32232_ _35658_/CLK _32232_/D VGND VGND VPWR VPWR _32232_/Q sky130_fd_sc_hd__dfxtp_1
X_35020_ _35661_/CLK _35020_/D VGND VGND VPWR VPWR _35020_/Q sky130_fd_sc_hd__dfxtp_1
X_17166_ _17157_/X _17164_/X _17165_/X VGND VGND VPWR VPWR _17167_/D sky130_fd_sc_hd__o21ba_1
XFILLER_128_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16117_ _32599_/Q _32535_/Q _32471_/Q _35927_/Q _17866_/A _17717_/A VGND VGND VPWR
+ VPWR _16117_/X sky130_fd_sc_hd__mux4_1
XFILLER_157_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32163_ _36210_/CLK _32163_/D VGND VGND VPWR VPWR _32163_/Q sky130_fd_sc_hd__dfxtp_1
X_17097_ _33395_/Q _33331_/Q _33267_/Q _33203_/Q _16774_/X _16775_/X VGND VGND VPWR
+ VPWR _17097_/X sky130_fd_sc_hd__mux4_1
XFILLER_143_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_1460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31114_ _35782_/Q input43/X _31116_/S VGND VGND VPWR VPWR _31115_/A sky130_fd_sc_hd__mux2_1
X_16048_ _17859_/A VGND VGND VPWR VPWR _16048_/X sky130_fd_sc_hd__clkbuf_4
X_32094_ _32869_/CLK _32094_/D VGND VGND VPWR VPWR _32094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_297_CLK clkbuf_6_56__f_CLK/X VGND VGND VPWR VPWR _36034_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_83_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35922_ _35922_/CLK _35922_/D VGND VGND VPWR VPWR _35922_/Q sky130_fd_sc_hd__dfxtp_1
X_31045_ _35749_/Q input7/X _31053_/S VGND VGND VPWR VPWR _31046_/A sky130_fd_sc_hd__mux2_1
X_19807_ _34686_/Q _34622_/Q _34558_/Q _34494_/Q _19592_/X _19593_/X VGND VGND VPWR
+ VPWR _19807_/X sky130_fd_sc_hd__mux4_1
XFILLER_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35853_ _35853_/CLK _35853_/D VGND VGND VPWR VPWR _35853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17999_ _17999_/A VGND VGND VPWR VPWR _17999_/X sky130_fd_sc_hd__buf_4
X_34804_ _35828_/CLK _34804_/D VGND VGND VPWR VPWR _34804_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19738_ _19453_/X _19736_/X _19737_/X _19456_/X VGND VGND VPWR VPWR _19738_/X sky130_fd_sc_hd__a22o_1
XFILLER_244_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35784_ _35785_/CLK _35784_/D VGND VGND VPWR VPWR _35784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32996_ _34593_/CLK _32996_/D VGND VGND VPWR VPWR _32996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34735_ _34926_/CLK _34735_/D VGND VGND VPWR VPWR _34735_/Q sky130_fd_sc_hd__dfxtp_1
X_31947_ _31947_/A VGND VGND VPWR VPWR _36176_/D sky130_fd_sc_hd__clkbuf_1
X_19669_ _19458_/X _19667_/X _19668_/X _19463_/X VGND VGND VPWR VPWR _19669_/X sky130_fd_sc_hd__a22o_1
XFILLER_64_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21700_ _21696_/X _21699_/X _21379_/X VGND VGND VPWR VPWR _21722_/A sky130_fd_sc_hd__o21ba_1
X_22680_ _32911_/Q _32847_/Q _32783_/Q _32719_/Q _20584_/X _20587_/X VGND VGND VPWR
+ VPWR _22680_/X sky130_fd_sc_hd__mux4_1
XFILLER_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34666_ _35564_/CLK _34666_/D VGND VGND VPWR VPWR _34666_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31878_ _31878_/A VGND VGND VPWR VPWR _36143_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33617_ _34441_/CLK _33617_/D VGND VGND VPWR VPWR _33617_/Q sky130_fd_sc_hd__dfxtp_1
X_21631_ _21306_/X _21629_/X _21630_/X _21312_/X VGND VGND VPWR VPWR _21631_/X sky130_fd_sc_hd__a22o_1
X_30829_ _30829_/A VGND VGND VPWR VPWR _35646_/D sky130_fd_sc_hd__clkbuf_1
X_34597_ _36136_/CLK _34597_/D VGND VGND VPWR VPWR _34597_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_221_CLK clkbuf_6_53__f_CLK/X VGND VGND VPWR VPWR _34956_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_240_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24350_ _23024_/X _32706_/Q _24360_/S VGND VGND VPWR VPWR _24351_/A sky130_fd_sc_hd__mux2_1
X_33548_ _34188_/CLK _33548_/D VGND VGND VPWR VPWR _33548_/Q sky130_fd_sc_hd__dfxtp_1
X_21562_ _21314_/X _21560_/X _21561_/X _21318_/X VGND VGND VPWR VPWR _21562_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23301_ _23301_/A VGND VGND VPWR VPWR _32172_/D sky130_fd_sc_hd__clkbuf_1
X_20513_ _34451_/Q _36179_/Q _34323_/Q _34259_/Q _20235_/X _20236_/X VGND VGND VPWR
+ VPWR _20513_/X sky130_fd_sc_hd__mux4_1
X_24281_ _22922_/X _32673_/Q _24297_/S VGND VGND VPWR VPWR _24282_/A sky130_fd_sc_hd__mux2_1
X_21493_ _21306_/X _21491_/X _21492_/X _21312_/X VGND VGND VPWR VPWR _21493_/X sky130_fd_sc_hd__a22o_1
X_33479_ _34185_/CLK _33479_/D VGND VGND VPWR VPWR _33479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26020_ _24905_/X _33464_/Q _26030_/S VGND VGND VPWR VPWR _26021_/A sky130_fd_sc_hd__mux2_1
X_23232_ _32150_/Q _23225_/X _23259_/S VGND VGND VPWR VPWR _23233_/A sky130_fd_sc_hd__mux2_1
X_35218_ _36114_/CLK _35218_/D VGND VGND VPWR VPWR _35218_/Q sky130_fd_sc_hd__dfxtp_1
X_20444_ _35665_/Q _35025_/Q _34385_/Q _33745_/Q _20150_/X _20151_/X VGND VGND VPWR
+ VPWR _20444_/X sky130_fd_sc_hd__mux4_1
XFILLER_153_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36198_ _36207_/CLK _36198_/D VGND VGND VPWR VPWR _36198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_1295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20375_ _20371_/X _20374_/X _20138_/X VGND VGND VPWR VPWR _20397_/A sky130_fd_sc_hd__o21ba_2
X_35149_ _35663_/CLK _35149_/D VGND VGND VPWR VPWR _35149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23163_ _22993_/X _32120_/Q _23173_/S VGND VGND VPWR VPWR _23164_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22114_ _22467_/A VGND VGND VPWR VPWR _22114_/X sky130_fd_sc_hd__clkbuf_4
XTAP_7139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27971_ _27834_/X _34324_/Q _27973_/S VGND VGND VPWR VPWR _27972_/A sky130_fd_sc_hd__mux2_1
X_23094_ _22891_/X _32087_/Q _23110_/S VGND VGND VPWR VPWR _23095_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_288_CLK clkbuf_6_58__f_CLK/X VGND VGND VPWR VPWR _36031_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_6438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22045_ _33661_/Q _33597_/Q _33533_/Q _33469_/Q _21800_/X _21801_/X VGND VGND VPWR
+ VPWR _22045_/X sky130_fd_sc_hd__mux4_1
X_26922_ _26922_/A VGND VGND VPWR VPWR _33888_/D sky130_fd_sc_hd__clkbuf_1
X_29710_ _35116_/Q _29398_/X _29724_/S VGND VGND VPWR VPWR _29711_/A sky130_fd_sc_hd__mux2_1
XTAP_6449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29641_ _29641_/A VGND VGND VPWR VPWR _35083_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26853_ _33856_/Q _23429_/X _26867_/S VGND VGND VPWR VPWR _26854_/A sky130_fd_sc_hd__mux2_1
XTAP_5759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_810 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25804_ _24985_/X _33362_/Q _25810_/S VGND VGND VPWR VPWR _25805_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29572_ _29572_/A VGND VGND VPWR VPWR _35050_/D sky130_fd_sc_hd__clkbuf_1
X_26784_ _26784_/A VGND VGND VPWR VPWR _33823_/D sky130_fd_sc_hd__clkbuf_1
X_23996_ _22909_/X _32541_/Q _24000_/S VGND VGND VPWR VPWR _23997_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28523_ _27652_/X _34585_/Q _28535_/S VGND VGND VPWR VPWR _28524_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25735_ _24883_/X _33329_/Q _25739_/S VGND VGND VPWR VPWR _25736_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22947_ _22946_/X _32041_/Q _22947_/S VGND VGND VPWR VPWR _22948_/A sky130_fd_sc_hd__mux2_1
XFILLER_244_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_460_CLK clkbuf_6_9__f_CLK/X VGND VGND VPWR VPWR _35433_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_83_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_616 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28454_ _28454_/A VGND VGND VPWR VPWR _34552_/D sky130_fd_sc_hd__clkbuf_1
X_25666_ _25666_/A VGND VGND VPWR VPWR _33296_/D sky130_fd_sc_hd__clkbuf_1
X_22878_ _22878_/A VGND VGND VPWR VPWR _36245_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27405_ _27405_/A VGND VGND VPWR VPWR _34086_/D sky130_fd_sc_hd__clkbuf_1
X_24617_ _24617_/A VGND VGND VPWR VPWR _32832_/D sky130_fd_sc_hd__clkbuf_1
X_28385_ _28385_/A VGND VGND VPWR VPWR _34519_/D sky130_fd_sc_hd__clkbuf_1
X_21829_ _22535_/A VGND VGND VPWR VPWR _21829_/X sky130_fd_sc_hd__buf_8
X_25597_ _25597_/A VGND VGND VPWR VPWR _33263_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_227_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_212_CLK clkbuf_6_52__f_CLK/X VGND VGND VPWR VPWR _35724_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_145_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27336_ _34054_/Q _27183_/X _27338_/S VGND VGND VPWR VPWR _27337_/A sky130_fd_sc_hd__mux2_1
XFILLER_200_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24548_ _24659_/S VGND VGND VPWR VPWR _24567_/S sky130_fd_sc_hd__buf_4
XFILLER_12_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27267_ _34021_/Q _27081_/X _27275_/S VGND VGND VPWR VPWR _27268_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24479_ _23015_/X _32767_/Q _24495_/S VGND VGND VPWR VPWR _24480_/A sky130_fd_sc_hd__mux2_1
XFILLER_221_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17020_ _33649_/Q _33585_/Q _33521_/Q _33457_/Q _16847_/X _16848_/X VGND VGND VPWR
+ VPWR _17020_/X sky130_fd_sc_hd__mux4_1
X_29006_ _34813_/Q _27155_/X _29006_/S VGND VGND VPWR VPWR _29007_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26218_ _26350_/S VGND VGND VPWR VPWR _26237_/S sky130_fd_sc_hd__buf_6
XFILLER_32_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27198_ _27198_/A VGND VGND VPWR VPWR _33994_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_5_15_0_CLK clkbuf_5_9_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_15_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_50_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26149_ _24896_/X _33525_/Q _26165_/S VGND VGND VPWR VPWR _26150_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_964 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18971_ _20150_/A VGND VGND VPWR VPWR _18971_/X sky130_fd_sc_hd__buf_4
XFILLER_234_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_279_CLK clkbuf_6_59__f_CLK/X VGND VGND VPWR VPWR _33921_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29908_ _35210_/Q _29491_/X _29922_/S VGND VGND VPWR VPWR _29909_/A sky130_fd_sc_hd__mux2_1
X_17922_ _32906_/Q _32842_/Q _32778_/Q _32714_/Q _17699_/X _17700_/X VGND VGND VPWR
+ VPWR _17922_/X sky130_fd_sc_hd__mux4_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17853_ _17704_/X _17849_/X _17852_/X _17707_/X VGND VGND VPWR VPWR _17853_/X sky130_fd_sc_hd__a22o_1
X_29839_ _29839_/A VGND VGND VPWR VPWR _35177_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16804_ _16800_/X _16801_/X _16802_/X _16803_/X VGND VGND VPWR VPWR _16804_/X sky130_fd_sc_hd__a22o_1
X_32850_ _32914_/CLK _32850_/D VGND VGND VPWR VPWR _32850_/Q sky130_fd_sc_hd__dfxtp_1
X_17784_ _17935_/A VGND VGND VPWR VPWR _17784_/X sky130_fd_sc_hd__buf_6
XFILLER_219_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31801_ _36107_/Q input49/X _31813_/S VGND VGND VPWR VPWR _31802_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19523_ _33078_/Q _32054_/Q _35830_/Q _35766_/Q _19378_/X _19379_/X VGND VGND VPWR
+ VPWR _19523_/X sky130_fd_sc_hd__mux4_1
XFILLER_47_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16735_ _16452_/X _16733_/X _16734_/X _16457_/X VGND VGND VPWR VPWR _16735_/X sky130_fd_sc_hd__a22o_1
X_32781_ _32909_/CLK _32781_/D VGND VGND VPWR VPWR _32781_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_451_CLK clkbuf_6_14__f_CLK/X VGND VGND VPWR VPWR _35822_/CLK sky130_fd_sc_hd__clkbuf_16
X_34520_ _34904_/CLK _34520_/D VGND VGND VPWR VPWR _34520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_235_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31732_ _36074_/Q input13/X _31750_/S VGND VGND VPWR VPWR _31733_/A sky130_fd_sc_hd__mux2_1
X_16666_ _16666_/A VGND VGND VPWR VPWR _31974_/D sky130_fd_sc_hd__clkbuf_1
X_19454_ _34676_/Q _34612_/Q _34548_/Q _34484_/Q _19239_/X _19240_/X VGND VGND VPWR
+ VPWR _19454_/X sky130_fd_sc_hd__mux4_1
XFILLER_35_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18405_ _18389_/X _18402_/X _18404_/X VGND VGND VPWR VPWR _18406_/D sky130_fd_sc_hd__o21ba_1
XFILLER_222_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34451_ _34963_/CLK _34451_/D VGND VGND VPWR VPWR _34451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31663_ _31663_/A VGND VGND VPWR VPWR _36041_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16597_ _33637_/Q _33573_/Q _33509_/Q _33445_/Q _16494_/X _16495_/X VGND VGND VPWR
+ VPWR _16597_/X sky130_fd_sc_hd__mux4_1
X_19385_ _19100_/X _19383_/X _19384_/X _19103_/X VGND VGND VPWR VPWR _19385_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_203_CLK clkbuf_6_51__f_CLK/X VGND VGND VPWR VPWR _35722_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33402_ _33914_/CLK _33402_/D VGND VGND VPWR VPWR _33402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30614_ _30614_/A VGND VGND VPWR VPWR _35544_/D sky130_fd_sc_hd__clkbuf_1
X_18336_ _18361_/A VGND VGND VPWR VPWR _20133_/A sky130_fd_sc_hd__buf_12
XFILLER_194_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34382_ _35664_/CLK _34382_/D VGND VGND VPWR VPWR _34382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31594_ _27701_/X _36009_/Q _31594_/S VGND VGND VPWR VPWR _31595_/A sky130_fd_sc_hd__mux2_1
X_36121_ _36121_/CLK _36121_/D VGND VGND VPWR VPWR _36121_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18267_ _33109_/Q _32085_/Q _35861_/Q _35797_/Q _16079_/X _16080_/X VGND VGND VPWR
+ VPWR _18267_/X sky130_fd_sc_hd__mux4_1
X_33333_ _34100_/CLK _33333_/D VGND VGND VPWR VPWR _33333_/Q sky130_fd_sc_hd__dfxtp_1
X_30545_ _35512_/Q _29435_/X _30555_/S VGND VGND VPWR VPWR _30546_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36052_ _36052_/CLK _36052_/D VGND VGND VPWR VPWR _36052_/Q sky130_fd_sc_hd__dfxtp_1
X_17218_ _17214_/X _17217_/X _17140_/X _17141_/X VGND VGND VPWR VPWR _17235_/B sky130_fd_sc_hd__o211a_1
XFILLER_239_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30476_ _35479_/Q _29333_/X _30492_/S VGND VGND VPWR VPWR _30477_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18198_ _17153_/A _18196_/X _18197_/X _17156_/A VGND VGND VPWR VPWR _18198_/X sky130_fd_sc_hd__a22o_1
X_33264_ _33904_/CLK _33264_/D VGND VGND VPWR VPWR _33264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35003_ _35644_/CLK _35003_/D VGND VGND VPWR VPWR _35003_/Q sky130_fd_sc_hd__dfxtp_1
X_17149_ _33076_/Q _32052_/Q _35828_/Q _35764_/Q _17078_/X _17079_/X VGND VGND VPWR
+ VPWR _17149_/X sky130_fd_sc_hd__mux4_1
X_32215_ _35581_/CLK _32215_/D VGND VGND VPWR VPWR _32215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33195_ _36075_/CLK _33195_/D VGND VGND VPWR VPWR _33195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_6_16__f_CLK clkbuf_5_8_0_CLK/X VGND VGND VPWR VPWR clkbuf_leaf_96_CLK/A sky130_fd_sc_hd__clkbuf_16
XFILLER_6_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20160_ _34696_/Q _34632_/Q _34568_/Q _34504_/Q _19945_/X _19946_/X VGND VGND VPWR
+ VPWR _20160_/X sky130_fd_sc_hd__mux4_1
XFILLER_196_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32146_ _35922_/CLK _32146_/D VGND VGND VPWR VPWR _32146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20091_ _19806_/X _20089_/X _20090_/X _19809_/X VGND VGND VPWR VPWR _20091_/X sky130_fd_sc_hd__a22o_1
XFILLER_157_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32077_ _35852_/CLK _32077_/D VGND VGND VPWR VPWR _32077_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31028_ _35741_/Q input62/X _31032_/S VGND VGND VPWR VPWR _31029_/A sky130_fd_sc_hd__mux2_1
X_35905_ _35969_/CLK _35905_/D VGND VGND VPWR VPWR _35905_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_245_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_218_719 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23850_ _22894_/X _32472_/Q _23864_/S VGND VGND VPWR VPWR _23851_/A sky130_fd_sc_hd__mux2_1
XTAP_3609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35836_ _36029_/CLK _35836_/D VGND VGND VPWR VPWR _35836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22801_ _21758_/A _22799_/X _22800_/X _21763_/A VGND VGND VPWR VPWR _22801_/X sky130_fd_sc_hd__a22o_1
XFILLER_242_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35767_ _35830_/CLK _35767_/D VGND VGND VPWR VPWR _35767_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23781_ _23781_/A VGND VGND VPWR VPWR _32376_/D sky130_fd_sc_hd__clkbuf_1
X_32979_ _35859_/CLK _32979_/D VGND VGND VPWR VPWR _32979_/Q sky130_fd_sc_hd__dfxtp_1
X_20993_ _20747_/X _20991_/X _20992_/X _20750_/X VGND VGND VPWR VPWR _20993_/X sky130_fd_sc_hd__a22o_1
XFILLER_53_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25520_ _24964_/X _33227_/Q _25532_/S VGND VGND VPWR VPWR _25521_/A sky130_fd_sc_hd__mux2_1
XFILLER_214_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_442_CLK clkbuf_6_37__f_CLK/X VGND VGND VPWR VPWR _35952_/CLK sky130_fd_sc_hd__clkbuf_16
X_34718_ _36245_/CLK _34718_/D VGND VGND VPWR VPWR _34718_/Q sky130_fd_sc_hd__dfxtp_1
X_22732_ _33425_/Q _33361_/Q _33297_/Q _33233_/Q _22433_/X _22434_/X VGND VGND VPWR
+ VPWR _22732_/X sky130_fd_sc_hd__mux4_2
XFILLER_26_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35698_ _35698_/CLK _35698_/D VGND VGND VPWR VPWR _35698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25451_ _24861_/X _33194_/Q _25469_/S VGND VGND VPWR VPWR _25452_/A sky130_fd_sc_hd__mux2_1
X_34649_ _34903_/CLK _34649_/D VGND VGND VPWR VPWR _34649_/Q sky130_fd_sc_hd__dfxtp_1
X_22663_ _34446_/Q _36174_/Q _34318_/Q _34254_/Q _22535_/X _22536_/X VGND VGND VPWR
+ VPWR _22663_/X sky130_fd_sc_hd__mux4_1
XFILLER_179_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24402_ _24402_/A VGND VGND VPWR VPWR _32730_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21614_ _34416_/Q _36144_/Q _34288_/Q _34224_/Q _21476_/X _21477_/X VGND VGND VPWR
+ VPWR _21614_/X sky130_fd_sc_hd__mux4_1
X_28170_ _27729_/X _34418_/Q _28172_/S VGND VGND VPWR VPWR _28171_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_1422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25382_ _25382_/A VGND VGND VPWR VPWR _33162_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22594_ _35468_/Q _35404_/Q _35340_/Q _35276_/Q _22560_/X _22561_/X VGND VGND VPWR
+ VPWR _22594_/X sky130_fd_sc_hd__mux4_1
XFILLER_146_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27121_ input21/X VGND VGND VPWR VPWR _27121_/X sky130_fd_sc_hd__buf_2
X_24333_ _22999_/X _32698_/Q _24339_/S VGND VGND VPWR VPWR _24334_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21545_ _34926_/Q _34862_/Q _34798_/Q _34734_/Q _21407_/X _21408_/X VGND VGND VPWR
+ VPWR _21545_/X sky130_fd_sc_hd__mux4_1
XFILLER_224_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27052_ _27052_/A VGND VGND VPWR VPWR _33947_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24264_ _22897_/X _32665_/Q _24276_/S VGND VGND VPWR VPWR _24265_/A sky130_fd_sc_hd__mux2_1
X_21476_ _22316_/A VGND VGND VPWR VPWR _21476_/X sky130_fd_sc_hd__buf_4
XFILLER_181_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26003_ _24880_/X _33456_/Q _26009_/S VGND VGND VPWR VPWR _26004_/A sky130_fd_sc_hd__mux2_1
X_23215_ _23070_/X _32145_/Q _23215_/S VGND VGND VPWR VPWR _23216_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20427_ _20427_/A _20427_/B _20427_/C _20427_/D VGND VGND VPWR VPWR _20428_/A sky130_fd_sc_hd__or4_1
XFILLER_4_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24195_ _32634_/Q _23408_/X _24201_/S VGND VGND VPWR VPWR _24196_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23146_ _22968_/X _32112_/Q _23152_/S VGND VGND VPWR VPWR _23147_/A sky130_fd_sc_hd__mux2_1
X_20358_ _18301_/X _20356_/X _20357_/X _18307_/X VGND VGND VPWR VPWR _20358_/X sky130_fd_sc_hd__a22o_1
XTAP_6202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27954_ _27954_/A VGND VGND VPWR VPWR _34315_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23077_ _23076_/X _32083_/Q _23083_/S VGND VGND VPWR VPWR _23078_/A sky130_fd_sc_hd__mux2_1
X_20289_ _20073_/X _20287_/X _20288_/X _20077_/X VGND VGND VPWR VPWR _20289_/X sky130_fd_sc_hd__a22o_1
XFILLER_121_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_1163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26905_ _26905_/A VGND VGND VPWR VPWR _33880_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22028_ _35644_/Q _35004_/Q _34364_/Q _33724_/Q _21744_/X _21745_/X VGND VGND VPWR
+ VPWR _22028_/X sky130_fd_sc_hd__mux4_1
XTAP_6279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27885_ _27885_/A VGND VGND VPWR VPWR _34282_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29624_ _29624_/A VGND VGND VPWR VPWR _35075_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26836_ _33848_/Q _23402_/X _26846_/S VGND VGND VPWR VPWR _26837_/A sky130_fd_sc_hd__mux2_1
XTAP_5589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26767_ _33815_/Q _23234_/X _26783_/S VGND VGND VPWR VPWR _26768_/A sky130_fd_sc_hd__mux2_1
XTAP_4888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29555_ _29555_/A VGND VGND VPWR VPWR _35042_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23979_ _27232_/B _25132_/A _28786_/A VGND VGND VPWR VPWR _31553_/A sky130_fd_sc_hd__nor3_4
XFILLER_56_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_433_CLK clkbuf_6_36__f_CLK/X VGND VGND VPWR VPWR _36147_/CLK sky130_fd_sc_hd__clkbuf_16
X_16520_ _34658_/Q _34594_/Q _34530_/Q _34466_/Q _16233_/X _16234_/X VGND VGND VPWR
+ VPWR _16520_/X sky130_fd_sc_hd__mux4_1
X_28506_ _28506_/A VGND VGND VPWR VPWR _34577_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_217_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25718_ _24858_/X _33321_/Q _25718_/S VGND VGND VPWR VPWR _25719_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29486_ _35016_/Q _29484_/X _29513_/S VGND VGND VPWR VPWR _29487_/A sky130_fd_sc_hd__mux2_1
XFILLER_189_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26698_ _26698_/A VGND VGND VPWR VPWR _33782_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16451_ _16447_/X _16448_/X _16449_/X _16450_/X VGND VGND VPWR VPWR _16451_/X sky130_fd_sc_hd__a22o_1
X_25649_ _24954_/X _33288_/Q _25667_/S VGND VGND VPWR VPWR _25650_/A sky130_fd_sc_hd__mux2_1
X_28437_ _28437_/A VGND VGND VPWR VPWR _34544_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19170_ _33068_/Q _32044_/Q _35820_/Q _35756_/Q _19025_/X _19026_/X VGND VGND VPWR
+ VPWR _19170_/X sky130_fd_sc_hd__mux4_1
X_16382_ _16091_/X _16380_/X _16381_/X _16101_/X VGND VGND VPWR VPWR _16382_/X sky130_fd_sc_hd__a22o_1
X_28368_ _27822_/X _34512_/Q _28370_/S VGND VGND VPWR VPWR _28369_/A sky130_fd_sc_hd__mux2_1
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18121_ _35216_/Q _35152_/Q _35088_/Q _32272_/Q _16092_/X _16094_/X VGND VGND VPWR
+ VPWR _18121_/X sky130_fd_sc_hd__mux4_1
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27319_ _27367_/S VGND VGND VPWR VPWR _27338_/S sky130_fd_sc_hd__buf_6
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28299_ _27720_/X _34479_/Q _28307_/S VGND VGND VPWR VPWR _28300_/A sky130_fd_sc_hd__mux2_1
X_30330_ _30330_/A VGND VGND VPWR VPWR _35410_/D sky130_fd_sc_hd__clkbuf_1
X_18052_ _18048_/X _18051_/X _17846_/X _17847_/X VGND VGND VPWR VPWR _18067_/B sky130_fd_sc_hd__o211a_1
XFILLER_172_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17003_ _17864_/A VGND VGND VPWR VPWR _17003_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_172_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30261_ _30261_/A VGND VGND VPWR VPWR _35377_/D sky130_fd_sc_hd__clkbuf_1
X_32000_ _36202_/CLK _32000_/D VGND VGND VPWR VPWR _32000_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30192_ _35345_/Q _29512_/X _30192_/S VGND VGND VPWR VPWR _30193_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18954_ _18950_/X _18951_/X _18952_/X _18953_/X VGND VGND VPWR VPWR _18954_/X sky130_fd_sc_hd__a22o_1
XFILLER_234_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17905_ _17905_/A VGND VGND VPWR VPWR _17905_/X sky130_fd_sc_hd__buf_4
X_33951_ _36207_/CLK _33951_/D VGND VGND VPWR VPWR _33951_/Q sky130_fd_sc_hd__dfxtp_1
X_18885_ _18881_/X _18884_/X _18745_/X VGND VGND VPWR VPWR _18895_/C sky130_fd_sc_hd__o21ba_1
XTAP_6780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32902_ _32903_/CLK _32902_/D VGND VGND VPWR VPWR _32902_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17836_ _33928_/Q _33864_/Q _33800_/Q _36104_/Q _17730_/X _17731_/X VGND VGND VPWR
+ VPWR _17836_/X sky130_fd_sc_hd__mux4_1
X_33882_ _36058_/CLK _33882_/D VGND VGND VPWR VPWR _33882_/Q sky130_fd_sc_hd__dfxtp_1
X_35621_ _35625_/CLK _35621_/D VGND VGND VPWR VPWR _35621_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32833_ _35970_/CLK _32833_/D VGND VGND VPWR VPWR _32833_/Q sky130_fd_sc_hd__dfxtp_1
X_17767_ _32646_/Q _32582_/Q _32518_/Q _35974_/Q _17629_/X _17766_/X VGND VGND VPWR
+ VPWR _17767_/X sky130_fd_sc_hd__mux4_1
XFILLER_130_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_424_CLK clkbuf_6_33__f_CLK/X VGND VGND VPWR VPWR _35764_/CLK sky130_fd_sc_hd__clkbuf_16
X_19506_ _20212_/A VGND VGND VPWR VPWR _19506_/X sky130_fd_sc_hd__buf_6
XFILLER_235_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35552_ _35553_/CLK _35552_/D VGND VGND VPWR VPWR _35552_/Q sky130_fd_sc_hd__dfxtp_1
X_16718_ _17915_/A VGND VGND VPWR VPWR _16718_/X sky130_fd_sc_hd__clkbuf_4
X_32764_ _32895_/CLK _32764_/D VGND VGND VPWR VPWR _32764_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17698_ _32132_/Q _32324_/Q _32388_/Q _35908_/Q _17633_/X _17421_/X VGND VGND VPWR
+ VPWR _17698_/X sky130_fd_sc_hd__mux4_1
XFILLER_63_974 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34503_ _34633_/CLK _34503_/D VGND VGND VPWR VPWR _34503_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31715_ _36066_/Q input4/X _31729_/S VGND VGND VPWR VPWR _31716_/A sky130_fd_sc_hd__mux2_1
X_19437_ _32116_/Q _32308_/Q _32372_/Q _35892_/Q _19227_/X _19368_/X VGND VGND VPWR
+ VPWR _19437_/X sky130_fd_sc_hd__mux4_1
X_35483_ _35547_/CLK _35483_/D VGND VGND VPWR VPWR _35483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16649_ _16645_/X _16646_/X _16647_/X _16648_/X VGND VGND VPWR VPWR _16649_/X sky130_fd_sc_hd__a22o_1
X_32695_ _32887_/CLK _32695_/D VGND VGND VPWR VPWR _32695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34434_ _34690_/CLK _34434_/D VGND VGND VPWR VPWR _34434_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31646_ _31646_/A VGND VGND VPWR VPWR _36033_/D sky130_fd_sc_hd__clkbuf_1
X_19368_ _20074_/A VGND VGND VPWR VPWR _19368_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_188_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18319_ _18361_/A VGND VGND VPWR VPWR _20282_/A sky130_fd_sc_hd__buf_12
X_34365_ _35644_/CLK _34365_/D VGND VGND VPWR VPWR _34365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31577_ _31577_/A VGND VGND VPWR VPWR _36000_/D sky130_fd_sc_hd__clkbuf_1
X_19299_ _35696_/Q _32204_/Q _35568_/Q _35504_/Q _19264_/X _19265_/X VGND VGND VPWR
+ VPWR _19299_/X sky130_fd_sc_hd__mux4_1
XFILLER_241_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36104_ _36104_/CLK _36104_/D VGND VGND VPWR VPWR _36104_/Q sky130_fd_sc_hd__dfxtp_1
X_33316_ _33828_/CLK _33316_/D VGND VGND VPWR VPWR _33316_/Q sky130_fd_sc_hd__dfxtp_1
X_21330_ _34664_/Q _34600_/Q _34536_/Q _34472_/Q _21186_/X _21187_/X VGND VGND VPWR
+ VPWR _21330_/X sky130_fd_sc_hd__mux4_1
XFILLER_176_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30528_ _35504_/Q _29410_/X _30534_/S VGND VGND VPWR VPWR _30529_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34296_ _35192_/CLK _34296_/D VGND VGND VPWR VPWR _34296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36035_ _36037_/CLK _36035_/D VGND VGND VPWR VPWR _36035_/Q sky130_fd_sc_hd__dfxtp_1
X_30459_ _30459_/A VGND VGND VPWR VPWR _35471_/D sky130_fd_sc_hd__clkbuf_1
X_33247_ _35615_/CLK _33247_/D VGND VGND VPWR VPWR _33247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21261_ _34406_/Q _36134_/Q _34278_/Q _34214_/Q _21123_/X _21124_/X VGND VGND VPWR
+ VPWR _21261_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23000_ _22999_/X _32058_/Q _23009_/S VGND VGND VPWR VPWR _23001_/A sky130_fd_sc_hd__mux2_1
X_20212_ _20212_/A VGND VGND VPWR VPWR _20212_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_117_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21192_ _34916_/Q _34852_/Q _34788_/Q _34724_/Q _21054_/X _21055_/X VGND VGND VPWR
+ VPWR _21192_/X sky130_fd_sc_hd__mux4_1
X_33178_ _36211_/CLK _33178_/D VGND VGND VPWR VPWR _33178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20143_ _32136_/Q _32328_/Q _32392_/Q _35912_/Q _19933_/X _20074_/X VGND VGND VPWR
+ VPWR _20143_/X sky130_fd_sc_hd__mux4_1
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32129_ _35969_/CLK _32129_/D VGND VGND VPWR VPWR _32129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24951_ input44/X VGND VGND VPWR VPWR _24951_/X sky130_fd_sc_hd__buf_4
X_20074_ _20074_/A VGND VGND VPWR VPWR _20074_/X sky130_fd_sc_hd__clkbuf_4
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23902_ _22971_/X _32497_/Q _23906_/S VGND VGND VPWR VPWR _23903_/A sky130_fd_sc_hd__mux2_1
XTAP_4129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27670_ input64/X VGND VGND VPWR VPWR _27670_/X sky130_fd_sc_hd__buf_4
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24882_ _24882_/A VGND VGND VPWR VPWR _32944_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26621_ _26621_/A VGND VGND VPWR VPWR _33748_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23833_ _23833_/A VGND VGND VPWR VPWR _32401_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35819_ _35820_/CLK _35819_/D VGND VGND VPWR VPWR _35819_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_415_CLK clkbuf_6_32__f_CLK/X VGND VGND VPWR VPWR _35632_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29340_ _34969_/Q _29339_/X _29358_/S VGND VGND VPWR VPWR _29341_/A sky130_fd_sc_hd__mux2_1
X_26552_ _26552_/A VGND VGND VPWR VPWR _33715_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23764_ _23764_/A VGND VGND VPWR VPWR _32368_/D sky130_fd_sc_hd__clkbuf_1
X_20976_ _20970_/X _20975_/X _20675_/X VGND VGND VPWR VPWR _20984_/C sky130_fd_sc_hd__o21ba_1
XFILLER_246_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25503_ _24939_/X _33219_/Q _25511_/S VGND VGND VPWR VPWR _25504_/A sky130_fd_sc_hd__mux2_1
XFILLER_198_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22715_ _20581_/X _22713_/X _22714_/X _20591_/X VGND VGND VPWR VPWR _22715_/X sky130_fd_sc_hd__a22o_1
XFILLER_183_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29271_ _29271_/A VGND VGND VPWR VPWR _34938_/D sky130_fd_sc_hd__clkbuf_1
X_26483_ _26483_/A VGND VGND VPWR VPWR _33683_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_207_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23695_ _23695_/A VGND VGND VPWR VPWR _32337_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28222_ _28222_/A VGND VGND VPWR VPWR _34442_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25434_ _24837_/X _33186_/Q _25448_/S VGND VGND VPWR VPWR _25435_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22646_ _32654_/Q _32590_/Q _32526_/Q _35982_/Q _22582_/X _22366_/X VGND VGND VPWR
+ VPWR _22646_/X sky130_fd_sc_hd__mux4_1
XFILLER_201_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28153_ _28243_/S VGND VGND VPWR VPWR _28172_/S sky130_fd_sc_hd__buf_4
X_25365_ _25365_/A VGND VGND VPWR VPWR _33154_/D sky130_fd_sc_hd__clkbuf_1
X_22577_ _22505_/X _22575_/X _22576_/X _22510_/X VGND VGND VPWR VPWR _22577_/X sky130_fd_sc_hd__a22o_1
XFILLER_51_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27104_ _33964_/Q _27103_/X _27125_/S VGND VGND VPWR VPWR _27105_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24316_ _22974_/X _32690_/Q _24318_/S VGND VGND VPWR VPWR _24317_/A sky130_fd_sc_hd__mux2_1
X_28084_ _34377_/Q _27193_/X _28100_/S VGND VGND VPWR VPWR _28085_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21528_ _32110_/Q _32302_/Q _32366_/Q _35886_/Q _21527_/X _21315_/X VGND VGND VPWR
+ VPWR _21528_/X sky130_fd_sc_hd__mux4_1
X_25296_ _25296_/A VGND VGND VPWR VPWR _33121_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27035_ _27230_/S VGND VGND VPWR VPWR _27063_/S sky130_fd_sc_hd__buf_8
X_24247_ _32659_/Q _23492_/X _24251_/S VGND VGND VPWR VPWR _24248_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21459_ _32620_/Q _32556_/Q _32492_/Q _35948_/Q _21170_/X _21307_/X VGND VGND VPWR
+ VPWR _21459_/X sky130_fd_sc_hd__mux4_1
XFILLER_135_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24178_ _32626_/Q _23381_/X _24180_/S VGND VGND VPWR VPWR _24179_/A sky130_fd_sc_hd__mux2_1
XTAP_6010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23129_ _22943_/X _32104_/Q _23131_/S VGND VGND VPWR VPWR _23130_/A sky130_fd_sc_hd__mux2_1
XTAP_6021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28986_ _28986_/A VGND VGND VPWR VPWR _34803_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_6_62__f_CLK clkbuf_5_31_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_62__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XTAP_6043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput97 _31974_/Q VGND VGND VPWR VPWR D1[16] sky130_fd_sc_hd__buf_2
XTAP_6065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27937_ _27937_/A VGND VGND VPWR VPWR _34307_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18670_ _18592_/X _18668_/X _18669_/X _18595_/X VGND VGND VPWR VPWR _18670_/X sky130_fd_sc_hd__a22o_1
XFILLER_209_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27868_ _27868_/A VGND VGND VPWR VPWR _34274_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_248_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17621_ _17621_/A VGND VGND VPWR VPWR _32001_/D sky130_fd_sc_hd__buf_4
XFILLER_36_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29607_ _29607_/A VGND VGND VPWR VPWR _35067_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_236_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26819_ _33840_/Q _23340_/X _26825_/S VGND VGND VPWR VPWR _26820_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27799_ _27797_/X _34248_/Q _27826_/S VGND VGND VPWR VPWR _27800_/A sky130_fd_sc_hd__mux2_1
XTAP_4685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_406_CLK clkbuf_6_34__f_CLK/X VGND VGND VPWR VPWR _36085_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17552_ _17905_/A VGND VGND VPWR VPWR _17552_/X sky130_fd_sc_hd__clkbuf_4
X_29538_ _29538_/A VGND VGND VPWR VPWR _35034_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16503_ _17869_/A VGND VGND VPWR VPWR _16503_/X sky130_fd_sc_hd__buf_4
XFILLER_60_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17483_ _33918_/Q _33854_/Q _33790_/Q _36094_/Q _17377_/X _17378_/X VGND VGND VPWR
+ VPWR _17483_/X sky130_fd_sc_hd__mux4_1
XFILLER_45_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29469_ input40/X VGND VGND VPWR VPWR _29469_/X sky130_fd_sc_hd__buf_2
XFILLER_225_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19222_ _19218_/X _19221_/X _19079_/X VGND VGND VPWR VPWR _19248_/A sky130_fd_sc_hd__o21ba_1
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31500_ _31500_/A VGND VGND VPWR VPWR _35964_/D sky130_fd_sc_hd__clkbuf_1
X_16434_ _17846_/A VGND VGND VPWR VPWR _16434_/X sky130_fd_sc_hd__buf_2
XFILLER_176_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32480_ _35938_/CLK _32480_/D VGND VGND VPWR VPWR _32480_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31431_ _31431_/A VGND VGND VPWR VPWR _35931_/D sky130_fd_sc_hd__clkbuf_1
X_16365_ _17915_/A VGND VGND VPWR VPWR _16365_/X sky130_fd_sc_hd__clkbuf_4
X_19153_ _20212_/A VGND VGND VPWR VPWR _19153_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_13_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_1243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18104_ _17912_/X _18102_/X _18103_/X _17915_/X VGND VGND VPWR VPWR _18104_/X sky130_fd_sc_hd__a22o_1
X_34150_ _34790_/CLK _34150_/D VGND VGND VPWR VPWR _34150_/Q sky130_fd_sc_hd__dfxtp_1
X_31362_ _27757_/X _35899_/Q _31366_/S VGND VGND VPWR VPWR _31363_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16296_ _16292_/X _16293_/X _16294_/X _16295_/X VGND VGND VPWR VPWR _16296_/X sky130_fd_sc_hd__a22o_1
X_19084_ _32106_/Q _32298_/Q _32362_/Q _35882_/Q _18874_/X _19015_/X VGND VGND VPWR
+ VPWR _19084_/X sky130_fd_sc_hd__mux4_1
XFILLER_9_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30313_ _35402_/Q _29491_/X _30327_/S VGND VGND VPWR VPWR _30314_/A sky130_fd_sc_hd__mux2_1
X_33101_ _35852_/CLK _33101_/D VGND VGND VPWR VPWR _33101_/Q sky130_fd_sc_hd__dfxtp_1
X_18035_ _17864_/X _18033_/X _18034_/X _17869_/X VGND VGND VPWR VPWR _18035_/X sky130_fd_sc_hd__a22o_1
X_31293_ _27655_/X _35866_/Q _31303_/S VGND VGND VPWR VPWR _31294_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34081_ _34594_/CLK _34081_/D VGND VGND VPWR VPWR _34081_/Q sky130_fd_sc_hd__dfxtp_1
X_33032_ _35785_/CLK _33032_/D VGND VGND VPWR VPWR _33032_/Q sky130_fd_sc_hd__dfxtp_1
X_30244_ _30244_/A VGND VGND VPWR VPWR _35369_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30175_ _30175_/A VGND VGND VPWR VPWR _35336_/D sky130_fd_sc_hd__clkbuf_1
X_19986_ _19986_/A _19986_/B _19986_/C _19986_/D VGND VGND VPWR VPWR _19987_/A sky130_fd_sc_hd__or4_4
XFILLER_119_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18937_ _33126_/Q _36006_/Q _32998_/Q _32934_/Q _18656_/X _18657_/X VGND VGND VPWR
+ VPWR _18937_/X sky130_fd_sc_hd__mux4_1
X_34983_ _35622_/CLK _34983_/D VGND VGND VPWR VPWR _34983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33934_ _33934_/CLK _33934_/D VGND VGND VPWR VPWR _33934_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18868_ _18800_/X _18866_/X _18867_/X _18803_/X VGND VGND VPWR VPWR _18868_/X sky130_fd_sc_hd__a22o_1
XFILLER_41_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17819_ _17709_/X _17817_/X _17818_/X _17712_/X VGND VGND VPWR VPWR _17819_/X sky130_fd_sc_hd__a22o_1
XFILLER_39_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33865_ _36105_/CLK _33865_/D VGND VGND VPWR VPWR _33865_/Q sky130_fd_sc_hd__dfxtp_1
X_18799_ _18793_/X _18796_/X _18797_/X _18798_/X VGND VGND VPWR VPWR _18799_/X sky130_fd_sc_hd__a22o_1
XFILLER_243_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_242_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35604_ _35668_/CLK _35604_/D VGND VGND VPWR VPWR _35604_/Q sky130_fd_sc_hd__dfxtp_1
X_20830_ _33050_/Q _32026_/Q _35802_/Q _35738_/Q _20667_/X _20669_/X VGND VGND VPWR
+ VPWR _20830_/X sky130_fd_sc_hd__mux4_1
X_32816_ _32909_/CLK _32816_/D VGND VGND VPWR VPWR _32816_/Q sky130_fd_sc_hd__dfxtp_1
X_33796_ _36097_/CLK _33796_/D VGND VGND VPWR VPWR _33796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35535_ _35727_/CLK _35535_/D VGND VGND VPWR VPWR _35535_/Q sky130_fd_sc_hd__dfxtp_1
X_20761_ _35608_/Q _34968_/Q _34328_/Q _33688_/Q _20653_/X _20655_/X VGND VGND VPWR
+ VPWR _20761_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32747_ _35946_/CLK _32747_/D VGND VGND VPWR VPWR _32747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22500_ _34953_/Q _34889_/Q _34825_/Q _34761_/Q _22466_/X _22467_/X VGND VGND VPWR
+ VPWR _22500_/X sky130_fd_sc_hd__mux4_1
X_23480_ _23480_/A VGND VGND VPWR VPWR _32238_/D sky130_fd_sc_hd__clkbuf_1
X_35466_ _35466_/CLK _35466_/D VGND VGND VPWR VPWR _35466_/Q sky130_fd_sc_hd__dfxtp_1
X_20692_ _22316_/A VGND VGND VPWR VPWR _20692_/X sky130_fd_sc_hd__clkbuf_8
X_32678_ _32873_/CLK _32678_/D VGND VGND VPWR VPWR _32678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22431_ _34184_/Q _34120_/Q _34056_/Q _33992_/Q _22399_/X _22400_/X VGND VGND VPWR
+ VPWR _22431_/X sky130_fd_sc_hd__mux4_1
XFILLER_56_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34417_ _36144_/CLK _34417_/D VGND VGND VPWR VPWR _34417_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31629_ _31629_/A VGND VGND VPWR VPWR _36025_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35397_ _35463_/CLK _35397_/D VGND VGND VPWR VPWR _35397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25150_ _33053_/Q _23252_/X _25154_/S VGND VGND VPWR VPWR _25151_/A sky130_fd_sc_hd__mux2_1
X_22362_ _33926_/Q _33862_/Q _33798_/Q _36102_/Q _22330_/X _22331_/X VGND VGND VPWR
+ VPWR _22362_/X sky130_fd_sc_hd__mux4_1
X_34348_ _35692_/CLK _34348_/D VGND VGND VPWR VPWR _34348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24101_ _23064_/X _32591_/Q _24105_/S VGND VGND VPWR VPWR _24102_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21313_ _21306_/X _21308_/X _21311_/X _21312_/X VGND VGND VPWR VPWR _21313_/X sky130_fd_sc_hd__a22o_1
X_25081_ _25081_/A VGND VGND VPWR VPWR _33021_/D sky130_fd_sc_hd__clkbuf_1
X_22293_ _22159_/X _22291_/X _22292_/X _22162_/X VGND VGND VPWR VPWR _22293_/X sky130_fd_sc_hd__a22o_1
XFILLER_184_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34279_ _35554_/CLK _34279_/D VGND VGND VPWR VPWR _34279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36018_ _36019_/CLK _36018_/D VGND VGND VPWR VPWR _36018_/Q sky130_fd_sc_hd__dfxtp_1
X_24032_ _22962_/X _32558_/Q _24042_/S VGND VGND VPWR VPWR _24033_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21244_ _21238_/X _21243_/X _21034_/X _21035_/X VGND VGND VPWR VPWR _21265_/B sky130_fd_sc_hd__o211a_1
XFILLER_137_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28840_ _34734_/Q _27109_/X _28850_/S VGND VGND VPWR VPWR _28841_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21175_ _32100_/Q _32292_/Q _32356_/Q _35876_/Q _21174_/X _20962_/X VGND VGND VPWR
+ VPWR _21175_/X sky130_fd_sc_hd__mux4_1
XFILLER_172_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20126_ _19811_/X _20124_/X _20125_/X _19816_/X VGND VGND VPWR VPWR _20126_/X sky130_fd_sc_hd__a22o_1
X_28771_ _28771_/A VGND VGND VPWR VPWR _34702_/D sky130_fd_sc_hd__clkbuf_1
X_25983_ _25983_/A VGND VGND VPWR VPWR _33446_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_219_803 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20057_ _20057_/A VGND VGND VPWR VPWR _32453_/D sky130_fd_sc_hd__clkbuf_4
X_24934_ _24933_/X _32961_/Q _24952_/S VGND VGND VPWR VPWR _24935_/A sky130_fd_sc_hd__mux2_1
X_27722_ _27722_/A VGND VGND VPWR VPWR _34223_/D sky130_fd_sc_hd__clkbuf_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27653_ _27652_/X _34201_/Q _27671_/S VGND VGND VPWR VPWR _27654_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24865_ input14/X VGND VGND VPWR VPWR _24865_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26604_ _24967_/X _33740_/Q _26614_/S VGND VGND VPWR VPWR _26605_/A sky130_fd_sc_hd__mux2_1
X_23816_ _23046_/X _32393_/Q _23832_/S VGND VGND VPWR VPWR _23817_/A sky130_fd_sc_hd__mux2_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27584_ _27584_/A VGND VGND VPWR VPWR _34171_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24796_ input1/X VGND VGND VPWR VPWR _24796_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29323_ _29323_/A VGND VGND VPWR VPWR _34963_/D sky130_fd_sc_hd__clkbuf_1
X_26535_ _24865_/X _33707_/Q _26551_/S VGND VGND VPWR VPWR _26536_/A sky130_fd_sc_hd__mux2_1
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23747_ _23747_/A VGND VGND VPWR VPWR _32360_/D sky130_fd_sc_hd__clkbuf_1
X_20959_ _22510_/A VGND VGND VPWR VPWR _20959_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_42_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_916 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26466_ _33675_/Q _23466_/X _26478_/S VGND VGND VPWR VPWR _26467_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29254_ _29254_/A VGND VGND VPWR VPWR _34930_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23678_ _23046_/X _32329_/Q _23694_/S VGND VGND VPWR VPWR _23679_/A sky130_fd_sc_hd__mux2_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28205_ _28205_/A VGND VGND VPWR VPWR _34434_/D sky130_fd_sc_hd__clkbuf_1
X_25417_ _24812_/X _33178_/Q _25427_/S VGND VGND VPWR VPWR _25418_/A sky130_fd_sc_hd__mux2_1
X_29185_ _34898_/Q _27220_/X _29191_/S VGND VGND VPWR VPWR _29186_/A sky130_fd_sc_hd__mux2_1
X_22629_ _22625_/X _22628_/X _22457_/X VGND VGND VPWR VPWR _22637_/C sky130_fd_sc_hd__o21ba_1
XFILLER_167_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26397_ _33642_/Q _23292_/X _26415_/S VGND VGND VPWR VPWR _26398_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28136_ _28136_/A VGND VGND VPWR VPWR _34401_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16150_ _17869_/A VGND VGND VPWR VPWR _16150_/X sky130_fd_sc_hd__buf_6
XFILLER_6_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25348_ _25348_/A VGND VGND VPWR VPWR _33146_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16081_ _34646_/Q _34582_/Q _34518_/Q _34454_/Q _16079_/X _16080_/X VGND VGND VPWR
+ VPWR _16081_/X sky130_fd_sc_hd__mux4_1
X_28067_ _34369_/Q _27168_/X _28079_/S VGND VGND VPWR VPWR _28068_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25279_ _25279_/A VGND VGND VPWR VPWR _33113_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27018_ _27018_/A VGND VGND VPWR VPWR _33934_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_1271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19840_ _33087_/Q _32063_/Q _35839_/Q _35775_/Q _19731_/X _19732_/X VGND VGND VPWR
+ VPWR _19840_/X sky130_fd_sc_hd__mux4_1
XFILLER_190_1236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19771_ _34429_/Q _36157_/Q _34301_/Q _34237_/Q _19529_/X _19530_/X VGND VGND VPWR
+ VPWR _19771_/X sky130_fd_sc_hd__mux4_1
X_16983_ _34160_/Q _34096_/Q _34032_/Q _33968_/Q _16740_/X _16741_/X VGND VGND VPWR
+ VPWR _16983_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28969_ _34795_/Q _27100_/X _28985_/S VGND VGND VPWR VPWR _28970_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18722_ _20100_/A VGND VGND VPWR VPWR _18722_/X sky130_fd_sc_hd__buf_4
XTAP_5150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31980_ _34790_/CLK _31980_/D VGND VGND VPWR VPWR _31980_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18653_ _20205_/A VGND VGND VPWR VPWR _18653_/X sky130_fd_sc_hd__clkbuf_4
X_30931_ _35695_/Q input18/X _30939_/S VGND VGND VPWR VPWR _30932_/A sky130_fd_sc_hd__mux2_1
XTAP_4460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17604_ _35713_/Q _32223_/Q _35585_/Q _35521_/Q _17317_/X _17318_/X VGND VGND VPWR
+ VPWR _17604_/X sky130_fd_sc_hd__mux4_1
XTAP_4493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33650_ _34098_/CLK _33650_/D VGND VGND VPWR VPWR _33650_/Q sky130_fd_sc_hd__dfxtp_1
X_30862_ _30862_/A VGND VGND VPWR VPWR _35662_/D sky130_fd_sc_hd__clkbuf_1
X_18584_ _33116_/Q _35996_/Q _32988_/Q _32924_/Q _18324_/X _18325_/X VGND VGND VPWR
+ VPWR _18584_/X sky130_fd_sc_hd__mux4_1
XTAP_3770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32601_ _34135_/CLK _32601_/D VGND VGND VPWR VPWR _32601_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17535_ _17531_/X _17534_/X _17493_/X _17494_/X VGND VGND VPWR VPWR _17550_/B sky130_fd_sc_hd__o211a_1
XFILLER_33_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33581_ _36077_/CLK _33581_/D VGND VGND VPWR VPWR _33581_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30793_ _30793_/A VGND VGND VPWR VPWR _35629_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35320_ _35320_/CLK _35320_/D VGND VGND VPWR VPWR _35320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_232_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32532_ _35988_/CLK _32532_/D VGND VGND VPWR VPWR _32532_/Q sky130_fd_sc_hd__dfxtp_1
X_17466_ _17356_/X _17464_/X _17465_/X _17359_/X VGND VGND VPWR VPWR _17466_/X sky130_fd_sc_hd__a22o_1
XFILLER_220_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19205_ _18950_/X _19203_/X _19204_/X _18953_/X VGND VGND VPWR VPWR _19205_/X sky130_fd_sc_hd__a22o_1
XFILLER_60_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16417_ _16417_/A VGND VGND VPWR VPWR _31967_/D sky130_fd_sc_hd__clkbuf_1
X_35251_ _35764_/CLK _35251_/D VGND VGND VPWR VPWR _35251_/Q sky130_fd_sc_hd__dfxtp_1
X_32463_ _33904_/CLK _32463_/D VGND VGND VPWR VPWR _32463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_1324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_919 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17397_ _35195_/Q _35131_/Q _35067_/Q _32251_/Q _17363_/X _17364_/X VGND VGND VPWR
+ VPWR _17397_/X sky130_fd_sc_hd__mux4_1
X_34202_ _36235_/CLK _34202_/D VGND VGND VPWR VPWR _34202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31414_ _27834_/X _35924_/Q _31416_/S VGND VGND VPWR VPWR _31415_/A sky130_fd_sc_hd__mux2_1
X_19136_ _19132_/X _19135_/X _19098_/X VGND VGND VPWR VPWR _19144_/C sky130_fd_sc_hd__o21ba_1
X_16348_ _16140_/X _16346_/X _16347_/X _16145_/X VGND VGND VPWR VPWR _16348_/X sky130_fd_sc_hd__a22o_1
X_35182_ _35183_/CLK _35182_/D VGND VGND VPWR VPWR _35182_/Q sky130_fd_sc_hd__dfxtp_1
X_32394_ _32907_/CLK _32394_/D VGND VGND VPWR VPWR _32394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_218_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34133_ _34773_/CLK _34133_/D VGND VGND VPWR VPWR _34133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16279_ _33372_/Q _33308_/Q _33244_/Q _33180_/Q _16002_/X _16003_/X VGND VGND VPWR
+ VPWR _16279_/X sky130_fd_sc_hd__mux4_1
X_19067_ _18752_/X _19065_/X _19066_/X _18757_/X VGND VGND VPWR VPWR _19067_/X sky130_fd_sc_hd__a22o_1
X_31345_ _27732_/X _35891_/Q _31345_/S VGND VGND VPWR VPWR _31346_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_805 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18018_ _17765_/X _18016_/X _18017_/X _17771_/X VGND VGND VPWR VPWR _18018_/X sky130_fd_sc_hd__a22o_1
X_34064_ _34064_/CLK _34064_/D VGND VGND VPWR VPWR _34064_/Q sky130_fd_sc_hd__dfxtp_1
X_31276_ _31276_/A VGND VGND VPWR VPWR _35858_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33015_ _34485_/CLK _33015_/D VGND VGND VPWR VPWR _33015_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30227_ _35361_/Q _29364_/X _30243_/S VGND VGND VPWR VPWR _30228_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30158_ _30158_/A VGND VGND VPWR VPWR _35328_/D sky130_fd_sc_hd__clkbuf_1
X_19969_ _19965_/X _19968_/X _19793_/X _19794_/X VGND VGND VPWR VPWR _19986_/B sky130_fd_sc_hd__o211a_1
XFILLER_234_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34966_ _35735_/CLK _34966_/D VGND VGND VPWR VPWR _34966_/Q sky130_fd_sc_hd__dfxtp_1
X_22980_ input24/X VGND VGND VPWR VPWR _22980_/X sky130_fd_sc_hd__clkbuf_4
X_30089_ _30200_/S VGND VGND VPWR VPWR _30108_/S sky130_fd_sc_hd__clkbuf_8
X_33917_ _36093_/CLK _33917_/D VGND VGND VPWR VPWR _33917_/Q sky130_fd_sc_hd__dfxtp_1
X_21931_ _21758_/X _21929_/X _21930_/X _21763_/X VGND VGND VPWR VPWR _21931_/X sky130_fd_sc_hd__a22o_1
XFILLER_95_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34897_ _34897_/CLK _34897_/D VGND VGND VPWR VPWR _34897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24650_ _24650_/A VGND VGND VPWR VPWR _32848_/D sky130_fd_sc_hd__clkbuf_1
X_33848_ _33911_/CLK _33848_/D VGND VGND VPWR VPWR _33848_/Q sky130_fd_sc_hd__dfxtp_1
X_21862_ _21753_/X _21860_/X _21861_/X _21756_/X VGND VGND VPWR VPWR _21862_/X sky130_fd_sc_hd__a22o_1
XFILLER_82_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23601_ _23601_/A VGND VGND VPWR VPWR _32292_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20813_ _33370_/Q _33306_/Q _33242_/Q _33178_/Q _20602_/X _20603_/X VGND VGND VPWR
+ VPWR _20813_/X sky130_fd_sc_hd__mux4_1
X_24581_ _24581_/A VGND VGND VPWR VPWR _32815_/D sky130_fd_sc_hd__clkbuf_1
X_33779_ _36085_/CLK _33779_/D VGND VGND VPWR VPWR _33779_/Q sky130_fd_sc_hd__dfxtp_1
X_21793_ _34421_/Q _36149_/Q _34293_/Q _34229_/Q _21476_/X _21477_/X VGND VGND VPWR
+ VPWR _21793_/X sky130_fd_sc_hd__mux4_1
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26320_ _26320_/A VGND VGND VPWR VPWR _33606_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_223_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23532_ _32261_/Q _23444_/X _23536_/S VGND VGND VPWR VPWR _23533_/A sky130_fd_sc_hd__mux2_1
X_35518_ _36095_/CLK _35518_/D VGND VGND VPWR VPWR _35518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_243_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20744_ _34136_/Q _34072_/Q _34008_/Q _33944_/Q _20609_/X _20611_/X VGND VGND VPWR
+ VPWR _20744_/X sky130_fd_sc_hd__mux4_1
XFILLER_223_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26251_ _26251_/A VGND VGND VPWR VPWR _33573_/D sky130_fd_sc_hd__clkbuf_1
X_23463_ input48/X VGND VGND VPWR VPWR _23463_/X sky130_fd_sc_hd__buf_4
X_35449_ _35449_/CLK _35449_/D VGND VGND VPWR VPWR _35449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20675_ _22457_/A VGND VGND VPWR VPWR _20675_/X sky130_fd_sc_hd__buf_4
XFILLER_52_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25202_ _25202_/A VGND VGND VPWR VPWR _33077_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22414_ _35719_/Q _32229_/Q _35591_/Q _35527_/Q _22270_/X _22271_/X VGND VGND VPWR
+ VPWR _22414_/X sky130_fd_sc_hd__mux4_1
XFILLER_155_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26182_ _24945_/X _33541_/Q _26186_/S VGND VGND VPWR VPWR _26183_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_824 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23394_ _32210_/Q _23393_/X _23418_/S VGND VGND VPWR VPWR _23395_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25133_ _25133_/A VGND VGND VPWR VPWR _30337_/A sky130_fd_sc_hd__buf_6
X_22345_ _35461_/Q _35397_/Q _35333_/Q _35269_/Q _22207_/X _22208_/X VGND VGND VPWR
+ VPWR _22345_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29941_ _29941_/A VGND VGND VPWR VPWR _35225_/D sky130_fd_sc_hd__clkbuf_1
X_25064_ _24896_/X _33013_/Q _25080_/S VGND VGND VPWR VPWR _25065_/A sky130_fd_sc_hd__mux2_1
X_22276_ _33091_/Q _32067_/Q _35843_/Q _35779_/Q _22031_/X _22032_/X VGND VGND VPWR
+ VPWR _22276_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24015_ _22937_/X _32550_/Q _24021_/S VGND VGND VPWR VPWR _24016_/A sky130_fd_sc_hd__mux2_1
X_21227_ _21227_/A _21227_/B _21227_/C _21227_/D VGND VGND VPWR VPWR _21228_/A sky130_fd_sc_hd__or4_1
XFILLER_176_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29872_ _35193_/Q _29438_/X _29880_/S VGND VGND VPWR VPWR _29873_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_754 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28823_ _34726_/Q _27084_/X _28829_/S VGND VGND VPWR VPWR _28824_/A sky130_fd_sc_hd__mux2_1
X_21158_ _34915_/Q _34851_/Q _34787_/Q _34723_/Q _21054_/X _21055_/X VGND VGND VPWR
+ VPWR _21158_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20109_ _20065_/X _20107_/X _20108_/X _20071_/X VGND VGND VPWR VPWR _20109_/X sky130_fd_sc_hd__a22o_1
XFILLER_28_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28754_ _28754_/A VGND VGND VPWR VPWR _34694_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_863 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25966_ _25966_/A VGND VGND VPWR VPWR _33438_/D sky130_fd_sc_hd__clkbuf_1
X_21089_ _21052_/X _21087_/X _21088_/X _21057_/X VGND VGND VPWR VPWR _21089_/X sky130_fd_sc_hd__a22o_1
XFILLER_247_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27705_ _27838_/S VGND VGND VPWR VPWR _27733_/S sky130_fd_sc_hd__buf_4
XTAP_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24917_ input32/X VGND VGND VPWR VPWR _24917_/X sky130_fd_sc_hd__clkbuf_4
X_25897_ _25945_/S VGND VGND VPWR VPWR _25916_/S sky130_fd_sc_hd__buf_4
X_28685_ _28685_/A VGND VGND VPWR VPWR _34661_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_233_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27636_ _27636_/A VGND VGND VPWR VPWR _34196_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_233_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24848_ _24848_/A VGND VGND VPWR VPWR _32933_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24779_ _24779_/A VGND VGND VPWR VPWR _32909_/D sky130_fd_sc_hd__clkbuf_1
X_27567_ _27567_/A VGND VGND VPWR VPWR _34163_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_730 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29306_ _34955_/Q _27199_/X _29318_/S VGND VGND VPWR VPWR _29307_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_1051 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17320_ _35641_/Q _35001_/Q _34361_/Q _33721_/Q _17144_/X _17145_/X VGND VGND VPWR
+ VPWR _17320_/X sky130_fd_sc_hd__mux4_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26518_ _24840_/X _33699_/Q _26530_/S VGND VGND VPWR VPWR _26519_/A sky130_fd_sc_hd__mux2_1
X_27498_ _34131_/Q _27223_/X _27502_/S VGND VGND VPWR VPWR _27499_/A sky130_fd_sc_hd__mux2_1
XFILLER_187_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17251_ _35703_/Q _32212_/Q _35575_/Q _35511_/Q _16964_/X _16965_/X VGND VGND VPWR
+ VPWR _17251_/X sky130_fd_sc_hd__mux4_1
X_29237_ _34922_/Q _27096_/X _29255_/S VGND VGND VPWR VPWR _29238_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26449_ _33667_/Q _23438_/X _26457_/S VGND VGND VPWR VPWR _26450_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16202_ _35161_/Q _35097_/Q _35033_/Q _32153_/Q _16083_/X _16085_/X VGND VGND VPWR
+ VPWR _16202_/X sky130_fd_sc_hd__mux4_1
XFILLER_224_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17182_ _17178_/X _17181_/X _17140_/X _17141_/X VGND VGND VPWR VPWR _17197_/B sky130_fd_sc_hd__o211a_1
X_29168_ _29168_/A VGND VGND VPWR VPWR _34889_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16133_ _16078_/X _16131_/X _16132_/X _16088_/X VGND VGND VPWR VPWR _16133_/X sky130_fd_sc_hd__a22o_1
XFILLER_31_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28119_ _28119_/A VGND VGND VPWR VPWR _34393_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29099_ _34857_/Q _27093_/X _29099_/S VGND VGND VPWR VPWR _29100_/A sky130_fd_sc_hd__mux2_1
X_16064_ _17851_/A VGND VGND VPWR VPWR _16064_/X sky130_fd_sc_hd__buf_4
X_31130_ _31130_/A VGND VGND VPWR VPWR _35789_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31061_ _31061_/A VGND VGND VPWR VPWR _35756_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_1180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30012_ _30012_/A VGND VGND VPWR VPWR _35259_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19823_ _34175_/Q _34111_/Q _34047_/Q _33983_/Q _19746_/X _19747_/X VGND VGND VPWR
+ VPWR _19823_/X sky130_fd_sc_hd__mux4_1
XFILLER_111_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1058 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34820_ _36164_/CLK _34820_/D VGND VGND VPWR VPWR _34820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19754_ _32637_/Q _32573_/Q _32509_/Q _35965_/Q _19576_/X _19713_/X VGND VGND VPWR
+ VPWR _19754_/X sky130_fd_sc_hd__mux4_1
XFILLER_133_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16966_ _35695_/Q _32203_/Q _35567_/Q _35503_/Q _16964_/X _16965_/X VGND VGND VPWR
+ VPWR _16966_/X sky130_fd_sc_hd__mux4_1
X_18705_ _35423_/Q _35359_/Q _35295_/Q _35231_/Q _18495_/X _18496_/X VGND VGND VPWR
+ VPWR _18705_/X sky130_fd_sc_hd__mux4_1
X_34751_ _34815_/CLK _34751_/D VGND VGND VPWR VPWR _34751_/Q sky130_fd_sc_hd__dfxtp_1
X_31963_ _34148_/CLK _31963_/D VGND VGND VPWR VPWR _31963_/Q sky130_fd_sc_hd__dfxtp_1
X_19685_ _32123_/Q _32315_/Q _32379_/Q _35899_/Q _19580_/X _19368_/X VGND VGND VPWR
+ VPWR _19685_/X sky130_fd_sc_hd__mux4_1
XFILLER_237_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16897_ _16893_/X _16896_/X _16787_/X _16788_/X VGND VGND VPWR VPWR _16914_/B sky130_fd_sc_hd__o211a_1
X_33702_ _35620_/CLK _33702_/D VGND VGND VPWR VPWR _33702_/Q sky130_fd_sc_hd__dfxtp_1
X_18636_ _18632_/X _18635_/X _18375_/X VGND VGND VPWR VPWR _18644_/C sky130_fd_sc_hd__o21ba_1
X_30914_ _35687_/Q input9/X _30918_/S VGND VGND VPWR VPWR _30915_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34682_ _35197_/CLK _34682_/D VGND VGND VPWR VPWR _34682_/Q sky130_fd_sc_hd__dfxtp_1
X_31894_ _23399_/X _36151_/Q _31906_/S VGND VGND VPWR VPWR _31895_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33633_ _34593_/CLK _33633_/D VGND VGND VPWR VPWR _33633_/Q sky130_fd_sc_hd__dfxtp_1
X_18567_ _34651_/Q _34587_/Q _34523_/Q _34459_/Q _18533_/X _18534_/X VGND VGND VPWR
+ VPWR _18567_/X sky130_fd_sc_hd__mux4_1
X_30845_ _30845_/A VGND VGND VPWR VPWR _35654_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17518_ _17871_/A VGND VGND VPWR VPWR _17518_/X sky130_fd_sc_hd__buf_2
XFILLER_127_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33564_ _36211_/CLK _33564_/D VGND VGND VPWR VPWR _33564_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18498_ _33049_/Q _32025_/Q _35801_/Q _35737_/Q _18367_/X _18369_/X VGND VGND VPWR
+ VPWR _18498_/X sky130_fd_sc_hd__mux4_1
X_30776_ _30776_/A VGND VGND VPWR VPWR _35621_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35303_ _35367_/CLK _35303_/D VGND VGND VPWR VPWR _35303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1029 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32515_ _35907_/CLK _32515_/D VGND VGND VPWR VPWR _32515_/Q sky130_fd_sc_hd__dfxtp_1
X_17449_ _17199_/X _17445_/X _17448_/X _17204_/X VGND VGND VPWR VPWR _17449_/X sky130_fd_sc_hd__a22o_1
X_33495_ _35995_/CLK _33495_/D VGND VGND VPWR VPWR _33495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35234_ _35553_/CLK _35234_/D VGND VGND VPWR VPWR _35234_/Q sky130_fd_sc_hd__dfxtp_1
X_20460_ _34194_/Q _34130_/Q _34066_/Q _34002_/Q _18349_/X _18350_/X VGND VGND VPWR
+ VPWR _20460_/X sky130_fd_sc_hd__mux4_1
X_32446_ _36075_/CLK _32446_/D VGND VGND VPWR VPWR _32446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19119_ _33387_/Q _33323_/Q _33259_/Q _33195_/Q _19074_/X _19075_/X VGND VGND VPWR
+ VPWR _19119_/X sky130_fd_sc_hd__mux4_1
X_35165_ _36219_/CLK _35165_/D VGND VGND VPWR VPWR _35165_/Q sky130_fd_sc_hd__dfxtp_1
X_20391_ _35215_/Q _35151_/Q _35087_/Q _32271_/Q _18392_/X _18394_/X VGND VGND VPWR
+ VPWR _20391_/X sky130_fd_sc_hd__mux4_1
XFILLER_173_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32377_ _32889_/CLK _32377_/D VGND VGND VPWR VPWR _32377_/Q sky130_fd_sc_hd__dfxtp_1
X_34116_ _34180_/CLK _34116_/D VGND VGND VPWR VPWR _34116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_996 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22130_ _33151_/Q _36031_/Q _33023_/Q _32959_/Q _22015_/X _22016_/X VGND VGND VPWR
+ VPWR _22130_/X sky130_fd_sc_hd__mux4_1
XFILLER_173_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31328_ _31328_/A VGND VGND VPWR VPWR _35882_/D sky130_fd_sc_hd__clkbuf_1
Xoutput210 _36242_/Q VGND VGND VPWR VPWR D2[60] sky130_fd_sc_hd__buf_2
X_35096_ _35162_/CLK _35096_/D VGND VGND VPWR VPWR _35096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput221 _32418_/Q VGND VGND VPWR VPWR D3[12] sky130_fd_sc_hd__buf_2
XFILLER_133_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput232 _32428_/Q VGND VGND VPWR VPWR D3[22] sky130_fd_sc_hd__buf_2
XFILLER_86_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34047_ _35454_/CLK _34047_/D VGND VGND VPWR VPWR _34047_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput243 _32438_/Q VGND VGND VPWR VPWR D3[32] sky130_fd_sc_hd__buf_2
X_22061_ _35709_/Q _32218_/Q _35581_/Q _35517_/Q _21917_/X _21918_/X VGND VGND VPWR
+ VPWR _22061_/X sky130_fd_sc_hd__mux4_1
XFILLER_245_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31259_ _27804_/X _35850_/Q _31273_/S VGND VGND VPWR VPWR _31260_/A sky130_fd_sc_hd__mux2_1
Xoutput254 _32448_/Q VGND VGND VPWR VPWR D3[42] sky130_fd_sc_hd__buf_2
XFILLER_114_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput265 _32458_/Q VGND VGND VPWR VPWR D3[52] sky130_fd_sc_hd__buf_2
Xoutput276 _32468_/Q VGND VGND VPWR VPWR D3[62] sky130_fd_sc_hd__buf_2
X_21012_ _34399_/Q _36127_/Q _34271_/Q _34207_/Q _20770_/X _20771_/X VGND VGND VPWR
+ VPWR _21012_/X sky130_fd_sc_hd__mux4_1
XFILLER_138_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25820_ _24809_/X _33369_/Q _25832_/S VGND VGND VPWR VPWR _25821_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35998_ _35998_/CLK _35998_/D VGND VGND VPWR VPWR _35998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25751_ _25751_/A VGND VGND VPWR VPWR _33336_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34949_ _34949_/CLK _34949_/D VGND VGND VPWR VPWR _34949_/Q sky130_fd_sc_hd__dfxtp_1
X_22963_ _22962_/X _32046_/Q _22978_/S VGND VGND VPWR VPWR _22964_/A sky130_fd_sc_hd__mux2_1
XFILLER_244_934 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21914_ _32889_/Q _32825_/Q _32761_/Q _32697_/Q _21593_/X _21594_/X VGND VGND VPWR
+ VPWR _21914_/X sky130_fd_sc_hd__mux4_1
X_24702_ _22946_/X _32873_/Q _24702_/S VGND VGND VPWR VPWR _24703_/A sky130_fd_sc_hd__mux2_1
X_28470_ _27773_/X _34560_/Q _28484_/S VGND VGND VPWR VPWR _28471_/A sky130_fd_sc_hd__mux2_1
X_25682_ _25682_/A VGND VGND VPWR VPWR _33303_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22894_ input23/X VGND VGND VPWR VPWR _22894_/X sky130_fd_sc_hd__buf_2
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24633_ _23042_/X _32840_/Q _24651_/S VGND VGND VPWR VPWR _24634_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27421_ _34094_/Q _27109_/X _27431_/S VGND VGND VPWR VPWR _27422_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21845_ _33143_/Q _36023_/Q _33015_/Q _32951_/Q _21662_/X _21663_/X VGND VGND VPWR
+ VPWR _21845_/X sky130_fd_sc_hd__mux4_1
XFILLER_93_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27352_ _27352_/A VGND VGND VPWR VPWR _34061_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24564_ _24564_/A VGND VGND VPWR VPWR _32807_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21776_ _32629_/Q _32565_/Q _32501_/Q _35957_/Q _21523_/X _21660_/X VGND VGND VPWR
+ VPWR _21776_/X sky130_fd_sc_hd__mux4_1
XFILLER_168_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26303_ _24923_/X _33598_/Q _26321_/S VGND VGND VPWR VPWR _26304_/A sky130_fd_sc_hd__mux2_1
X_23515_ _32253_/Q _23417_/X _23515_/S VGND VGND VPWR VPWR _23516_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20727_ _35415_/Q _35351_/Q _35287_/Q _35223_/Q _20662_/X _20664_/X VGND VGND VPWR
+ VPWR _20727_/X sky130_fd_sc_hd__mux4_1
XFILLER_180_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27283_ _27283_/A VGND VGND VPWR VPWR _34028_/D sky130_fd_sc_hd__clkbuf_1
X_24495_ _23039_/X _32775_/Q _24495_/S VGND VGND VPWR VPWR _24496_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29022_ _29022_/A VGND VGND VPWR VPWR _34820_/D sky130_fd_sc_hd__clkbuf_1
X_26234_ _26234_/A VGND VGND VPWR VPWR _33565_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23446_ _23446_/A VGND VGND VPWR VPWR _32227_/D sky130_fd_sc_hd__clkbuf_1
X_20658_ _22462_/A VGND VGND VPWR VPWR _20658_/X sky130_fd_sc_hd__buf_4
XFILLER_184_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26165_ _24920_/X _33533_/Q _26165_/S VGND VGND VPWR VPWR _26166_/A sky130_fd_sc_hd__mux2_1
XFILLER_221_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23377_ _32204_/Q _23340_/X _23385_/S VGND VGND VPWR VPWR _23378_/A sky130_fd_sc_hd__mux2_1
X_20589_ input73/X input74/X VGND VGND VPWR VPWR _22371_/A sky130_fd_sc_hd__nor2_4
XFILLER_165_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25116_ _24973_/X _33038_/Q _25122_/S VGND VGND VPWR VPWR _25117_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22328_ _22152_/X _22326_/X _22327_/X _22157_/X VGND VGND VPWR VPWR _22328_/X sky130_fd_sc_hd__a22o_1
X_26096_ _24818_/X _33500_/Q _26102_/S VGND VGND VPWR VPWR _26097_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29924_ _35218_/Q _29515_/X _29930_/S VGND VGND VPWR VPWR _29925_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25047_ _24871_/X _33005_/Q _25059_/S VGND VGND VPWR VPWR _25048_/A sky130_fd_sc_hd__mux2_1
XFILLER_219_1150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22259_ _33411_/Q _33347_/Q _33283_/Q _33219_/Q _22080_/X _22081_/X VGND VGND VPWR
+ VPWR _22259_/X sky130_fd_sc_hd__mux4_1
XFILLER_191_1331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29855_ _35185_/Q _29413_/X _29859_/S VGND VGND VPWR VPWR _29856_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28806_ _34718_/Q _27059_/X _28808_/S VGND VGND VPWR VPWR _28807_/A sky130_fd_sc_hd__mux2_1
X_16820_ _33899_/Q _33835_/Q _33771_/Q _36075_/Q _16671_/X _16672_/X VGND VGND VPWR
+ VPWR _16820_/X sky130_fd_sc_hd__mux4_1
X_29786_ _29786_/A VGND VGND VPWR VPWR _35152_/D sky130_fd_sc_hd__clkbuf_1
X_26998_ _33925_/Q _23444_/X _27002_/S VGND VGND VPWR VPWR _26999_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28737_ _34686_/Q _27158_/X _28755_/S VGND VGND VPWR VPWR _28738_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16751_ _32105_/Q _32297_/Q _32361_/Q _35881_/Q _16574_/X _16715_/X VGND VGND VPWR
+ VPWR _16751_/X sky130_fd_sc_hd__mux4_1
X_25949_ _24796_/X _33430_/Q _25967_/S VGND VGND VPWR VPWR _25950_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_1136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19470_ _34165_/Q _34101_/Q _34037_/Q _33973_/Q _19393_/X _19394_/X VGND VGND VPWR
+ VPWR _19470_/X sky130_fd_sc_hd__mux4_1
XFILLER_47_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28668_ _28668_/A VGND VGND VPWR VPWR _34653_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16682_ _16678_/X _16681_/X _16434_/X _16435_/X VGND VGND VPWR VPWR _16697_/B sky130_fd_sc_hd__o211a_1
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_235_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_1018 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18421_ _32855_/Q _32791_/Q _32727_/Q _32663_/Q _18337_/X _18339_/X VGND VGND VPWR
+ VPWR _18421_/X sky130_fd_sc_hd__mux4_1
XFILLER_74_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27619_ _34188_/Q _27202_/X _27629_/S VGND VGND VPWR VPWR _27620_/A sky130_fd_sc_hd__mux2_1
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28599_ _28599_/A VGND VGND VPWR VPWR _34621_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18352_ _20282_/A VGND VGND VPWR VPWR _20298_/A sky130_fd_sc_hd__buf_12
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30630_ _35552_/Q _29360_/X _30648_/S VGND VGND VPWR VPWR _30631_/A sky130_fd_sc_hd__mux2_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ _33657_/Q _33593_/Q _33529_/Q _33465_/Q _17200_/X _17201_/X VGND VGND VPWR
+ VPWR _17303_/X sky130_fd_sc_hd__mux4_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_875 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18283_ _18361_/A VGND VGND VPWR VPWR _20206_/A sky130_fd_sc_hd__buf_12
X_30561_ _30561_/A VGND VGND VPWR VPWR _35519_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_230_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_587 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32300_ _32875_/CLK _32300_/D VGND VGND VPWR VPWR _32300_/Q sky130_fd_sc_hd__dfxtp_1
X_17234_ _17228_/X _17233_/X _17165_/X VGND VGND VPWR VPWR _17235_/D sky130_fd_sc_hd__o21ba_1
X_33280_ _33921_/CLK _33280_/D VGND VGND VPWR VPWR _33280_/Q sky130_fd_sc_hd__dfxtp_1
X_30492_ _35487_/Q _29357_/X _30492_/S VGND VGND VPWR VPWR _30493_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32231_ _35124_/CLK _32231_/D VGND VGND VPWR VPWR _32231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17165_ _17871_/A VGND VGND VPWR VPWR _17165_/X sky130_fd_sc_hd__buf_2
XFILLER_127_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16116_ _16110_/X _16115_/X _16015_/X VGND VGND VPWR VPWR _16138_/A sky130_fd_sc_hd__o21ba_1
X_32162_ _36197_/CLK _32162_/D VGND VGND VPWR VPWR _32162_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17096_ _16846_/X _17092_/X _17095_/X _16851_/X VGND VGND VPWR VPWR _17096_/X sky130_fd_sc_hd__a22o_1
XFILLER_182_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31113_ _31113_/A VGND VGND VPWR VPWR _35781_/D sky130_fd_sc_hd__clkbuf_1
X_16047_ _16028_/X _16042_/X _16044_/X _16046_/X VGND VGND VPWR VPWR _16106_/B sky130_fd_sc_hd__o211a_1
XFILLER_100_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32093_ _32797_/CLK _32093_/D VGND VGND VPWR VPWR _32093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35921_ _35921_/CLK _35921_/D VGND VGND VPWR VPWR _35921_/Q sky130_fd_sc_hd__dfxtp_1
X_31044_ _31044_/A VGND VGND VPWR VPWR _35748_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19806_ _20159_/A VGND VGND VPWR VPWR _19806_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35852_ _35852_/CLK _35852_/D VGND VGND VPWR VPWR _35852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17998_ _17998_/A VGND VGND VPWR VPWR _17998_/X sky130_fd_sc_hd__buf_6
XFILLER_238_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34803_ _34927_/CLK _34803_/D VGND VGND VPWR VPWR _34803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19737_ _35196_/Q _35132_/Q _35068_/Q _32252_/Q _19663_/X _19664_/X VGND VGND VPWR
+ VPWR _19737_/X sky130_fd_sc_hd__mux4_1
XFILLER_211_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35783_ _35845_/CLK _35783_/D VGND VGND VPWR VPWR _35783_/Q sky130_fd_sc_hd__dfxtp_1
X_16949_ _16949_/A VGND VGND VPWR VPWR _31982_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32995_ _34593_/CLK _32995_/D VGND VGND VPWR VPWR _32995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34734_ _35183_/CLK _34734_/D VGND VGND VPWR VPWR _34734_/Q sky130_fd_sc_hd__dfxtp_1
X_31946_ _23481_/X _36176_/Q _31948_/S VGND VGND VPWR VPWR _31947_/A sky130_fd_sc_hd__mux2_1
X_19668_ _34938_/Q _34874_/Q _34810_/Q _34746_/Q _19460_/X _19461_/X VGND VGND VPWR
+ VPWR _19668_/X sky130_fd_sc_hd__mux4_1
XFILLER_25_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_1344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18619_ _20151_/A VGND VGND VPWR VPWR _18619_/X sky130_fd_sc_hd__buf_4
XFILLER_241_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34665_ _34913_/CLK _34665_/D VGND VGND VPWR VPWR _34665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19599_ _19458_/X _19597_/X _19598_/X _19463_/X VGND VGND VPWR VPWR _19599_/X sky130_fd_sc_hd__a22o_1
XFILLER_53_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31877_ _23316_/X _36143_/Q _31885_/S VGND VGND VPWR VPWR _31878_/A sky130_fd_sc_hd__mux2_1
X_33616_ _34192_/CLK _33616_/D VGND VGND VPWR VPWR _33616_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_6_39__f_CLK clkbuf_5_19_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_39__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_21630_ _33137_/Q _36017_/Q _33009_/Q _32945_/Q _21309_/X _21310_/X VGND VGND VPWR
+ VPWR _21630_/X sky130_fd_sc_hd__mux4_1
XFILLER_178_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30828_ _35646_/Q input35/X _30846_/S VGND VGND VPWR VPWR _30829_/A sky130_fd_sc_hd__mux2_1
X_34596_ _35490_/CLK _34596_/D VGND VGND VPWR VPWR _34596_/Q sky130_fd_sc_hd__dfxtp_1
X_33547_ _34188_/CLK _33547_/D VGND VGND VPWR VPWR _33547_/Q sky130_fd_sc_hd__dfxtp_1
X_21561_ _32879_/Q _32815_/Q _32751_/Q _32687_/Q _21240_/X _21241_/X VGND VGND VPWR
+ VPWR _21561_/X sky130_fd_sc_hd__mux4_1
X_30759_ _30759_/A VGND VGND VPWR VPWR _35613_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_1074 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23300_ _32172_/Q _23299_/X _23424_/S VGND VGND VPWR VPWR _23301_/A sky130_fd_sc_hd__mux2_1
X_20512_ _18348_/X _20510_/X _20511_/X _18358_/X VGND VGND VPWR VPWR _20512_/X sky130_fd_sc_hd__a22o_1
X_24280_ _24280_/A VGND VGND VPWR VPWR _32672_/D sky130_fd_sc_hd__clkbuf_1
X_33478_ _34179_/CLK _33478_/D VGND VGND VPWR VPWR _33478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21492_ _33133_/Q _36013_/Q _33005_/Q _32941_/Q _21309_/X _21310_/X VGND VGND VPWR
+ VPWR _21492_/X sky130_fd_sc_hd__mux4_1
XFILLER_53_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35217_ _35217_/CLK _35217_/D VGND VGND VPWR VPWR _35217_/Q sky130_fd_sc_hd__dfxtp_1
X_23231_ _23565_/S VGND VGND VPWR VPWR _23259_/S sky130_fd_sc_hd__buf_6
X_20443_ _35729_/Q _32240_/Q _35601_/Q _35537_/Q _18293_/X _18295_/X VGND VGND VPWR
+ VPWR _20443_/X sky130_fd_sc_hd__mux4_1
XFILLER_181_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32429_ _33895_/CLK _32429_/D VGND VGND VPWR VPWR _32429_/Q sky130_fd_sc_hd__dfxtp_1
X_36197_ _36197_/CLK _36197_/D VGND VGND VPWR VPWR _36197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35148_ _35213_/CLK _35148_/D VGND VGND VPWR VPWR _35148_/Q sky130_fd_sc_hd__dfxtp_1
X_23162_ _23162_/A VGND VGND VPWR VPWR _32119_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20374_ _20212_/X _20372_/X _20373_/X _20215_/X VGND VGND VPWR VPWR _20374_/X sky130_fd_sc_hd__a22o_1
XFILLER_109_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22113_ _22466_/A VGND VGND VPWR VPWR _22113_/X sky130_fd_sc_hd__buf_4
XTAP_7129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27970_ _27970_/A VGND VGND VPWR VPWR _34323_/D sky130_fd_sc_hd__clkbuf_1
X_23093_ _23093_/A VGND VGND VPWR VPWR _32086_/D sky130_fd_sc_hd__clkbuf_1
X_35079_ _35721_/CLK _35079_/D VGND VGND VPWR VPWR _35079_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26921_ _33888_/Q _23261_/X _26939_/S VGND VGND VPWR VPWR _26922_/A sky130_fd_sc_hd__mux2_1
X_22044_ _22044_/A VGND VGND VPWR VPWR _36220_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_248_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29640_ _35083_/Q _29494_/X _29652_/S VGND VGND VPWR VPWR _29641_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26852_ _26852_/A VGND VGND VPWR VPWR _33855_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25803_ _25803_/A VGND VGND VPWR VPWR _33361_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29571_ _35050_/Q _29391_/X _29589_/S VGND VGND VPWR VPWR _29572_/A sky130_fd_sc_hd__mux2_1
X_23995_ _23995_/A VGND VGND VPWR VPWR _32540_/D sky130_fd_sc_hd__clkbuf_1
X_26783_ _33823_/Q _23258_/X _26783_/S VGND VGND VPWR VPWR _26784_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28522_ _28522_/A VGND VGND VPWR VPWR _34584_/D sky130_fd_sc_hd__clkbuf_1
X_25734_ _25734_/A VGND VGND VPWR VPWR _33328_/D sky130_fd_sc_hd__clkbuf_1
X_22946_ input11/X VGND VGND VPWR VPWR _22946_/X sky130_fd_sc_hd__buf_2
XFILLER_244_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28453_ _27748_/X _34552_/Q _28463_/S VGND VGND VPWR VPWR _28454_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_245_1018 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25665_ _24979_/X _33296_/Q _25667_/S VGND VGND VPWR VPWR _25666_/A sky130_fd_sc_hd__mux2_1
X_22877_ _22877_/A _22877_/B _22877_/C _22877_/D VGND VGND VPWR VPWR _22878_/A sky130_fd_sc_hd__or4_4
XFILLER_186_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27404_ _34086_/Q _27084_/X _27410_/S VGND VGND VPWR VPWR _27405_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24616_ _23018_/X _32832_/Q _24630_/S VGND VGND VPWR VPWR _24617_/A sky130_fd_sc_hd__mux2_1
X_21828_ _21753_/X _21826_/X _21827_/X _21756_/X VGND VGND VPWR VPWR _21828_/X sky130_fd_sc_hd__a22o_1
X_28384_ _27646_/X _34519_/Q _28400_/S VGND VGND VPWR VPWR _28385_/A sky130_fd_sc_hd__mux2_1
X_25596_ _24877_/X _33263_/Q _25604_/S VGND VGND VPWR VPWR _25597_/A sky130_fd_sc_hd__mux2_1
XFILLER_227_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27335_ _27335_/A VGND VGND VPWR VPWR _34053_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24547_ _24547_/A VGND VGND VPWR VPWR _32799_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21759_ _34420_/Q _36148_/Q _34292_/Q _34228_/Q _21476_/X _21477_/X VGND VGND VPWR
+ VPWR _21759_/X sky130_fd_sc_hd__mux4_1
XFILLER_19_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24478_ _24478_/A VGND VGND VPWR VPWR _32766_/D sky130_fd_sc_hd__clkbuf_1
X_27266_ _27266_/A VGND VGND VPWR VPWR _34020_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29005_ _29005_/A VGND VGND VPWR VPWR _34812_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23429_ input37/X VGND VGND VPWR VPWR _23429_/X sky130_fd_sc_hd__buf_4
X_26217_ _31553_/A _26352_/B VGND VGND VPWR VPWR _26350_/S sky130_fd_sc_hd__nand2_8
X_27197_ _33994_/Q _27196_/X _27218_/S VGND VGND VPWR VPWR _27198_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26148_ _26148_/A VGND VGND VPWR VPWR _33524_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26079_ _26079_/A VGND VGND VPWR VPWR _33492_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18970_ _33383_/Q _33319_/Q _33255_/Q _33191_/Q _18721_/X _18722_/X VGND VGND VPWR
+ VPWR _18970_/X sky130_fd_sc_hd__mux4_1
XFILLER_98_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_700 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29907_ _29907_/A VGND VGND VPWR VPWR _35209_/D sky130_fd_sc_hd__clkbuf_1
X_17921_ _32138_/Q _32330_/Q _32394_/Q _35914_/Q _17633_/X _17774_/X VGND VGND VPWR
+ VPWR _17921_/X sky130_fd_sc_hd__mux4_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17852_ _35656_/Q _35016_/Q _34376_/Q _33736_/Q _17850_/X _17851_/X VGND VGND VPWR
+ VPWR _17852_/X sky130_fd_sc_hd__mux4_1
X_29838_ _35177_/Q _29388_/X _29838_/S VGND VGND VPWR VPWR _29839_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16803_ _17156_/A VGND VGND VPWR VPWR _16803_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_120_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29769_ _35144_/Q _29484_/X _29787_/S VGND VGND VPWR VPWR _29770_/A sky130_fd_sc_hd__mux2_1
X_17783_ _35462_/Q _35398_/Q _35334_/Q _35270_/Q _17607_/X _17608_/X VGND VGND VPWR
+ VPWR _17783_/X sky130_fd_sc_hd__mux4_1
XFILLER_130_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31800_ _31800_/A VGND VGND VPWR VPWR _36106_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_219_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19522_ _35446_/Q _35382_/Q _35318_/Q _35254_/Q _19201_/X _19202_/X VGND VGND VPWR
+ VPWR _19522_/X sky130_fd_sc_hd__mux4_1
X_16734_ _34920_/Q _34856_/Q _34792_/Q _34728_/Q _16454_/X _16455_/X VGND VGND VPWR
+ VPWR _16734_/X sky130_fd_sc_hd__mux4_1
XFILLER_93_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32780_ _32879_/CLK _32780_/D VGND VGND VPWR VPWR _32780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31731_ _31821_/S VGND VGND VPWR VPWR _31750_/S sky130_fd_sc_hd__buf_4
X_19453_ _19453_/A VGND VGND VPWR VPWR _19453_/X sky130_fd_sc_hd__clkbuf_4
X_16665_ _16665_/A _16665_/B _16665_/C _16665_/D VGND VGND VPWR VPWR _16666_/A sky130_fd_sc_hd__or4_2
XFILLER_61_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18404_ _20171_/A VGND VGND VPWR VPWR _18404_/X sky130_fd_sc_hd__clkbuf_4
X_34450_ _36180_/CLK _34450_/D VGND VGND VPWR VPWR _34450_/Q sky130_fd_sc_hd__dfxtp_1
X_31662_ _27801_/X _36041_/Q _31678_/S VGND VGND VPWR VPWR _31663_/A sky130_fd_sc_hd__mux2_1
X_19384_ _35186_/Q _35122_/Q _35058_/Q _32209_/Q _19310_/X _19311_/X VGND VGND VPWR
+ VPWR _19384_/X sky130_fd_sc_hd__mux4_1
X_16596_ _16596_/A VGND VGND VPWR VPWR _31972_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33401_ _33914_/CLK _33401_/D VGND VGND VPWR VPWR _33401_/Q sky130_fd_sc_hd__dfxtp_1
X_30613_ _35544_/Q _29336_/X _30627_/S VGND VGND VPWR VPWR _30614_/A sky130_fd_sc_hd__mux2_1
X_18335_ _32086_/Q _32278_/Q _32342_/Q _35862_/Q _18332_/X _20167_/A VGND VGND VPWR
+ VPWR _18335_/X sky130_fd_sc_hd__mux4_1
XFILLER_128_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34381_ _35663_/CLK _34381_/D VGND VGND VPWR VPWR _34381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31593_ _31593_/A VGND VGND VPWR VPWR _36008_/D sky130_fd_sc_hd__clkbuf_1
X_36120_ _36121_/CLK _36120_/D VGND VGND VPWR VPWR _36120_/Q sky130_fd_sc_hd__dfxtp_1
X_33332_ _34100_/CLK _33332_/D VGND VGND VPWR VPWR _33332_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18266_ _35477_/Q _35413_/Q _35349_/Q _35285_/Q _16009_/X _16011_/X VGND VGND VPWR
+ VPWR _18266_/X sky130_fd_sc_hd__mux4_1
X_30544_ _30544_/A VGND VGND VPWR VPWR _35511_/D sky130_fd_sc_hd__clkbuf_1
X_36051_ _36051_/CLK _36051_/D VGND VGND VPWR VPWR _36051_/Q sky130_fd_sc_hd__dfxtp_1
X_17217_ _17067_/X _17215_/X _17216_/X _17071_/X VGND VGND VPWR VPWR _17217_/X sky130_fd_sc_hd__a22o_1
XFILLER_198_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33263_ _36079_/CLK _33263_/D VGND VGND VPWR VPWR _33263_/Q sky130_fd_sc_hd__dfxtp_1
X_30475_ _30475_/A VGND VGND VPWR VPWR _35478_/D sky130_fd_sc_hd__clkbuf_1
X_18197_ _33171_/Q _36051_/Q _33043_/Q _32979_/Q _16032_/X _17161_/A VGND VGND VPWR
+ VPWR _18197_/X sky130_fd_sc_hd__mux4_1
X_35002_ _35645_/CLK _35002_/D VGND VGND VPWR VPWR _35002_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32214_ _35835_/CLK _32214_/D VGND VGND VPWR VPWR _32214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17148_ _35444_/Q _35380_/Q _35316_/Q _35252_/Q _16901_/X _16902_/X VGND VGND VPWR
+ VPWR _17148_/X sky130_fd_sc_hd__mux4_1
X_33194_ _34091_/CLK _33194_/D VGND VGND VPWR VPWR _33194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32145_ _32913_/CLK _32145_/D VGND VGND VPWR VPWR _32145_/Q sky130_fd_sc_hd__dfxtp_1
X_17079_ _17936_/A VGND VGND VPWR VPWR _17079_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_171_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20090_ _35206_/Q _35142_/Q _35078_/Q _32262_/Q _20016_/X _20017_/X VGND VGND VPWR
+ VPWR _20090_/X sky130_fd_sc_hd__mux4_1
XFILLER_170_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32076_ _36042_/CLK _32076_/D VGND VGND VPWR VPWR _32076_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31027_ _31027_/A VGND VGND VPWR VPWR _35740_/D sky130_fd_sc_hd__clkbuf_1
X_35904_ _35969_/CLK _35904_/D VGND VGND VPWR VPWR _35904_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_1387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35835_ _35835_/CLK _35835_/D VGND VGND VPWR VPWR _35835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22800_ _32915_/Q _32851_/Q _32787_/Q _32723_/Q _20584_/X _20587_/X VGND VGND VPWR
+ VPWR _22800_/X sky130_fd_sc_hd__mux4_1
XFILLER_84_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23780_ _22993_/X _32376_/Q _23790_/S VGND VGND VPWR VPWR _23781_/A sky130_fd_sc_hd__mux2_1
X_32978_ _35858_/CLK _32978_/D VGND VGND VPWR VPWR _32978_/Q sky130_fd_sc_hd__dfxtp_1
X_20992_ _33887_/Q _33823_/Q _33759_/Q _36063_/Q _20918_/X _20919_/X VGND VGND VPWR
+ VPWR _20992_/X sky130_fd_sc_hd__mux4_1
X_35766_ _35830_/CLK _35766_/D VGND VGND VPWR VPWR _35766_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22731_ _22505_/X _22729_/X _22730_/X _22510_/X VGND VGND VPWR VPWR _22731_/X sky130_fd_sc_hd__a22o_1
X_34717_ _36242_/CLK _34717_/D VGND VGND VPWR VPWR _34717_/Q sky130_fd_sc_hd__dfxtp_1
X_31929_ _31956_/S VGND VGND VPWR VPWR _31948_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_129_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35697_ _35697_/CLK _35697_/D VGND VGND VPWR VPWR _35697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25450_ _25540_/S VGND VGND VPWR VPWR _25469_/S sky130_fd_sc_hd__buf_4
XFILLER_53_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34648_ _34903_/CLK _34648_/D VGND VGND VPWR VPWR _34648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22662_ _22459_/X _22660_/X _22661_/X _22462_/X VGND VGND VPWR VPWR _22662_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24401_ _22900_/X _32730_/Q _24411_/S VGND VGND VPWR VPWR _24402_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21613_ _21400_/X _21609_/X _21612_/X _21403_/X VGND VGND VPWR VPWR _21613_/X sky130_fd_sc_hd__a22o_1
XFILLER_197_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25381_ _33162_/Q _23463_/X _25395_/S VGND VGND VPWR VPWR _25382_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_222_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34579_ _34708_/CLK _34579_/D VGND VGND VPWR VPWR _34579_/Q sky130_fd_sc_hd__dfxtp_1
X_22593_ _22304_/X _22591_/X _22592_/X _22307_/X VGND VGND VPWR VPWR _22593_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_1434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27120_ _27120_/A VGND VGND VPWR VPWR _33969_/D sky130_fd_sc_hd__clkbuf_1
X_24332_ _24332_/A VGND VGND VPWR VPWR _32697_/D sky130_fd_sc_hd__clkbuf_1
X_21544_ _34414_/Q _36142_/Q _34286_/Q _34222_/Q _21476_/X _21477_/X VGND VGND VPWR
+ VPWR _21544_/X sky130_fd_sc_hd__mux4_1
X_27051_ _33947_/Q _27050_/X _27063_/S VGND VGND VPWR VPWR _27052_/A sky130_fd_sc_hd__mux2_1
X_24263_ _24263_/A VGND VGND VPWR VPWR _32664_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21475_ _21400_/X _21473_/X _21474_/X _21403_/X VGND VGND VPWR VPWR _21475_/X sky130_fd_sc_hd__a22o_1
XFILLER_217_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26002_ _26002_/A VGND VGND VPWR VPWR _33455_/D sky130_fd_sc_hd__clkbuf_1
X_23214_ _23214_/A VGND VGND VPWR VPWR _32144_/D sky130_fd_sc_hd__clkbuf_1
X_20426_ _20422_/X _20425_/X _20171_/X VGND VGND VPWR VPWR _20427_/D sky130_fd_sc_hd__o21ba_1
X_24194_ _24194_/A VGND VGND VPWR VPWR _32633_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23145_ _23145_/A VGND VGND VPWR VPWR _32111_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20357_ _33102_/Q _32078_/Q _35854_/Q _35790_/Q _20084_/X _20085_/X VGND VGND VPWR
+ VPWR _20357_/X sky130_fd_sc_hd__mux4_1
XFILLER_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27953_ _27807_/X _34315_/Q _27965_/S VGND VGND VPWR VPWR _27954_/A sky130_fd_sc_hd__mux2_1
XFILLER_216_1120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23076_ input58/X VGND VGND VPWR VPWR _23076_/X sky130_fd_sc_hd__clkbuf_2
XTAP_6236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20288_ _32908_/Q _32844_/Q _32780_/Q _32716_/Q _19999_/X _20000_/X VGND VGND VPWR
+ VPWR _20288_/X sky130_fd_sc_hd__mux4_1
XTAP_5502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26904_ _33880_/Q _23237_/X _26918_/S VGND VGND VPWR VPWR _26905_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22027_ _35708_/Q _32217_/Q _35580_/Q _35516_/Q _21917_/X _21918_/X VGND VGND VPWR
+ VPWR _22027_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_130_CLK clkbuf_6_23__f_CLK/X VGND VGND VPWR VPWR _35160_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_6269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27884_ _27704_/X _34282_/Q _27902_/S VGND VGND VPWR VPWR _27885_/A sky130_fd_sc_hd__mux2_1
XTAP_5546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29623_ _35075_/Q _29469_/X _29631_/S VGND VGND VPWR VPWR _29624_/A sky130_fd_sc_hd__mux2_1
XTAP_5568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26835_ _26835_/A VGND VGND VPWR VPWR _33847_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29554_ _35042_/Q _29367_/X _29568_/S VGND VGND VPWR VPWR _29555_/A sky130_fd_sc_hd__mux2_1
XTAP_4878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26766_ _26766_/A VGND VGND VPWR VPWR _33814_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23978_ _23978_/A VGND VGND VPWR VPWR _32533_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28505_ _27825_/X _34577_/Q _28505_/S VGND VGND VPWR VPWR _28506_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25717_ _25717_/A VGND VGND VPWR VPWR _33320_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29485_ _29525_/S VGND VGND VPWR VPWR _29513_/S sky130_fd_sc_hd__buf_4
XFILLER_16_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22929_ _22928_/X _32035_/Q _22947_/S VGND VGND VPWR VPWR _22930_/A sky130_fd_sc_hd__mux2_1
XFILLER_232_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26697_ _33782_/Q _23396_/X _26711_/S VGND VGND VPWR VPWR _26698_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28436_ _27723_/X _34544_/Q _28442_/S VGND VGND VPWR VPWR _28437_/A sky130_fd_sc_hd__mux2_1
X_16450_ _17156_/A VGND VGND VPWR VPWR _16450_/X sky130_fd_sc_hd__buf_4
X_25648_ _25675_/S VGND VGND VPWR VPWR _25667_/S sky130_fd_sc_hd__buf_4
XFILLER_182_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16381_ _34910_/Q _34846_/Q _34782_/Q _34718_/Q _16096_/X _16098_/X VGND VGND VPWR
+ VPWR _16381_/X sky130_fd_sc_hd__mux4_1
X_28367_ _28367_/A VGND VGND VPWR VPWR _34511_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_22__f_CLK clkbuf_5_11_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_22__f_CLK/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_197_CLK clkbuf_6_49__f_CLK/X VGND VGND VPWR VPWR _35727_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25579_ _24852_/X _33255_/Q _25583_/S VGND VGND VPWR VPWR _25580_/A sky130_fd_sc_hd__mux2_1
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18120_ _34704_/Q _34640_/Q _34576_/Q _34512_/Q _17998_/X _17999_/X VGND VGND VPWR
+ VPWR _18120_/X sky130_fd_sc_hd__mux4_1
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27318_ _27318_/A VGND VGND VPWR VPWR _34045_/D sky130_fd_sc_hd__clkbuf_1
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28298_ _28298_/A VGND VGND VPWR VPWR _34478_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18051_ _17773_/X _18049_/X _18050_/X _17777_/X VGND VGND VPWR VPWR _18051_/X sky130_fd_sc_hd__a22o_1
XFILLER_200_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27249_ _27249_/A VGND VGND VPWR VPWR _34012_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_240_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17002_ _16998_/X _16999_/X _17000_/X _17001_/X VGND VGND VPWR VPWR _17002_/X sky130_fd_sc_hd__a22o_1
XFILLER_126_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30260_ _35377_/Q _29413_/X _30264_/S VGND VGND VPWR VPWR _30261_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30191_ _30191_/A VGND VGND VPWR VPWR _35344_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18953_ _20169_/A VGND VGND VPWR VPWR _18953_/X sky130_fd_sc_hd__buf_4
XFILLER_193_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17904_ _17904_/A VGND VGND VPWR VPWR _32009_/D sky130_fd_sc_hd__clkbuf_4
X_33950_ _36188_/CLK _33950_/D VGND VGND VPWR VPWR _33950_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_121_CLK clkbuf_6_21__f_CLK/X VGND VGND VPWR VPWR _36127_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_121_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18884_ _18597_/X _18882_/X _18883_/X _18600_/X VGND VGND VPWR VPWR _18884_/X sky130_fd_sc_hd__a22o_1
XTAP_6770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32901_ _32901_/CLK _32901_/D VGND VGND VPWR VPWR _32901_/Q sky130_fd_sc_hd__dfxtp_1
X_17835_ _33416_/Q _33352_/Q _33288_/Q _33224_/Q _17833_/X _17834_/X VGND VGND VPWR
+ VPWR _17835_/X sky130_fd_sc_hd__mux4_1
XTAP_6792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33881_ _34009_/CLK _33881_/D VGND VGND VPWR VPWR _33881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32832_ _32896_/CLK _32832_/D VGND VGND VPWR VPWR _32832_/Q sky130_fd_sc_hd__dfxtp_1
X_35620_ _35620_/CLK _35620_/D VGND VGND VPWR VPWR _35620_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17766_ _17766_/A VGND VGND VPWR VPWR _17766_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_47_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19505_ _19499_/X _19502_/X _19503_/X _19504_/X VGND VGND VPWR VPWR _19505_/X sky130_fd_sc_hd__a22o_1
XFILLER_235_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35551_ _35551_/CLK _35551_/D VGND VGND VPWR VPWR _35551_/Q sky130_fd_sc_hd__dfxtp_1
X_16717_ _32872_/Q _32808_/Q _32744_/Q _32680_/Q _16640_/X _16641_/X VGND VGND VPWR
+ VPWR _16717_/X sky130_fd_sc_hd__mux4_1
X_32763_ _32891_/CLK _32763_/D VGND VGND VPWR VPWR _32763_/Q sky130_fd_sc_hd__dfxtp_1
X_17697_ _17412_/X _17695_/X _17696_/X _17418_/X VGND VGND VPWR VPWR _17697_/X sky130_fd_sc_hd__a22o_1
XFILLER_35_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34502_ _35657_/CLK _34502_/D VGND VGND VPWR VPWR _34502_/Q sky130_fd_sc_hd__dfxtp_1
X_31714_ _31714_/A VGND VGND VPWR VPWR _36065_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_986 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19436_ _19359_/X _19434_/X _19435_/X _19365_/X VGND VGND VPWR VPWR _19436_/X sky130_fd_sc_hd__a22o_1
X_35482_ _35482_/CLK _35482_/D VGND VGND VPWR VPWR _35482_/Q sky130_fd_sc_hd__dfxtp_1
X_16648_ _17862_/A VGND VGND VPWR VPWR _16648_/X sky130_fd_sc_hd__clkbuf_4
X_32694_ _32903_/CLK _32694_/D VGND VGND VPWR VPWR _32694_/Q sky130_fd_sc_hd__dfxtp_1
X_34433_ _34690_/CLK _34433_/D VGND VGND VPWR VPWR _34433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31645_ _27776_/X _36033_/Q _31657_/S VGND VGND VPWR VPWR _31646_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_188_CLK clkbuf_leaf_65_CLK/A VGND VGND VPWR VPWR _35982_/CLK sky130_fd_sc_hd__clkbuf_16
X_19367_ _20212_/A VGND VGND VPWR VPWR _19367_/X sky130_fd_sc_hd__clkbuf_4
X_16579_ _35684_/Q _32191_/Q _35556_/Q _35492_/Q _16258_/X _16259_/X VGND VGND VPWR
+ VPWR _16579_/X sky130_fd_sc_hd__mux4_1
XFILLER_128_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18318_ _20205_/A VGND VGND VPWR VPWR _18318_/X sky130_fd_sc_hd__buf_4
X_34364_ _35644_/CLK _34364_/D VGND VGND VPWR VPWR _34364_/Q sky130_fd_sc_hd__dfxtp_1
X_31576_ _27673_/X _36000_/Q _31594_/S VGND VGND VPWR VPWR _31577_/A sky130_fd_sc_hd__mux2_1
X_19298_ _20159_/A VGND VGND VPWR VPWR _19298_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_148_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36103_ _36103_/CLK _36103_/D VGND VGND VPWR VPWR _36103_/Q sky130_fd_sc_hd__dfxtp_1
X_33315_ _33573_/CLK _33315_/D VGND VGND VPWR VPWR _33315_/Q sky130_fd_sc_hd__dfxtp_1
X_18249_ _33685_/Q _33621_/Q _33557_/Q _33493_/Q _16024_/X _16025_/X VGND VGND VPWR
+ VPWR _18249_/X sky130_fd_sc_hd__mux4_1
X_30527_ _30527_/A VGND VGND VPWR VPWR _35503_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34295_ _36150_/CLK _34295_/D VGND VGND VPWR VPWR _34295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36034_ _36034_/CLK _36034_/D VGND VGND VPWR VPWR _36034_/Q sky130_fd_sc_hd__dfxtp_1
X_33246_ _36191_/CLK _33246_/D VGND VGND VPWR VPWR _33246_/Q sky130_fd_sc_hd__dfxtp_1
X_21260_ _21047_/X _21256_/X _21259_/X _21050_/X VGND VGND VPWR VPWR _21260_/X sky130_fd_sc_hd__a22o_1
X_30458_ _35471_/Q _29506_/X _30462_/S VGND VGND VPWR VPWR _30459_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20211_ _20205_/X _20208_/X _20209_/X _20210_/X VGND VGND VPWR VPWR _20211_/X sky130_fd_sc_hd__a22o_1
XFILLER_117_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33177_ _33753_/CLK _33177_/D VGND VGND VPWR VPWR _33177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21191_ _34404_/Q _36132_/Q _34276_/Q _34212_/Q _21123_/X _21124_/X VGND VGND VPWR
+ VPWR _21191_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_360_CLK clkbuf_6_46__f_CLK/X VGND VGND VPWR VPWR _35577_/CLK sky130_fd_sc_hd__clkbuf_16
X_30389_ _35438_/Q _29404_/X _30399_/S VGND VGND VPWR VPWR _30390_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20142_ _20065_/X _20140_/X _20141_/X _20071_/X VGND VGND VPWR VPWR _20142_/X sky130_fd_sc_hd__a22o_1
X_32128_ _35969_/CLK _32128_/D VGND VGND VPWR VPWR _32128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_1140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_112_CLK clkbuf_6_22__f_CLK/X VGND VGND VPWR VPWR _35673_/CLK sky130_fd_sc_hd__clkbuf_16
X_24950_ _24950_/A VGND VGND VPWR VPWR _32966_/D sky130_fd_sc_hd__clkbuf_1
X_20073_ _20073_/A VGND VGND VPWR VPWR _20073_/X sky130_fd_sc_hd__clkbuf_4
X_32059_ _35835_/CLK _32059_/D VGND VGND VPWR VPWR _32059_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23901_ _23901_/A VGND VGND VPWR VPWR _32496_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_245_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_246_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24881_ _24880_/X _32944_/Q _24890_/S VGND VGND VPWR VPWR _24882_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26620_ _24991_/X _33748_/Q _26622_/S VGND VGND VPWR VPWR _26621_/A sky130_fd_sc_hd__mux2_1
XTAP_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23832_ _23070_/X _32401_/Q _23832_/S VGND VGND VPWR VPWR _23833_/A sky130_fd_sc_hd__mux2_1
X_35818_ _35820_/CLK _35818_/D VGND VGND VPWR VPWR _35818_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_14_0_CLK clkbuf_5_9_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_14_0_CLK/X sky130_fd_sc_hd__clkbuf_8
X_26551_ _24889_/X _33715_/Q _26551_/S VGND VGND VPWR VPWR _26552_/A sky130_fd_sc_hd__mux2_1
X_23763_ _22968_/X _32368_/Q _23769_/S VGND VGND VPWR VPWR _23764_/A sky130_fd_sc_hd__mux2_1
X_20975_ _20897_/X _20971_/X _20974_/X _20900_/X VGND VGND VPWR VPWR _20975_/X sky130_fd_sc_hd__a22o_1
X_35749_ _35814_/CLK _35749_/D VGND VGND VPWR VPWR _35749_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25502_ _25502_/A VGND VGND VPWR VPWR _33218_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22714_ _35664_/Q _35024_/Q _34384_/Q _33744_/Q _22450_/X _22451_/X VGND VGND VPWR
+ VPWR _22714_/X sky130_fd_sc_hd__mux4_1
X_29270_ _34938_/Q _27146_/X _29276_/S VGND VGND VPWR VPWR _29271_/A sky130_fd_sc_hd__mux2_1
X_26482_ _33683_/Q _23492_/X _26486_/S VGND VGND VPWR VPWR _26483_/A sky130_fd_sc_hd__mux2_1
XFILLER_214_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23694_ _23070_/X _32337_/Q _23694_/S VGND VGND VPWR VPWR _23695_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28221_ _27804_/X _34442_/Q _28235_/S VGND VGND VPWR VPWR _28222_/A sky130_fd_sc_hd__mux2_1
XFILLER_214_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22645_ _22641_/X _22644_/X _22438_/X VGND VGND VPWR VPWR _22667_/A sky130_fd_sc_hd__o21ba_1
XFILLER_201_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25433_ _25433_/A VGND VGND VPWR VPWR _33185_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_179_CLK clkbuf_6_27__f_CLK/X VGND VGND VPWR VPWR _35026_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_213_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_5_29_0_CLK clkbuf_2_3_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_29_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_185_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25364_ _33154_/Q _23435_/X _25374_/S VGND VGND VPWR VPWR _25365_/A sky130_fd_sc_hd__mux2_1
X_28152_ _28152_/A VGND VGND VPWR VPWR _34409_/D sky130_fd_sc_hd__clkbuf_1
X_22576_ _34188_/Q _34124_/Q _34060_/Q _33996_/Q _22399_/X _22400_/X VGND VGND VPWR
+ VPWR _22576_/X sky130_fd_sc_hd__mux4_1
XFILLER_167_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27103_ input15/X VGND VGND VPWR VPWR _27103_/X sky130_fd_sc_hd__buf_2
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21527_ _22586_/A VGND VGND VPWR VPWR _21527_/X sky130_fd_sc_hd__buf_6
X_24315_ _24315_/A VGND VGND VPWR VPWR _32689_/D sky130_fd_sc_hd__clkbuf_1
X_28083_ _28083_/A VGND VGND VPWR VPWR _34376_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25295_ _33121_/Q _23265_/X _25311_/S VGND VGND VPWR VPWR _25296_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27034_ _30472_/A _31688_/B VGND VGND VPWR VPWR _27230_/S sky130_fd_sc_hd__nor2_8
X_24246_ _24246_/A VGND VGND VPWR VPWR _32658_/D sky130_fd_sc_hd__clkbuf_1
X_21458_ _21452_/X _21457_/X _21379_/X VGND VGND VPWR VPWR _21482_/A sky130_fd_sc_hd__o21ba_1
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20409_ _32144_/Q _32336_/Q _32400_/Q _35920_/Q _20286_/X _19311_/A VGND VGND VPWR
+ VPWR _20409_/X sky130_fd_sc_hd__mux4_1
X_24177_ _24177_/A VGND VGND VPWR VPWR _32625_/D sky130_fd_sc_hd__clkbuf_1
X_21389_ _21383_/X _21386_/X _21387_/X _21388_/X VGND VGND VPWR VPWR _21414_/B sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_351_CLK clkbuf_6_47__f_CLK/X VGND VGND VPWR VPWR _35708_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_162_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23128_ _23128_/A VGND VGND VPWR VPWR _32103_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28985_ _34803_/Q _27124_/X _28985_/S VGND VGND VPWR VPWR _28986_/A sky130_fd_sc_hd__mux2_1
XTAP_6022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27936_ _27782_/X _34307_/Q _27944_/S VGND VGND VPWR VPWR _27937_/A sky130_fd_sc_hd__mux2_1
XTAP_5310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_103_CLK clkbuf_leaf_99_CLK/A VGND VGND VPWR VPWR _34331_/CLK sky130_fd_sc_hd__clkbuf_16
X_23059_ _23058_/X _32077_/Q _23071_/S VGND VGND VPWR VPWR _23060_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput98 _31975_/Q VGND VGND VPWR VPWR D1[17] sky130_fd_sc_hd__buf_2
XTAP_6066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27867_ _27680_/X _34274_/Q _27881_/S VGND VGND VPWR VPWR _27868_/A sky130_fd_sc_hd__mux2_1
XTAP_5376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17620_ _17620_/A _17620_/B _17620_/C _17620_/D VGND VGND VPWR VPWR _17621_/A sky130_fd_sc_hd__or4_1
XTAP_4642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29606_ _35067_/Q _29444_/X _29610_/S VGND VGND VPWR VPWR _29607_/A sky130_fd_sc_hd__mux2_1
XTAP_5398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26818_ _26818_/A VGND VGND VPWR VPWR _33839_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27798_ _27838_/S VGND VGND VPWR VPWR _27826_/S sky130_fd_sc_hd__buf_4
XTAP_4675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29537_ _35034_/Q _29342_/X _29547_/S VGND VGND VPWR VPWR _29538_/A sky130_fd_sc_hd__mux2_1
XTAP_4697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17551_ _17551_/A VGND VGND VPWR VPWR _31999_/D sky130_fd_sc_hd__buf_4
XFILLER_16_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26749_ _33807_/Q _23478_/X _26753_/S VGND VGND VPWR VPWR _26750_/A sky130_fd_sc_hd__mux2_1
XTAP_3963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16502_ _33890_/Q _33826_/Q _33762_/Q _36066_/Q _16318_/X _16319_/X VGND VGND VPWR
+ VPWR _16502_/X sky130_fd_sc_hd__mux4_1
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29468_ _29468_/A VGND VGND VPWR VPWR _35010_/D sky130_fd_sc_hd__clkbuf_1
X_17482_ _33406_/Q _33342_/Q _33278_/Q _33214_/Q _17480_/X _17481_/X VGND VGND VPWR
+ VPWR _17482_/X sky130_fd_sc_hd__mux4_1
XFILLER_189_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19221_ _19153_/X _19219_/X _19220_/X _19156_/X VGND VGND VPWR VPWR _19221_/X sky130_fd_sc_hd__a22o_1
X_16433_ _16361_/X _16431_/X _16432_/X _16365_/X VGND VGND VPWR VPWR _16433_/X sky130_fd_sc_hd__a22o_1
X_28419_ _27698_/X _34536_/Q _28421_/S VGND VGND VPWR VPWR _28420_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29399_ _34988_/Q _29398_/X _29420_/S VGND VGND VPWR VPWR _29400_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31430_ _27658_/X _35931_/Q _31438_/S VGND VGND VPWR VPWR _31431_/A sky130_fd_sc_hd__mux2_1
X_19152_ _19146_/X _19149_/X _19150_/X _19151_/X VGND VGND VPWR VPWR _19152_/X sky130_fd_sc_hd__a22o_1
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16364_ _32862_/Q _32798_/Q _32734_/Q _32670_/Q _16287_/X _16288_/X VGND VGND VPWR
+ VPWR _16364_/X sky130_fd_sc_hd__mux4_1
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18103_ _33936_/Q _33872_/Q _33808_/Q _36112_/Q _16062_/X _16064_/X VGND VGND VPWR
+ VPWR _18103_/X sky130_fd_sc_hd__mux4_1
XFILLER_200_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19083_ _19006_/X _19081_/X _19082_/X _19012_/X VGND VGND VPWR VPWR _19083_/X sky130_fd_sc_hd__a22o_1
X_31361_ _31361_/A VGND VGND VPWR VPWR _35898_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16295_ _17862_/A VGND VGND VPWR VPWR _16295_/X sky130_fd_sc_hd__buf_4
XFILLER_201_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33100_ _35852_/CLK _33100_/D VGND VGND VPWR VPWR _33100_/Q sky130_fd_sc_hd__dfxtp_1
X_18034_ _34957_/Q _34893_/Q _34829_/Q _34765_/Q _17866_/X _17867_/X VGND VGND VPWR
+ VPWR _18034_/X sky130_fd_sc_hd__mux4_1
X_30312_ _30312_/A VGND VGND VPWR VPWR _35401_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_1252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34080_ _36202_/CLK _34080_/D VGND VGND VPWR VPWR _34080_/Q sky130_fd_sc_hd__dfxtp_1
X_31292_ _31292_/A VGND VGND VPWR VPWR _35865_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33031_ _33160_/CLK _33031_/D VGND VGND VPWR VPWR _33031_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30243_ _35369_/Q _29388_/X _30243_/S VGND VGND VPWR VPWR _30244_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_342_CLK clkbuf_6_45__f_CLK/X VGND VGND VPWR VPWR _32896_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_114_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19985_ _19981_/X _19984_/X _19818_/X VGND VGND VPWR VPWR _19986_/D sky130_fd_sc_hd__o21ba_1
X_30174_ _35336_/Q _29484_/X _30192_/S VGND VGND VPWR VPWR _30175_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18936_ _32614_/Q _32550_/Q _32486_/Q _35942_/Q _18870_/X _18654_/X VGND VGND VPWR
+ VPWR _18936_/X sky130_fd_sc_hd__mux4_1
XFILLER_132_1302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34982_ _35559_/CLK _34982_/D VGND VGND VPWR VPWR _34982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33933_ _36109_/CLK _33933_/D VGND VGND VPWR VPWR _33933_/Q sky130_fd_sc_hd__dfxtp_1
X_18867_ _33892_/Q _33828_/Q _33764_/Q _36068_/Q _18618_/X _18619_/X VGND VGND VPWR
+ VPWR _18867_/X sky130_fd_sc_hd__mux4_1
XFILLER_41_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17818_ _33095_/Q _32071_/Q _35847_/Q _35783_/Q _17784_/X _17785_/X VGND VGND VPWR
+ VPWR _17818_/X sky130_fd_sc_hd__mux4_1
X_33864_ _36104_/CLK _33864_/D VGND VGND VPWR VPWR _33864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_212_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_1379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18798_ _20162_/A VGND VGND VPWR VPWR _18798_/X sky130_fd_sc_hd__buf_4
XFILLER_167_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35603_ _35730_/CLK _35603_/D VGND VGND VPWR VPWR _35603_/Q sky130_fd_sc_hd__dfxtp_1
X_32815_ _32879_/CLK _32815_/D VGND VGND VPWR VPWR _32815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17749_ _34693_/Q _34629_/Q _34565_/Q _34501_/Q _17645_/X _17646_/X VGND VGND VPWR
+ VPWR _17749_/X sky130_fd_sc_hd__mux4_1
XFILLER_208_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33795_ _36100_/CLK _33795_/D VGND VGND VPWR VPWR _33795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20760_ _35672_/Q _32178_/Q _35544_/Q _35480_/Q _20649_/X _20650_/X VGND VGND VPWR
+ VPWR _20760_/X sky130_fd_sc_hd__mux4_1
X_35534_ _35599_/CLK _35534_/D VGND VGND VPWR VPWR _35534_/Q sky130_fd_sc_hd__dfxtp_1
X_32746_ _32875_/CLK _32746_/D VGND VGND VPWR VPWR _32746_/Q sky130_fd_sc_hd__dfxtp_1
X_19419_ _34931_/Q _34867_/Q _34803_/Q _34739_/Q _19107_/X _19108_/X VGND VGND VPWR
+ VPWR _19419_/X sky130_fd_sc_hd__mux4_1
X_35465_ _35721_/CLK _35465_/D VGND VGND VPWR VPWR _35465_/Q sky130_fd_sc_hd__dfxtp_1
X_20691_ _21758_/A VGND VGND VPWR VPWR _20691_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_195_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32677_ _32869_/CLK _32677_/D VGND VGND VPWR VPWR _32677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22430_ _33672_/Q _33608_/Q _33544_/Q _33480_/Q _22153_/X _22154_/X VGND VGND VPWR
+ VPWR _22430_/X sky130_fd_sc_hd__mux4_1
X_34416_ _36144_/CLK _34416_/D VGND VGND VPWR VPWR _34416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31628_ _27751_/X _36025_/Q _31636_/S VGND VGND VPWR VPWR _31629_/A sky130_fd_sc_hd__mux2_1
X_35396_ _35843_/CLK _35396_/D VGND VGND VPWR VPWR _35396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22361_ _33414_/Q _33350_/Q _33286_/Q _33222_/Q _22080_/X _22081_/X VGND VGND VPWR
+ VPWR _22361_/X sky130_fd_sc_hd__mux4_1
X_34347_ _34987_/CLK _34347_/D VGND VGND VPWR VPWR _34347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_248_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31559_ _27649_/X _35992_/Q _31573_/S VGND VGND VPWR VPWR _31560_/A sky130_fd_sc_hd__mux2_1
XFILLER_241_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24100_ _24100_/A VGND VGND VPWR VPWR _32590_/D sky130_fd_sc_hd__clkbuf_1
X_21312_ _22510_/A VGND VGND VPWR VPWR _21312_/X sky130_fd_sc_hd__clkbuf_4
X_25080_ _24920_/X _33021_/Q _25080_/S VGND VGND VPWR VPWR _25081_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22292_ _33924_/Q _33860_/Q _33796_/Q _36100_/Q _21977_/X _21978_/X VGND VGND VPWR
+ VPWR _22292_/X sky130_fd_sc_hd__mux4_1
X_34278_ _34914_/CLK _34278_/D VGND VGND VPWR VPWR _34278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36017_ _36017_/CLK _36017_/D VGND VGND VPWR VPWR _36017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24031_ _24031_/A VGND VGND VPWR VPWR _32557_/D sky130_fd_sc_hd__clkbuf_1
X_33229_ _34186_/CLK _33229_/D VGND VGND VPWR VPWR _33229_/Q sky130_fd_sc_hd__dfxtp_1
X_21243_ _20961_/X _21239_/X _21242_/X _20965_/X VGND VGND VPWR VPWR _21243_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_333_CLK clkbuf_6_44__f_CLK/X VGND VGND VPWR VPWR _36024_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_102_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21174_ _22586_/A VGND VGND VPWR VPWR _21174_/X sky130_fd_sc_hd__buf_4
XFILLER_78_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20125_ _34951_/Q _34887_/Q _34823_/Q _34759_/Q _19813_/X _19814_/X VGND VGND VPWR
+ VPWR _20125_/X sky130_fd_sc_hd__mux4_1
X_28770_ _34702_/Q _27208_/X _28776_/S VGND VGND VPWR VPWR _28771_/A sky130_fd_sc_hd__mux2_1
X_25982_ _24849_/X _33446_/Q _25988_/S VGND VGND VPWR VPWR _25983_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_1443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27721_ _27720_/X _34223_/Q _27733_/S VGND VGND VPWR VPWR _27722_/A sky130_fd_sc_hd__mux2_1
X_20056_ _20056_/A _20056_/B _20056_/C _20056_/D VGND VGND VPWR VPWR _20057_/A sky130_fd_sc_hd__or4_1
X_24933_ input38/X VGND VGND VPWR VPWR _24933_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_133_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27652_ input34/X VGND VGND VPWR VPWR _27652_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24864_ _24864_/A VGND VGND VPWR VPWR _32938_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26603_ _26603_/A VGND VGND VPWR VPWR _33739_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23815_ _23815_/A VGND VGND VPWR VPWR _32392_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27583_ _34171_/Q _27149_/X _27587_/S VGND VGND VPWR VPWR _27584_/A sky130_fd_sc_hd__mux2_1
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24795_ _24795_/A VGND VGND VPWR VPWR _32917_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29322_ _34963_/Q _27223_/X _29326_/S VGND VGND VPWR VPWR _29323_/A sky130_fd_sc_hd__mux2_1
XFILLER_242_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26534_ _26534_/A VGND VGND VPWR VPWR _33706_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20958_ _33118_/Q _35998_/Q _32990_/Q _32926_/Q _20956_/X _20957_/X VGND VGND VPWR
+ VPWR _20958_/X sky130_fd_sc_hd__mux4_1
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23746_ _22943_/X _32360_/Q _23748_/S VGND VGND VPWR VPWR _23747_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29253_ _34930_/Q _27121_/X _29255_/S VGND VGND VPWR VPWR _29254_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26465_ _26465_/A VGND VGND VPWR VPWR _33674_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20889_ _32860_/Q _32796_/Q _32732_/Q _32668_/Q _20887_/X _20888_/X VGND VGND VPWR
+ VPWR _20889_/X sky130_fd_sc_hd__mux4_1
X_23677_ _23677_/A VGND VGND VPWR VPWR _32328_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28204_ _27779_/X _34434_/Q _28214_/S VGND VGND VPWR VPWR _28205_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25416_ _25416_/A VGND VGND VPWR VPWR _33177_/D sky130_fd_sc_hd__clkbuf_1
X_29184_ _29184_/A VGND VGND VPWR VPWR _34897_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_224_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22628_ _22309_/X _22626_/X _22627_/X _22312_/X VGND VGND VPWR VPWR _22628_/X sky130_fd_sc_hd__a22o_1
X_26396_ _26486_/S VGND VGND VPWR VPWR _26415_/S sky130_fd_sc_hd__buf_4
XFILLER_22_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28135_ _27677_/X _34401_/Q _28151_/S VGND VGND VPWR VPWR _28136_/A sky130_fd_sc_hd__mux2_1
X_22559_ _22304_/X _22557_/X _22558_/X _22307_/X VGND VGND VPWR VPWR _22559_/X sky130_fd_sc_hd__a22o_1
XFILLER_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25347_ _33146_/Q _23408_/X _25353_/S VGND VGND VPWR VPWR _25348_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16080_ _17936_/A VGND VGND VPWR VPWR _16080_/X sky130_fd_sc_hd__buf_6
X_28066_ _28066_/A VGND VGND VPWR VPWR _34368_/D sky130_fd_sc_hd__clkbuf_1
X_25278_ _33113_/Q _23240_/X _25290_/S VGND VGND VPWR VPWR _25279_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27017_ _33934_/Q _23475_/X _27023_/S VGND VGND VPWR VPWR _27018_/A sky130_fd_sc_hd__mux2_1
X_24229_ _32650_/Q _23463_/X _24243_/S VGND VGND VPWR VPWR _24230_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_1283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_324_CLK clkbuf_6_39__f_CLK/X VGND VGND VPWR VPWR _32903_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_68_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19770_ _19453_/X _19768_/X _19769_/X _19456_/X VGND VGND VPWR VPWR _19770_/X sky130_fd_sc_hd__a22o_1
XFILLER_231_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16982_ _33648_/Q _33584_/Q _33520_/Q _33456_/Q _16847_/X _16848_/X VGND VGND VPWR
+ VPWR _16982_/X sky130_fd_sc_hd__mux4_1
X_28968_ _28968_/A VGND VGND VPWR VPWR _34794_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18721_ _20099_/A VGND VGND VPWR VPWR _18721_/X sky130_fd_sc_hd__buf_4
XFILLER_49_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27919_ _27757_/X _34299_/Q _27923_/S VGND VGND VPWR VPWR _27920_/A sky130_fd_sc_hd__mux2_1
X_28899_ _34762_/Q _27196_/X _28913_/S VGND VGND VPWR VPWR _28900_/A sky130_fd_sc_hd__mux2_1
XTAP_5151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18652_ _18648_/X _18651_/X _18315_/X VGND VGND VPWR VPWR _18684_/A sky130_fd_sc_hd__o21ba_1
X_30930_ _30930_/A VGND VGND VPWR VPWR _35694_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17603_ _17599_/X _17602_/X _17493_/X _17494_/X VGND VGND VPWR VPWR _17620_/B sky130_fd_sc_hd__o211a_1
XFILLER_18_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30861_ _35662_/Q input52/X _30867_/S VGND VGND VPWR VPWR _30862_/A sky130_fd_sc_hd__mux2_1
X_18583_ _32604_/Q _32540_/Q _32476_/Q _35932_/Q _18517_/X _20017_/A VGND VGND VPWR
+ VPWR _18583_/X sky130_fd_sc_hd__mux4_1
XTAP_4494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32600_ _35735_/CLK _32600_/D VGND VGND VPWR VPWR _32600_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17534_ _17420_/X _17532_/X _17533_/X _17424_/X VGND VGND VPWR VPWR _17534_/X sky130_fd_sc_hd__a22o_1
XTAP_3793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33580_ _34093_/CLK _33580_/D VGND VGND VPWR VPWR _33580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30792_ _35629_/Q input16/X _30804_/S VGND VGND VPWR VPWR _30793_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32531_ _36051_/CLK _32531_/D VGND VGND VPWR VPWR _32531_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17465_ _33085_/Q _32061_/Q _35837_/Q _35773_/Q _17431_/X _17432_/X VGND VGND VPWR
+ VPWR _17465_/X sky130_fd_sc_hd__mux4_1
XFILLER_33_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19204_ _33069_/Q _32045_/Q _35821_/Q _35757_/Q _19025_/X _19026_/X VGND VGND VPWR
+ VPWR _19204_/X sky130_fd_sc_hd__mux4_1
X_16416_ _16416_/A _16416_/B _16416_/C _16416_/D VGND VGND VPWR VPWR _16417_/A sky130_fd_sc_hd__or4_4
X_35250_ _35764_/CLK _35250_/D VGND VGND VPWR VPWR _35250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32462_ _36079_/CLK _32462_/D VGND VGND VPWR VPWR _32462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17396_ _34683_/Q _34619_/Q _34555_/Q _34491_/Q _17292_/X _17293_/X VGND VGND VPWR
+ VPWR _17396_/X sky130_fd_sc_hd__mux4_1
X_34201_ _36121_/CLK _34201_/D VGND VGND VPWR VPWR _34201_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31413_ _31413_/A VGND VGND VPWR VPWR _35923_/D sky130_fd_sc_hd__clkbuf_1
X_19135_ _18950_/X _19133_/X _19134_/X _18953_/X VGND VGND VPWR VPWR _19135_/X sky130_fd_sc_hd__a22o_1
XFILLER_192_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16347_ _34142_/Q _34078_/Q _34014_/Q _33950_/Q _16009_/X _16011_/X VGND VGND VPWR
+ VPWR _16347_/X sky130_fd_sc_hd__mux4_1
X_35181_ _35181_/CLK _35181_/D VGND VGND VPWR VPWR _35181_/Q sky130_fd_sc_hd__dfxtp_1
X_32393_ _35978_/CLK _32393_/D VGND VGND VPWR VPWR _32393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34132_ _34773_/CLK _34132_/D VGND VGND VPWR VPWR _34132_/Q sky130_fd_sc_hd__dfxtp_1
X_19066_ _34921_/Q _34857_/Q _34793_/Q _34729_/Q _18754_/X _18755_/X VGND VGND VPWR
+ VPWR _19066_/X sky130_fd_sc_hd__mux4_1
X_31344_ _31344_/A VGND VGND VPWR VPWR _35890_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16278_ _16140_/X _16276_/X _16277_/X _16145_/X VGND VGND VPWR VPWR _16278_/X sky130_fd_sc_hd__a22o_1
XFILLER_218_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18017_ _33165_/Q _36045_/Q _33037_/Q _32973_/Q _17768_/X _17769_/X VGND VGND VPWR
+ VPWR _18017_/X sky130_fd_sc_hd__mux4_1
X_34063_ _34193_/CLK _34063_/D VGND VGND VPWR VPWR _34063_/Q sky130_fd_sc_hd__dfxtp_1
X_31275_ _27828_/X _35858_/Q _31281_/S VGND VGND VPWR VPWR _31276_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_315_CLK clkbuf_6_48__f_CLK/X VGND VGND VPWR VPWR _35980_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_172_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33014_ _34485_/CLK _33014_/D VGND VGND VPWR VPWR _33014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30226_ _30226_/A VGND VGND VPWR VPWR _35360_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30157_ _35328_/Q _29460_/X _30171_/S VGND VGND VPWR VPWR _30158_/A sky130_fd_sc_hd__mux2_1
X_19968_ _19720_/X _19966_/X _19967_/X _19724_/X VGND VGND VPWR VPWR _19968_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18919_ _18915_/X _18918_/X _18745_/X VGND VGND VPWR VPWR _18927_/C sky130_fd_sc_hd__o21ba_1
XFILLER_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34965_ _36181_/CLK _34965_/D VGND VGND VPWR VPWR _34965_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30088_ _30088_/A VGND VGND VPWR VPWR _35295_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19899_ _19712_/X _19897_/X _19898_/X _19718_/X VGND VGND VPWR VPWR _19899_/X sky130_fd_sc_hd__a22o_1
X_33916_ _36093_/CLK _33916_/D VGND VGND VPWR VPWR _33916_/Q sky130_fd_sc_hd__dfxtp_1
X_21930_ _34937_/Q _34873_/Q _34809_/Q _34745_/Q _21760_/X _21761_/X VGND VGND VPWR
+ VPWR _21930_/X sky130_fd_sc_hd__mux4_1
X_34896_ _34961_/CLK _34896_/D VGND VGND VPWR VPWR _34896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21861_ _35191_/Q _35127_/Q _35063_/Q _32247_/Q _21610_/X _21611_/X VGND VGND VPWR
+ VPWR _21861_/X sky130_fd_sc_hd__mux4_1
XFILLER_94_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33847_ _33910_/CLK _33847_/D VGND VGND VPWR VPWR _33847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20812_ _20740_/X _20810_/X _20811_/X _20745_/X VGND VGND VPWR VPWR _20812_/X sky130_fd_sc_hd__a22o_1
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23600_ _22931_/X _32292_/Q _23610_/S VGND VGND VPWR VPWR _23601_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33778_ _36082_/CLK _33778_/D VGND VGND VPWR VPWR _33778_/Q sky130_fd_sc_hd__dfxtp_1
X_21792_ _21753_/X _21790_/X _21791_/X _21756_/X VGND VGND VPWR VPWR _21792_/X sky130_fd_sc_hd__a22o_1
X_24580_ _22965_/X _32815_/Q _24588_/S VGND VGND VPWR VPWR _24581_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23531_ _23531_/A VGND VGND VPWR VPWR _32260_/D sky130_fd_sc_hd__clkbuf_1
X_20743_ _33624_/Q _33560_/Q _33496_/Q _33432_/Q _20741_/X _20742_/X VGND VGND VPWR
+ VPWR _20743_/X sky130_fd_sc_hd__mux4_1
X_35517_ _35708_/CLK _35517_/D VGND VGND VPWR VPWR _35517_/Q sky130_fd_sc_hd__dfxtp_1
X_32729_ _35865_/CLK _32729_/D VGND VGND VPWR VPWR _32729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23462_ _23462_/A VGND VGND VPWR VPWR _32232_/D sky130_fd_sc_hd__clkbuf_1
X_26250_ _24846_/X _33573_/Q _26258_/S VGND VGND VPWR VPWR _26251_/A sky130_fd_sc_hd__mux2_1
X_20674_ input75/X input76/X VGND VGND VPWR VPWR _22457_/A sky130_fd_sc_hd__or2_4
XFILLER_23_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35448_ _35448_/CLK _35448_/D VGND VGND VPWR VPWR _35448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22413_ _22409_/X _22412_/X _22093_/X _22094_/X VGND VGND VPWR VPWR _22428_/B sky130_fd_sc_hd__o211a_1
X_25201_ _33077_/Q _23393_/X _25217_/S VGND VGND VPWR VPWR _25202_/A sky130_fd_sc_hd__mux2_1
X_26181_ _26181_/A VGND VGND VPWR VPWR _33540_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23393_ input25/X VGND VGND VPWR VPWR _23393_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_12_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35379_ _35764_/CLK _35379_/D VGND VGND VPWR VPWR _35379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22344_ _22304_/X _22342_/X _22343_/X _22307_/X VGND VGND VPWR VPWR _22344_/X sky130_fd_sc_hd__a22o_1
X_25132_ _25132_/A _27232_/A _27232_/B VGND VGND VPWR VPWR _25133_/A sky130_fd_sc_hd__or3b_1
XFILLER_12_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_1308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29940_ _35225_/Q _29339_/X _29952_/S VGND VGND VPWR VPWR _29941_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25063_ _25063_/A VGND VGND VPWR VPWR _33012_/D sky130_fd_sc_hd__clkbuf_1
X_22275_ _35459_/Q _35395_/Q _35331_/Q _35267_/Q _22207_/X _22208_/X VGND VGND VPWR
+ VPWR _22275_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_306_CLK clkbuf_6_50__f_CLK/X VGND VGND VPWR VPWR _33160_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_178_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24014_ _24014_/A VGND VGND VPWR VPWR _32549_/D sky130_fd_sc_hd__clkbuf_1
X_21226_ _21222_/X _21225_/X _21059_/X VGND VGND VPWR VPWR _21227_/D sky130_fd_sc_hd__o21ba_1
X_29871_ _29871_/A VGND VGND VPWR VPWR _35192_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28822_ _28822_/A VGND VGND VPWR VPWR _34725_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21157_ _34403_/Q _36131_/Q _34275_/Q _34211_/Q _21123_/X _21124_/X VGND VGND VPWR
+ VPWR _21157_/X sky130_fd_sc_hd__mux4_1
XFILLER_104_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20108_ _33159_/Q _36039_/Q _33031_/Q _32967_/Q _20068_/X _20069_/X VGND VGND VPWR
+ VPWR _20108_/X sky130_fd_sc_hd__mux4_1
X_28753_ _34694_/Q _27183_/X _28755_/S VGND VGND VPWR VPWR _28754_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25965_ _24824_/X _33438_/Q _25967_/S VGND VGND VPWR VPWR _25966_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21088_ _34913_/Q _34849_/Q _34785_/Q _34721_/Q _21054_/X _21055_/X VGND VGND VPWR
+ VPWR _21088_/X sky130_fd_sc_hd__mux4_2
XFILLER_4_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_875 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27704_ input13/X VGND VGND VPWR VPWR _27704_/X sky130_fd_sc_hd__buf_2
X_20039_ _32901_/Q _32837_/Q _32773_/Q _32709_/Q _19999_/X _20000_/X VGND VGND VPWR
+ VPWR _20039_/X sky130_fd_sc_hd__mux4_1
X_24916_ _24916_/A VGND VGND VPWR VPWR _32955_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28684_ _34661_/Q _27081_/X _28692_/S VGND VGND VPWR VPWR _28685_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25896_ _25896_/A VGND VGND VPWR VPWR _33405_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27635_ _34196_/Q _27226_/X _27637_/S VGND VGND VPWR VPWR _27636_/A sky130_fd_sc_hd__mux2_1
XFILLER_206_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24847_ _24846_/X _32933_/Q _24859_/S VGND VGND VPWR VPWR _24848_/A sky130_fd_sc_hd__mux2_1
XTAP_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27566_ _34163_/Q _27124_/X _27566_/S VGND VGND VPWR VPWR _27567_/A sky130_fd_sc_hd__mux2_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24778_ _23058_/X _32909_/Q _24786_/S VGND VGND VPWR VPWR _24779_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29305_ _29305_/A VGND VGND VPWR VPWR _34954_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26517_ _26517_/A VGND VGND VPWR VPWR _33698_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23729_ _23840_/S VGND VGND VPWR VPWR _23748_/S sky130_fd_sc_hd__buf_4
X_27497_ _27497_/A VGND VGND VPWR VPWR _34130_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29236_ _29326_/S VGND VGND VPWR VPWR _29255_/S sky130_fd_sc_hd__buf_4
X_17250_ _17246_/X _17249_/X _17140_/X _17141_/X VGND VGND VPWR VPWR _17267_/B sky130_fd_sc_hd__o211a_1
X_26448_ _26448_/A VGND VGND VPWR VPWR _33666_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16201_ _34649_/Q _34585_/Q _34521_/Q _34457_/Q _16079_/X _16080_/X VGND VGND VPWR
+ VPWR _16201_/X sky130_fd_sc_hd__mux4_1
XFILLER_174_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29167_ _34889_/Q _27193_/X _29183_/S VGND VGND VPWR VPWR _29168_/A sky130_fd_sc_hd__mux2_1
X_17181_ _17067_/X _17179_/X _17180_/X _17071_/X VGND VGND VPWR VPWR _17181_/X sky130_fd_sc_hd__a22o_1
XFILLER_224_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26379_ _26379_/A VGND VGND VPWR VPWR _33633_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28118_ _27652_/X _34393_/Q _28130_/S VGND VGND VPWR VPWR _28119_/A sky130_fd_sc_hd__mux2_1
X_16132_ _35159_/Q _35095_/Q _35031_/Q _32151_/Q _16083_/X _16085_/X VGND VGND VPWR
+ VPWR _16132_/X sky130_fd_sc_hd__mux4_1
XFILLER_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29098_ _29098_/A VGND VGND VPWR VPWR _34856_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16063_ _16063_/A VGND VGND VPWR VPWR _17851_/A sky130_fd_sc_hd__buf_12
XFILLER_157_1419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28049_ _28049_/A VGND VGND VPWR VPWR _34360_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31060_ _35756_/Q input15/X _31074_/S VGND VGND VPWR VPWR _31061_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_1192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30011_ _35259_/Q _29444_/X _30015_/S VGND VGND VPWR VPWR _30012_/A sky130_fd_sc_hd__mux2_1
X_19822_ _33663_/Q _33599_/Q _33535_/Q _33471_/Q _19500_/X _19501_/X VGND VGND VPWR
+ VPWR _19822_/X sky130_fd_sc_hd__mux4_1
XFILLER_29_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19753_ _19749_/X _19752_/X _19432_/X VGND VGND VPWR VPWR _19775_/A sky130_fd_sc_hd__o21ba_1
X_16965_ _17800_/A VGND VGND VPWR VPWR _16965_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_209_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18704_ _18592_/X _18702_/X _18703_/X _18595_/X VGND VGND VPWR VPWR _18704_/X sky130_fd_sc_hd__a22o_1
X_34750_ _34945_/CLK _34750_/D VGND VGND VPWR VPWR _34750_/Q sky130_fd_sc_hd__dfxtp_1
X_31962_ _34148_/CLK _31962_/D VGND VGND VPWR VPWR _31962_/Q sky130_fd_sc_hd__dfxtp_1
X_19684_ _19359_/X _19682_/X _19683_/X _19365_/X VGND VGND VPWR VPWR _19684_/X sky130_fd_sc_hd__a22o_1
X_16896_ _16714_/X _16894_/X _16895_/X _16718_/X VGND VGND VPWR VPWR _16896_/X sky130_fd_sc_hd__a22o_1
X_18635_ _18597_/X _18633_/X _18634_/X _18600_/X VGND VGND VPWR VPWR _18635_/X sky130_fd_sc_hd__a22o_1
X_30913_ _30913_/A VGND VGND VPWR VPWR _35686_/D sky130_fd_sc_hd__clkbuf_1
X_33701_ _35620_/CLK _33701_/D VGND VGND VPWR VPWR _33701_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34681_ _36152_/CLK _34681_/D VGND VGND VPWR VPWR _34681_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31893_ _31893_/A VGND VGND VPWR VPWR _36150_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33632_ _34594_/CLK _33632_/D VGND VGND VPWR VPWR _33632_/Q sky130_fd_sc_hd__dfxtp_1
X_18566_ _18562_/X _18565_/X _18375_/X VGND VGND VPWR VPWR _18574_/C sky130_fd_sc_hd__o21ba_1
X_30844_ _35654_/Q input43/X _30846_/S VGND VGND VPWR VPWR _30845_/A sky130_fd_sc_hd__mux2_1
XTAP_3590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17517_ _17511_/X _17512_/X _17515_/X _17516_/X VGND VGND VPWR VPWR _17517_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33563_ _36211_/CLK _33563_/D VGND VGND VPWR VPWR _33563_/Q sky130_fd_sc_hd__dfxtp_1
X_18497_ _35417_/Q _35353_/Q _35289_/Q _35225_/Q _18495_/X _18496_/X VGND VGND VPWR
+ VPWR _18497_/X sky130_fd_sc_hd__mux4_1
X_30775_ _35621_/Q input7/X _30783_/S VGND VGND VPWR VPWR _30776_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32514_ _36037_/CLK _32514_/D VGND VGND VPWR VPWR _32514_/Q sky130_fd_sc_hd__dfxtp_1
X_35302_ _35367_/CLK _35302_/D VGND VGND VPWR VPWR _35302_/Q sky130_fd_sc_hd__dfxtp_1
X_17448_ _34173_/Q _34109_/Q _34045_/Q _33981_/Q _17446_/X _17447_/X VGND VGND VPWR
+ VPWR _17448_/X sky130_fd_sc_hd__mux4_1
XFILLER_162_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33494_ _35861_/CLK _33494_/D VGND VGND VPWR VPWR _33494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32445_ _33895_/CLK _32445_/D VGND VGND VPWR VPWR _32445_/Q sky130_fd_sc_hd__dfxtp_1
X_35233_ _35297_/CLK _35233_/D VGND VGND VPWR VPWR _35233_/Q sky130_fd_sc_hd__dfxtp_1
X_17379_ _33915_/Q _33851_/Q _33787_/Q _36091_/Q _17377_/X _17378_/X VGND VGND VPWR
+ VPWR _17379_/X sky130_fd_sc_hd__mux4_1
XFILLER_146_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_92_CLK clkbuf_leaf_96_CLK/A VGND VGND VPWR VPWR _33821_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_118_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19118_ _18793_/X _19116_/X _19117_/X _18798_/X VGND VGND VPWR VPWR _19118_/X sky130_fd_sc_hd__a22o_1
X_35164_ _35610_/CLK _35164_/D VGND VGND VPWR VPWR _35164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20390_ _34703_/Q _34639_/Q _34575_/Q _34511_/Q _20298_/X _20299_/X VGND VGND VPWR
+ VPWR _20390_/X sky130_fd_sc_hd__mux4_1
X_32376_ _32889_/CLK _32376_/D VGND VGND VPWR VPWR _32376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34115_ _34179_/CLK _34115_/D VGND VGND VPWR VPWR _34115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_817 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19049_ _33129_/Q _36009_/Q _33001_/Q _32937_/Q _19009_/X _19010_/X VGND VGND VPWR
+ VPWR _19049_/X sky130_fd_sc_hd__mux4_1
X_31327_ _27704_/X _35882_/Q _31345_/S VGND VGND VPWR VPWR _31328_/A sky130_fd_sc_hd__mux2_1
X_35095_ _35799_/CLK _35095_/D VGND VGND VPWR VPWR _35095_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput200 _36233_/Q VGND VGND VPWR VPWR D2[51] sky130_fd_sc_hd__buf_2
XFILLER_146_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput211 _36243_/Q VGND VGND VPWR VPWR D2[61] sky130_fd_sc_hd__buf_2
XFILLER_173_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput222 _32419_/Q VGND VGND VPWR VPWR D3[13] sky130_fd_sc_hd__buf_2
XFILLER_133_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34046_ _35454_/CLK _34046_/D VGND VGND VPWR VPWR _34046_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput233 _32429_/Q VGND VGND VPWR VPWR D3[23] sky130_fd_sc_hd__buf_2
X_22060_ _22056_/X _22059_/X _21740_/X _21741_/X VGND VGND VPWR VPWR _22075_/B sky130_fd_sc_hd__o211a_1
X_31258_ _31258_/A VGND VGND VPWR VPWR _35849_/D sky130_fd_sc_hd__clkbuf_1
Xoutput244 _32439_/Q VGND VGND VPWR VPWR D3[33] sky130_fd_sc_hd__buf_2
XFILLER_86_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput255 _32449_/Q VGND VGND VPWR VPWR D3[43] sky130_fd_sc_hd__buf_2
X_21011_ _20678_/X _21009_/X _21010_/X _20688_/X VGND VGND VPWR VPWR _21011_/X sky130_fd_sc_hd__a22o_1
Xoutput266 _32459_/Q VGND VGND VPWR VPWR D3[53] sky130_fd_sc_hd__buf_2
X_30209_ _30209_/A VGND VGND VPWR VPWR _35352_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput277 _32469_/Q VGND VGND VPWR VPWR D3[63] sky130_fd_sc_hd__buf_2
XFILLER_58_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_245_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31189_ _27701_/X _35817_/Q _31189_/S VGND VGND VPWR VPWR _31190_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35997_ _35997_/CLK _35997_/D VGND VGND VPWR VPWR _35997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25750_ _24905_/X _33336_/Q _25760_/S VGND VGND VPWR VPWR _25751_/A sky130_fd_sc_hd__mux2_1
X_34948_ _34949_/CLK _34948_/D VGND VGND VPWR VPWR _34948_/Q sky130_fd_sc_hd__dfxtp_1
X_22962_ input17/X VGND VGND VPWR VPWR _22962_/X sky130_fd_sc_hd__buf_2
XFILLER_56_834 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24701_ _24701_/A VGND VGND VPWR VPWR _32872_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21913_ _32121_/Q _32313_/Q _32377_/Q _35897_/Q _21880_/X _21668_/X VGND VGND VPWR
+ VPWR _21913_/X sky130_fd_sc_hd__mux4_1
XFILLER_244_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25681_ _24803_/X _33303_/Q _25697_/S VGND VGND VPWR VPWR _25682_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22893_ _22893_/A VGND VGND VPWR VPWR _32023_/D sky130_fd_sc_hd__clkbuf_1
X_34879_ _36161_/CLK _34879_/D VGND VGND VPWR VPWR _34879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27420_ _27420_/A VGND VGND VPWR VPWR _34093_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24632_ _24659_/S VGND VGND VPWR VPWR _24651_/S sky130_fd_sc_hd__buf_4
XFILLER_130_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21844_ _32631_/Q _32567_/Q _32503_/Q _35959_/Q _21523_/X _21660_/X VGND VGND VPWR
+ VPWR _21844_/X sky130_fd_sc_hd__mux4_1
XFILLER_215_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27351_ _34061_/Q _27205_/X _27359_/S VGND VGND VPWR VPWR _27352_/A sky130_fd_sc_hd__mux2_1
X_24563_ _22940_/X _32807_/Q _24567_/S VGND VGND VPWR VPWR _24564_/A sky130_fd_sc_hd__mux2_1
X_21775_ _21771_/X _21774_/X _21732_/X VGND VGND VPWR VPWR _21797_/A sky130_fd_sc_hd__o21ba_1
XFILLER_12_904 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26302_ _26350_/S VGND VGND VPWR VPWR _26321_/S sky130_fd_sc_hd__buf_6
XFILLER_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20726_ _20648_/X _20724_/X _20725_/X _20658_/X VGND VGND VPWR VPWR _20726_/X sky130_fd_sc_hd__a22o_1
XFILLER_168_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23514_ _23514_/A VGND VGND VPWR VPWR _32252_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27282_ _34028_/Q _27103_/X _27296_/S VGND VGND VPWR VPWR _27283_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24494_ _24494_/A VGND VGND VPWR VPWR _32774_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29021_ _34820_/Q _27177_/X _29027_/S VGND VGND VPWR VPWR _29022_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26233_ _24821_/X _33565_/Q _26237_/S VGND VGND VPWR VPWR _26234_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23445_ _32227_/Q _23444_/X _23451_/S VGND VGND VPWR VPWR _23446_/A sky130_fd_sc_hd__mux2_1
X_20657_ _22371_/A VGND VGND VPWR VPWR _22462_/A sky130_fd_sc_hd__buf_12
XFILLER_109_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_83_CLK clkbuf_leaf_88_CLK/A VGND VGND VPWR VPWR _35998_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_20_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26164_ _26164_/A VGND VGND VPWR VPWR _33532_/D sky130_fd_sc_hd__clkbuf_1
X_23376_ _23376_/A VGND VGND VPWR VPWR _32203_/D sky130_fd_sc_hd__clkbuf_1
X_20588_ _33622_/Q _33558_/Q _33494_/Q _33430_/Q _20584_/X _20587_/X VGND VGND VPWR
+ VPWR _20588_/X sky130_fd_sc_hd__mux4_1
XFILLER_137_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25115_ _25115_/A VGND VGND VPWR VPWR _33037_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22327_ _34181_/Q _34117_/Q _34053_/Q _33989_/Q _22046_/X _22047_/X VGND VGND VPWR
+ VPWR _22327_/X sky130_fd_sc_hd__mux4_1
XFILLER_180_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26095_ _26095_/A VGND VGND VPWR VPWR _33499_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_945 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22258_ _22152_/X _22256_/X _22257_/X _22157_/X VGND VGND VPWR VPWR _22258_/X sky130_fd_sc_hd__a22o_1
X_29923_ _29923_/A VGND VGND VPWR VPWR _35217_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25046_ _25046_/A VGND VGND VPWR VPWR _33004_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_1162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21209_ _20961_/X _21207_/X _21208_/X _20965_/X VGND VGND VPWR VPWR _21209_/X sky130_fd_sc_hd__a22o_1
X_29854_ _29854_/A VGND VGND VPWR VPWR _35184_/D sky130_fd_sc_hd__clkbuf_1
X_22189_ _22189_/A VGND VGND VPWR VPWR _36224_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_239_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28805_ _28805_/A VGND VGND VPWR VPWR _34717_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_238_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29785_ _35152_/Q _29509_/X _29787_/S VGND VGND VPWR VPWR _29786_/A sky130_fd_sc_hd__mux2_1
X_26997_ _26997_/A VGND VGND VPWR VPWR _33924_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28736_ _28784_/S VGND VGND VPWR VPWR _28755_/S sky130_fd_sc_hd__buf_4
XFILLER_150_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16750_ _16706_/X _16748_/X _16749_/X _16712_/X VGND VGND VPWR VPWR _16750_/X sky130_fd_sc_hd__a22o_1
X_25948_ _26080_/S VGND VGND VPWR VPWR _25967_/S sky130_fd_sc_hd__buf_6
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_992 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28667_ _34653_/Q _27056_/X _28671_/S VGND VGND VPWR VPWR _28668_/A sky130_fd_sc_hd__mux2_1
X_16681_ _16361_/X _16679_/X _16680_/X _16365_/X VGND VGND VPWR VPWR _16681_/X sky130_fd_sc_hd__a22o_1
X_25879_ _24896_/X _33397_/Q _25895_/S VGND VGND VPWR VPWR _25880_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18420_ _32087_/Q _32279_/Q _32343_/Q _35863_/Q _18332_/X _20167_/A VGND VGND VPWR
+ VPWR _18420_/X sky130_fd_sc_hd__mux4_1
X_27618_ _27618_/A VGND VGND VPWR VPWR _34187_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28598_ _27763_/X _34621_/Q _28598_/S VGND VGND VPWR VPWR _28599_/A sky130_fd_sc_hd__mux2_1
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18351_ _35670_/Q _32175_/Q _35542_/Q _35478_/Q _18349_/X _18350_/X VGND VGND VPWR
+ VPWR _18351_/X sky130_fd_sc_hd__mux4_1
XFILLER_163_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27549_ _27549_/A VGND VGND VPWR VPWR _34154_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ _17302_/A VGND VGND VPWR VPWR _31992_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18282_ input77/X VGND VGND VPWR VPWR _18361_/A sky130_fd_sc_hd__buf_6
X_30560_ _35519_/Q _29457_/X _30576_/S VGND VGND VPWR VPWR _30561_/A sky130_fd_sc_hd__mux2_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29219_ _29219_/A VGND VGND VPWR VPWR _34913_/D sky130_fd_sc_hd__clkbuf_1
X_17233_ _17158_/X _17231_/X _17232_/X _17163_/X VGND VGND VPWR VPWR _17233_/X sky130_fd_sc_hd__a22o_1
XFILLER_230_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30491_ _30491_/A VGND VGND VPWR VPWR _35486_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_74_CLK clkbuf_leaf_77_CLK/A VGND VGND VPWR VPWR _36052_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32230_ _35722_/CLK _32230_/D VGND VGND VPWR VPWR _32230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17164_ _17158_/X _17159_/X _17162_/X _17163_/X VGND VGND VPWR VPWR _17164_/X sky130_fd_sc_hd__a22o_1
XFILLER_196_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16115_ _16001_/X _16111_/X _16114_/X _16007_/X VGND VGND VPWR VPWR _16115_/X sky130_fd_sc_hd__a22o_1
XFILLER_155_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32161_ _35297_/CLK _32161_/D VGND VGND VPWR VPWR _32161_/Q sky130_fd_sc_hd__dfxtp_1
X_17095_ _34163_/Q _34099_/Q _34035_/Q _33971_/Q _17093_/X _17094_/X VGND VGND VPWR
+ VPWR _17095_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31112_ _35781_/Q input42/X _31116_/S VGND VGND VPWR VPWR _31113_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16046_ _17847_/A VGND VGND VPWR VPWR _16046_/X sky130_fd_sc_hd__buf_4
XFILLER_142_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32092_ _36052_/CLK _32092_/D VGND VGND VPWR VPWR _32092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35920_ _35985_/CLK _35920_/D VGND VGND VPWR VPWR _35920_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_1015 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31043_ _35748_/Q input6/X _31053_/S VGND VGND VPWR VPWR _31044_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19805_ _19800_/X _19803_/X _19804_/X VGND VGND VPWR VPWR _19820_/C sky130_fd_sc_hd__o21ba_1
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35851_ _35852_/CLK _35851_/D VGND VGND VPWR VPWR _35851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17997_ _17993_/X _17996_/X _17857_/X VGND VGND VPWR VPWR _18007_/C sky130_fd_sc_hd__o21ba_1
XFILLER_38_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34802_ _35439_/CLK _34802_/D VGND VGND VPWR VPWR _34802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16948_ _16948_/A _16948_/B _16948_/C _16948_/D VGND VGND VPWR VPWR _16949_/A sky130_fd_sc_hd__or4_4
X_19736_ _34684_/Q _34620_/Q _34556_/Q _34492_/Q _19592_/X _19593_/X VGND VGND VPWR
+ VPWR _19736_/X sky130_fd_sc_hd__mux4_1
X_35782_ _35845_/CLK _35782_/D VGND VGND VPWR VPWR _35782_/Q sky130_fd_sc_hd__dfxtp_1
X_32994_ _36129_/CLK _32994_/D VGND VGND VPWR VPWR _32994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34733_ _35566_/CLK _34733_/D VGND VGND VPWR VPWR _34733_/Q sky130_fd_sc_hd__dfxtp_1
X_31945_ _31945_/A VGND VGND VPWR VPWR _36175_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16879_ _34924_/Q _34860_/Q _34796_/Q _34732_/Q _16807_/X _16808_/X VGND VGND VPWR
+ VPWR _16879_/X sky130_fd_sc_hd__mux4_1
X_19667_ _34426_/Q _36154_/Q _34298_/Q _34234_/Q _19529_/X _19530_/X VGND VGND VPWR
+ VPWR _19667_/X sky130_fd_sc_hd__mux4_1
XFILLER_226_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18618_ _20150_/A VGND VGND VPWR VPWR _18618_/X sky130_fd_sc_hd__buf_6
XFILLER_80_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34664_ _34921_/CLK _34664_/D VGND VGND VPWR VPWR _34664_/Q sky130_fd_sc_hd__dfxtp_1
X_19598_ _34936_/Q _34872_/Q _34808_/Q _34744_/Q _19460_/X _19461_/X VGND VGND VPWR
+ VPWR _19598_/X sky130_fd_sc_hd__mux4_1
X_31876_ _31876_/A VGND VGND VPWR VPWR _36142_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33615_ _34064_/CLK _33615_/D VGND VGND VPWR VPWR _33615_/Q sky130_fd_sc_hd__dfxtp_1
X_30827_ _30875_/S VGND VGND VPWR VPWR _30846_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_52_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18549_ _18447_/X _18547_/X _18548_/X _18450_/X VGND VGND VPWR VPWR _18549_/X sky130_fd_sc_hd__a22o_1
XFILLER_90_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34595_ _36209_/CLK _34595_/D VGND VGND VPWR VPWR _34595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21560_ _32111_/Q _32303_/Q _32367_/Q _35887_/Q _21527_/X _21315_/X VGND VGND VPWR
+ VPWR _21560_/X sky130_fd_sc_hd__mux4_1
X_33546_ _33869_/CLK _33546_/D VGND VGND VPWR VPWR _33546_/Q sky130_fd_sc_hd__dfxtp_1
X_30758_ _35613_/Q input62/X _30762_/S VGND VGND VPWR VPWR _30759_/A sky130_fd_sc_hd__mux2_1
XFILLER_221_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20511_ _35219_/Q _35155_/Q _35091_/Q _32275_/Q _18392_/X _18394_/X VGND VGND VPWR
+ VPWR _20511_/X sky130_fd_sc_hd__mux4_1
XFILLER_127_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33477_ _34179_/CLK _33477_/D VGND VGND VPWR VPWR _33477_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_509_CLK clkbuf_leaf_2_CLK/A VGND VGND VPWR VPWR _34149_/CLK sky130_fd_sc_hd__clkbuf_16
X_21491_ _32621_/Q _32557_/Q _32493_/Q _35949_/Q _21170_/X _21307_/X VGND VGND VPWR
+ VPWR _21491_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_65_CLK clkbuf_leaf_65_CLK/A VGND VGND VPWR VPWR _35986_/CLK sky130_fd_sc_hd__clkbuf_16
X_30689_ _30689_/A VGND VGND VPWR VPWR _35580_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_1018 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23230_ _29797_/A _30472_/A VGND VGND VPWR VPWR _23565_/S sky130_fd_sc_hd__nor2_8
X_35216_ _35217_/CLK _35216_/D VGND VGND VPWR VPWR _35216_/Q sky130_fd_sc_hd__dfxtp_1
X_20442_ _20438_/X _20441_/X _20146_/X _20147_/X VGND VGND VPWR VPWR _20457_/B sky130_fd_sc_hd__o211a_1
XFILLER_119_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32428_ _36068_/CLK _32428_/D VGND VGND VPWR VPWR _32428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36196_ _36202_/CLK _36196_/D VGND VGND VPWR VPWR _36196_/Q sky130_fd_sc_hd__dfxtp_1
X_23161_ _22990_/X _32119_/Q _23173_/S VGND VGND VPWR VPWR _23162_/A sky130_fd_sc_hd__mux2_1
X_20373_ _33935_/Q _33871_/Q _33807_/Q _36111_/Q _18362_/X _18364_/X VGND VGND VPWR
+ VPWR _20373_/X sky130_fd_sc_hd__mux4_1
X_35147_ _35147_/CLK _35147_/D VGND VGND VPWR VPWR _35147_/Q sky130_fd_sc_hd__dfxtp_1
X_32359_ _32552_/CLK _32359_/D VGND VGND VPWR VPWR _32359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22112_ _34430_/Q _36158_/Q _34302_/Q _34238_/Q _21829_/X _21830_/X VGND VGND VPWR
+ VPWR _22112_/X sky130_fd_sc_hd__mux4_1
XTAP_7119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23092_ _22879_/X _32086_/Q _23110_/S VGND VGND VPWR VPWR _23093_/A sky130_fd_sc_hd__mux2_1
X_35078_ _35721_/CLK _35078_/D VGND VGND VPWR VPWR _35078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34029_ _35693_/CLK _34029_/D VGND VGND VPWR VPWR _34029_/Q sky130_fd_sc_hd__dfxtp_1
X_26920_ _27031_/S VGND VGND VPWR VPWR _26939_/S sky130_fd_sc_hd__buf_4
XFILLER_47_1032 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22043_ _22043_/A _22043_/B _22043_/C _22043_/D VGND VGND VPWR VPWR _22044_/A sky130_fd_sc_hd__or4_4
XTAP_6429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1013 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26851_ _33855_/Q _23426_/X _26867_/S VGND VGND VPWR VPWR _26852_/A sky130_fd_sc_hd__mux2_1
XFILLER_134_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25802_ _24982_/X _33361_/Q _25802_/S VGND VGND VPWR VPWR _25803_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29570_ _29660_/S VGND VGND VPWR VPWR _29589_/S sky130_fd_sc_hd__buf_6
X_26782_ _26782_/A VGND VGND VPWR VPWR _33822_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23994_ _22906_/X _32540_/Q _24000_/S VGND VGND VPWR VPWR _23995_/A sky130_fd_sc_hd__mux2_1
XFILLER_228_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28521_ _27649_/X _34584_/Q _28535_/S VGND VGND VPWR VPWR _28522_/A sky130_fd_sc_hd__mux2_1
X_25733_ _24880_/X _33328_/Q _25739_/S VGND VGND VPWR VPWR _25734_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22945_ _22945_/A VGND VGND VPWR VPWR _32040_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_216_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28452_ _28452_/A VGND VGND VPWR VPWR _34551_/D sky130_fd_sc_hd__clkbuf_1
X_25664_ _25664_/A VGND VGND VPWR VPWR _33295_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_189_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22876_ _22872_/X _22875_/X _22471_/A VGND VGND VPWR VPWR _22877_/D sky130_fd_sc_hd__o21ba_1
X_27403_ _27403_/A VGND VGND VPWR VPWR _34085_/D sky130_fd_sc_hd__clkbuf_1
X_24615_ _24615_/A VGND VGND VPWR VPWR _32831_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28383_ _28383_/A VGND VGND VPWR VPWR _34518_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21827_ _35190_/Q _35126_/Q _35062_/Q _32246_/Q _21610_/X _21611_/X VGND VGND VPWR
+ VPWR _21827_/X sky130_fd_sc_hd__mux4_1
X_25595_ _25595_/A VGND VGND VPWR VPWR _33262_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27334_ _34053_/Q _27180_/X _27338_/S VGND VGND VPWR VPWR _27335_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24546_ _22915_/X _32799_/Q _24546_/S VGND VGND VPWR VPWR _24547_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21758_ _21758_/A VGND VGND VPWR VPWR _21758_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_238_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20709_ _34135_/Q _34071_/Q _34007_/Q _33943_/Q _20609_/X _20611_/X VGND VGND VPWR
+ VPWR _20709_/X sky130_fd_sc_hd__mux4_1
X_27265_ _34020_/Q _27078_/X _27275_/S VGND VGND VPWR VPWR _27266_/A sky130_fd_sc_hd__mux2_1
X_24477_ _23011_/X _32766_/Q _24495_/S VGND VGND VPWR VPWR _24478_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_56_CLK clkbuf_leaf_57_CLK/A VGND VGND VPWR VPWR _32808_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_12_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21689_ _21685_/X _21688_/X _21412_/X VGND VGND VPWR VPWR _21690_/D sky130_fd_sc_hd__o21ba_1
X_29004_ _34812_/Q _27152_/X _29006_/S VGND VGND VPWR VPWR _29005_/A sky130_fd_sc_hd__mux2_1
X_26216_ _26216_/A VGND VGND VPWR VPWR _33557_/D sky130_fd_sc_hd__clkbuf_1
X_23428_ _23428_/A VGND VGND VPWR VPWR _32221_/D sky130_fd_sc_hd__clkbuf_1
X_27196_ input48/X VGND VGND VPWR VPWR _27196_/X sky130_fd_sc_hd__buf_4
XFILLER_11_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26147_ _24892_/X _33524_/Q _26165_/S VGND VGND VPWR VPWR _26148_/A sky130_fd_sc_hd__mux2_1
X_23359_ _32196_/Q _23289_/X _23359_/S VGND VGND VPWR VPWR _23360_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26078_ _24991_/X _33492_/Q _26080_/S VGND VGND VPWR VPWR _26079_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29906_ _35209_/Q _29488_/X _29922_/S VGND VGND VPWR VPWR _29907_/A sky130_fd_sc_hd__mux2_1
X_17920_ _17765_/X _17918_/X _17919_/X _17771_/X VGND VGND VPWR VPWR _17920_/X sky130_fd_sc_hd__a22o_1
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25029_ _25029_/A VGND VGND VPWR VPWR _32996_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17851_ _17851_/A VGND VGND VPWR VPWR _17851_/X sky130_fd_sc_hd__clkbuf_4
XTAP_6963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29837_ _29837_/A VGND VGND VPWR VPWR _35176_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_6_45__f_CLK clkbuf_5_22_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_45__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XTAP_6985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16802_ _35178_/Q _35114_/Q _35050_/Q _32170_/Q _16657_/X _16658_/X VGND VGND VPWR
+ VPWR _16802_/X sky130_fd_sc_hd__mux4_1
XTAP_6996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17782_ _17704_/X _17780_/X _17781_/X _17707_/X VGND VGND VPWR VPWR _17782_/X sky130_fd_sc_hd__a22o_1
XFILLER_226_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29768_ _29795_/S VGND VGND VPWR VPWR _29787_/S sky130_fd_sc_hd__buf_4
XFILLER_219_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19521_ _19298_/X _19519_/X _19520_/X _19301_/X VGND VGND VPWR VPWR _19521_/X sky130_fd_sc_hd__a22o_1
X_16733_ _34408_/Q _36136_/Q _34280_/Q _34216_/Q _16523_/X _16524_/X VGND VGND VPWR
+ VPWR _16733_/X sky130_fd_sc_hd__mux4_1
X_28719_ _28719_/A VGND VGND VPWR VPWR _34677_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29699_ _35111_/Q _29382_/X _29703_/S VGND VGND VPWR VPWR _29700_/A sky130_fd_sc_hd__mux2_1
XFILLER_235_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31730_ _31730_/A VGND VGND VPWR VPWR _36073_/D sky130_fd_sc_hd__clkbuf_1
X_19452_ _19447_/X _19450_/X _19451_/X VGND VGND VPWR VPWR _19467_/C sky130_fd_sc_hd__o21ba_1
X_16664_ _16660_/X _16663_/X _16459_/X VGND VGND VPWR VPWR _16665_/D sky130_fd_sc_hd__o21ba_1
XFILLER_234_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18403_ input82/X input81/X VGND VGND VPWR VPWR _20171_/A sky130_fd_sc_hd__or2b_4
XFILLER_201_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31661_ _31661_/A VGND VGND VPWR VPWR _36040_/D sky130_fd_sc_hd__clkbuf_1
X_19383_ _34674_/Q _34610_/Q _34546_/Q _34482_/Q _19239_/X _19240_/X VGND VGND VPWR
+ VPWR _19383_/X sky130_fd_sc_hd__mux4_1
XFILLER_76_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16595_ _16595_/A _16595_/B _16595_/C _16595_/D VGND VGND VPWR VPWR _16596_/A sky130_fd_sc_hd__or4_2
XFILLER_76_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30612_ _30612_/A VGND VGND VPWR VPWR _35543_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18334_ _20074_/A VGND VGND VPWR VPWR _20167_/A sky130_fd_sc_hd__buf_8
X_33400_ _36090_/CLK _33400_/D VGND VGND VPWR VPWR _33400_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34380_ _35661_/CLK _34380_/D VGND VGND VPWR VPWR _34380_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31592_ _27698_/X _36008_/Q _31594_/S VGND VGND VPWR VPWR _31593_/A sky130_fd_sc_hd__mux2_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33331_ _33393_/CLK _33331_/D VGND VGND VPWR VPWR _33331_/Q sky130_fd_sc_hd__dfxtp_1
X_18265_ _15981_/X _18263_/X _18264_/X _15991_/X VGND VGND VPWR VPWR _18265_/X sky130_fd_sc_hd__a22o_1
XFILLER_163_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30543_ _35511_/Q _29432_/X _30555_/S VGND VGND VPWR VPWR _30544_/A sky130_fd_sc_hd__mux2_1
XFILLER_198_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_47_CLK clkbuf_leaf_49_CLK/A VGND VGND VPWR VPWR _35755_/CLK sky130_fd_sc_hd__clkbuf_16
X_17216_ _32886_/Q _32822_/Q _32758_/Q _32694_/Q _16993_/X _16994_/X VGND VGND VPWR
+ VPWR _17216_/X sky130_fd_sc_hd__mux4_1
XFILLER_175_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36050_ _36051_/CLK _36050_/D VGND VGND VPWR VPWR _36050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33262_ _36079_/CLK _33262_/D VGND VGND VPWR VPWR _33262_/Q sky130_fd_sc_hd__dfxtp_1
X_30474_ _35478_/Q _29328_/X _30492_/S VGND VGND VPWR VPWR _30475_/A sky130_fd_sc_hd__mux2_1
X_18196_ _32659_/Q _32595_/Q _32531_/Q _35987_/Q _17982_/X _16877_/A VGND VGND VPWR
+ VPWR _18196_/X sky130_fd_sc_hd__mux4_1
X_32213_ _35704_/CLK _32213_/D VGND VGND VPWR VPWR _32213_/Q sky130_fd_sc_hd__dfxtp_1
X_35001_ _35769_/CLK _35001_/D VGND VGND VPWR VPWR _35001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17147_ _16998_/X _17143_/X _17146_/X _17001_/X VGND VGND VPWR VPWR _17147_/X sky130_fd_sc_hd__a22o_1
X_33193_ _36073_/CLK _33193_/D VGND VGND VPWR VPWR _33193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32144_ _35921_/CLK _32144_/D VGND VGND VPWR VPWR _32144_/Q sky130_fd_sc_hd__dfxtp_1
X_17078_ _17935_/A VGND VGND VPWR VPWR _17078_/X sky130_fd_sc_hd__buf_6
XFILLER_226_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16029_ _17773_/A VGND VGND VPWR VPWR _17912_/A sky130_fd_sc_hd__buf_12
X_32075_ _36042_/CLK _32075_/D VGND VGND VPWR VPWR _32075_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31026_ _35740_/Q input61/X _31032_/S VGND VGND VPWR VPWR _31027_/A sky130_fd_sc_hd__mux2_1
X_35903_ _35903_/CLK _35903_/D VGND VGND VPWR VPWR _35903_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_1238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35834_ _36026_/CLK _35834_/D VGND VGND VPWR VPWR _35834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19719_ _19712_/X _19714_/X _19717_/X _19718_/X VGND VGND VPWR VPWR _19719_/X sky130_fd_sc_hd__a22o_1
X_20991_ _33375_/Q _33311_/Q _33247_/Q _33183_/Q _20602_/X _20603_/X VGND VGND VPWR
+ VPWR _20991_/X sky130_fd_sc_hd__mux4_1
X_35765_ _35765_/CLK _35765_/D VGND VGND VPWR VPWR _35765_/Q sky130_fd_sc_hd__dfxtp_1
X_32977_ _35855_/CLK _32977_/D VGND VGND VPWR VPWR _32977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22730_ _34193_/Q _34129_/Q _34065_/Q _34001_/Q _20649_/X _20650_/X VGND VGND VPWR
+ VPWR _22730_/X sky130_fd_sc_hd__mux4_1
X_34716_ _36242_/CLK _34716_/D VGND VGND VPWR VPWR _34716_/Q sky130_fd_sc_hd__dfxtp_1
X_31928_ _31928_/A VGND VGND VPWR VPWR _36167_/D sky130_fd_sc_hd__clkbuf_1
X_35696_ _35697_/CLK _35696_/D VGND VGND VPWR VPWR _35696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34647_ _34647_/CLK _34647_/D VGND VGND VPWR VPWR _34647_/Q sky130_fd_sc_hd__dfxtp_1
X_22661_ _35214_/Q _35150_/Q _35086_/Q _32270_/Q _20692_/X _20694_/X VGND VGND VPWR
+ VPWR _22661_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31859_ _31859_/A VGND VGND VPWR VPWR _36134_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24400_ _24400_/A VGND VGND VPWR VPWR _32729_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21612_ _35184_/Q _35120_/Q _35056_/Q _32187_/Q _21610_/X _21611_/X VGND VGND VPWR
+ VPWR _21612_/X sky130_fd_sc_hd__mux4_1
X_25380_ _25380_/A VGND VGND VPWR VPWR _33161_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_240_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34578_ _34708_/CLK _34578_/D VGND VGND VPWR VPWR _34578_/Q sky130_fd_sc_hd__dfxtp_1
X_22592_ _35660_/Q _35020_/Q _34380_/Q _33740_/Q _22450_/X _22451_/X VGND VGND VPWR
+ VPWR _22592_/X sky130_fd_sc_hd__mux4_1
XFILLER_187_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24331_ _22996_/X _32697_/Q _24339_/S VGND VGND VPWR VPWR _24332_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33529_ _35641_/CLK _33529_/D VGND VGND VPWR VPWR _33529_/Q sky130_fd_sc_hd__dfxtp_1
X_21543_ _21400_/X _21541_/X _21542_/X _21403_/X VGND VGND VPWR VPWR _21543_/X sky130_fd_sc_hd__a22o_1
XFILLER_107_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_38_CLK clkbuf_6_7__f_CLK/X VGND VGND VPWR VPWR _35875_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_193_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27050_ input56/X VGND VGND VPWR VPWR _27050_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_138_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24262_ _22894_/X _32664_/Q _24276_/S VGND VGND VPWR VPWR _24263_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21474_ _35180_/Q _35116_/Q _35052_/Q _32172_/Q _21257_/X _21258_/X VGND VGND VPWR
+ VPWR _21474_/X sky130_fd_sc_hd__mux4_1
XFILLER_222_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26001_ _24877_/X _33455_/Q _26009_/S VGND VGND VPWR VPWR _26002_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_1064 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20425_ _20164_/X _20423_/X _20424_/X _20169_/X VGND VGND VPWR VPWR _20425_/X sky130_fd_sc_hd__a22o_1
XFILLER_140_1072 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23213_ _23067_/X _32144_/Q _23215_/S VGND VGND VPWR VPWR _23214_/A sky130_fd_sc_hd__mux2_1
XFILLER_134_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36179_ _36179_/CLK _36179_/D VGND VGND VPWR VPWR _36179_/Q sky130_fd_sc_hd__dfxtp_1
X_24193_ _32633_/Q _23405_/X _24201_/S VGND VGND VPWR VPWR _24194_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20356_ _35470_/Q _35406_/Q _35342_/Q _35278_/Q _20260_/X _20261_/X VGND VGND VPWR
+ VPWR _20356_/X sky130_fd_sc_hd__mux4_1
X_23144_ _22965_/X _32111_/Q _23152_/S VGND VGND VPWR VPWR _23145_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27952_ _27952_/A VGND VGND VPWR VPWR _34314_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23075_ _23075_/A VGND VGND VPWR VPWR _32082_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20287_ _32140_/Q _32332_/Q _32396_/Q _35916_/Q _20286_/X _20074_/X VGND VGND VPWR
+ VPWR _20287_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_1132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26903_ _26903_/A VGND VGND VPWR VPWR _33879_/D sky130_fd_sc_hd__clkbuf_1
X_22026_ _22019_/X _22025_/X _21740_/X _21741_/X VGND VGND VPWR VPWR _22043_/B sky130_fd_sc_hd__o211a_1
XFILLER_96_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27883_ _27973_/S VGND VGND VPWR VPWR _27902_/S sky130_fd_sc_hd__buf_4
XTAP_5536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29622_ _29622_/A VGND VGND VPWR VPWR _35074_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26834_ _33847_/Q _23399_/X _26846_/S VGND VGND VPWR VPWR _26835_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_248_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29553_ _29553_/A VGND VGND VPWR VPWR _35041_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26765_ _33814_/Q _23225_/X _26783_/S VGND VGND VPWR VPWR _26766_/A sky130_fd_sc_hd__mux2_1
XTAP_4879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23977_ _23082_/X _32533_/Q _23977_/S VGND VGND VPWR VPWR _23978_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_1152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28504_ _28504_/A VGND VGND VPWR VPWR _34576_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_216_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25716_ _24855_/X _33320_/Q _25718_/S VGND VGND VPWR VPWR _25717_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29484_ input46/X VGND VGND VPWR VPWR _29484_/X sky130_fd_sc_hd__clkbuf_4
X_22928_ input5/X VGND VGND VPWR VPWR _22928_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_205_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26696_ _26696_/A VGND VGND VPWR VPWR _33781_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_954 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28435_ _28435_/A VGND VGND VPWR VPWR _34543_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25647_ _25647_/A VGND VGND VPWR VPWR _33287_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22859_ _32149_/Q _32341_/Q _32405_/Q _35925_/Q _22586_/X _21611_/A VGND VGND VPWR
+ VPWR _22859_/X sky130_fd_sc_hd__mux4_1
XFILLER_227_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16380_ _34398_/Q _36126_/Q _34270_/Q _34206_/Q _16170_/X _16171_/X VGND VGND VPWR
+ VPWR _16380_/X sky130_fd_sc_hd__mux4_1
X_28366_ _27819_/X _34511_/Q _28370_/S VGND VGND VPWR VPWR _28367_/A sky130_fd_sc_hd__mux2_1
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25578_ _25578_/A VGND VGND VPWR VPWR _33254_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27317_ _34045_/Q _27155_/X _27317_/S VGND VGND VPWR VPWR _27318_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24529_ _24529_/A VGND VGND VPWR VPWR _32790_/D sky130_fd_sc_hd__clkbuf_1
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28297_ _27717_/X _34478_/Q _28307_/S VGND VGND VPWR VPWR _28298_/A sky130_fd_sc_hd__mux2_1
XPHY_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_29_CLK clkbuf_6_5__f_CLK/X VGND VGND VPWR VPWR _36202_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_240_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18050_ _32910_/Q _32846_/Q _32782_/Q _32718_/Q _15984_/X _15987_/X VGND VGND VPWR
+ VPWR _18050_/X sky130_fd_sc_hd__mux4_1
X_27248_ _34012_/Q _27053_/X _27254_/S VGND VGND VPWR VPWR _27249_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17001_ _17862_/A VGND VGND VPWR VPWR _17001_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_177_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27179_ _27179_/A VGND VGND VPWR VPWR _33988_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30190_ _35344_/Q _29509_/X _30192_/S VGND VGND VPWR VPWR _30191_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18952_ _33062_/Q _32038_/Q _35814_/Q _35750_/Q _18672_/X _18673_/X VGND VGND VPWR
+ VPWR _18952_/X sky130_fd_sc_hd__mux4_1
XFILLER_140_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17903_ _17903_/A _17903_/B _17903_/C _17903_/D VGND VGND VPWR VPWR _17904_/A sky130_fd_sc_hd__or4_2
XFILLER_105_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18883_ _33060_/Q _32036_/Q _35812_/Q _35748_/Q _18672_/X _18673_/X VGND VGND VPWR
+ VPWR _18883_/X sky130_fd_sc_hd__mux4_1
XTAP_6760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32900_ _35973_/CLK _32900_/D VGND VGND VPWR VPWR _32900_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17834_ _17834_/A VGND VGND VPWR VPWR _17834_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_66_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33880_ _36057_/CLK _33880_/D VGND VGND VPWR VPWR _33880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32831_ _32895_/CLK _32831_/D VGND VGND VPWR VPWR _32831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17765_ _17765_/A VGND VGND VPWR VPWR _17765_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_19_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19504_ _20210_/A VGND VGND VPWR VPWR _19504_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_169_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35550_ _35551_/CLK _35550_/D VGND VGND VPWR VPWR _35550_/Q sky130_fd_sc_hd__dfxtp_1
X_16716_ _32104_/Q _32296_/Q _32360_/Q _35880_/Q _16574_/X _16715_/X VGND VGND VPWR
+ VPWR _16716_/X sky130_fd_sc_hd__mux4_1
X_17696_ _33156_/Q _36036_/Q _33028_/Q _32964_/Q _17415_/X _17416_/X VGND VGND VPWR
+ VPWR _17696_/X sky130_fd_sc_hd__mux4_1
X_32762_ _32891_/CLK _32762_/D VGND VGND VPWR VPWR _32762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34501_ _34694_/CLK _34501_/D VGND VGND VPWR VPWR _34501_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31713_ _36065_/Q input3/X _31729_/S VGND VGND VPWR VPWR _31714_/A sky130_fd_sc_hd__mux2_1
X_16647_ _35622_/Q _34982_/Q _34342_/Q _33702_/Q _16438_/X _16439_/X VGND VGND VPWR
+ VPWR _16647_/X sky130_fd_sc_hd__mux4_1
X_19435_ _33140_/Q _36020_/Q _33012_/Q _32948_/Q _19362_/X _19363_/X VGND VGND VPWR
+ VPWR _19435_/X sky130_fd_sc_hd__mux4_1
X_35481_ _35482_/CLK _35481_/D VGND VGND VPWR VPWR _35481_/Q sky130_fd_sc_hd__dfxtp_1
X_32693_ _32904_/CLK _32693_/D VGND VGND VPWR VPWR _32693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34432_ _34815_/CLK _34432_/D VGND VGND VPWR VPWR _34432_/Q sky130_fd_sc_hd__dfxtp_1
X_31644_ _31644_/A VGND VGND VPWR VPWR _36032_/D sky130_fd_sc_hd__clkbuf_1
X_19366_ _19359_/X _19361_/X _19364_/X _19365_/X VGND VGND VPWR VPWR _19366_/X sky130_fd_sc_hd__a22o_1
X_16578_ _16573_/X _16577_/X _16434_/X _16435_/X VGND VGND VPWR VPWR _16595_/B sky130_fd_sc_hd__o211a_1
XFILLER_241_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18317_ _20065_/A VGND VGND VPWR VPWR _20205_/A sky130_fd_sc_hd__buf_12
X_34363_ _36154_/CLK _34363_/D VGND VGND VPWR VPWR _34363_/Q sky130_fd_sc_hd__dfxtp_1
X_31575_ _31686_/S VGND VGND VPWR VPWR _31594_/S sky130_fd_sc_hd__buf_4
X_19297_ _19291_/X _19296_/X _19087_/X _19088_/X VGND VGND VPWR VPWR _19318_/B sky130_fd_sc_hd__o211a_1
XFILLER_198_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36102_ _36102_/CLK _36102_/D VGND VGND VPWR VPWR _36102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18248_ _18248_/A VGND VGND VPWR VPWR _32020_/D sky130_fd_sc_hd__clkbuf_2
X_33314_ _33827_/CLK _33314_/D VGND VGND VPWR VPWR _33314_/Q sky130_fd_sc_hd__dfxtp_1
X_30526_ _35503_/Q _29407_/X _30534_/S VGND VGND VPWR VPWR _30527_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34294_ _35126_/CLK _34294_/D VGND VGND VPWR VPWR _34294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36033_ _36033_/CLK _36033_/D VGND VGND VPWR VPWR _36033_/Q sky130_fd_sc_hd__dfxtp_1
X_18179_ _18175_/X _18178_/X _17857_/A VGND VGND VPWR VPWR _18187_/C sky130_fd_sc_hd__o21ba_1
X_30457_ _30457_/A VGND VGND VPWR VPWR _35470_/D sky130_fd_sc_hd__clkbuf_1
X_33245_ _36205_/CLK _33245_/D VGND VGND VPWR VPWR _33245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20210_ _20210_/A VGND VGND VPWR VPWR _20210_/X sky130_fd_sc_hd__buf_4
X_33176_ _36057_/CLK _33176_/D VGND VGND VPWR VPWR _33176_/Q sky130_fd_sc_hd__dfxtp_1
X_21190_ _21047_/X _21188_/X _21189_/X _21050_/X VGND VGND VPWR VPWR _21190_/X sky130_fd_sc_hd__a22o_1
X_30388_ _30388_/A VGND VGND VPWR VPWR _35437_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20141_ _33160_/Q _36040_/Q _33032_/Q _32968_/Q _20068_/X _20069_/X VGND VGND VPWR
+ VPWR _20141_/X sky130_fd_sc_hd__mux4_1
X_32127_ _32575_/CLK _32127_/D VGND VGND VPWR VPWR _32127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20072_ _20065_/X _20067_/X _20070_/X _20071_/X VGND VGND VPWR VPWR _20072_/X sky130_fd_sc_hd__a22o_1
X_32058_ _35835_/CLK _32058_/D VGND VGND VPWR VPWR _32058_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31009_ _31009_/A VGND VGND VPWR VPWR _35732_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23900_ _22968_/X _32496_/Q _23906_/S VGND VGND VPWR VPWR _23901_/A sky130_fd_sc_hd__mux2_1
XFILLER_246_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24880_ input19/X VGND VGND VPWR VPWR _24880_/X sky130_fd_sc_hd__clkbuf_4
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23831_ _23831_/A VGND VGND VPWR VPWR _32400_/D sky130_fd_sc_hd__clkbuf_1
X_35817_ _35817_/CLK _35817_/D VGND VGND VPWR VPWR _35817_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26550_ _26550_/A VGND VGND VPWR VPWR _33714_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35748_ _35812_/CLK _35748_/D VGND VGND VPWR VPWR _35748_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23762_ _23762_/A VGND VGND VPWR VPWR _32367_/D sky130_fd_sc_hd__clkbuf_1
X_20974_ _33054_/Q _32030_/Q _35806_/Q _35742_/Q _20972_/X _20973_/X VGND VGND VPWR
+ VPWR _20974_/X sky130_fd_sc_hd__mux4_1
XFILLER_26_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25501_ _24936_/X _33218_/Q _25511_/S VGND VGND VPWR VPWR _25502_/A sky130_fd_sc_hd__mux2_1
X_22713_ _35728_/Q _32239_/Q _35600_/Q _35536_/Q _20593_/X _20595_/X VGND VGND VPWR
+ VPWR _22713_/X sky130_fd_sc_hd__mux4_1
XFILLER_246_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26481_ _26481_/A VGND VGND VPWR VPWR _33682_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_213_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23693_ _23693_/A VGND VGND VPWR VPWR _32336_/D sky130_fd_sc_hd__clkbuf_1
X_35679_ _35743_/CLK _35679_/D VGND VGND VPWR VPWR _35679_/Q sky130_fd_sc_hd__dfxtp_1
X_28220_ _28220_/A VGND VGND VPWR VPWR _34441_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_214_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25432_ _24834_/X _33185_/Q _25448_/S VGND VGND VPWR VPWR _25433_/A sky130_fd_sc_hd__mux2_1
X_22644_ _22512_/X _22642_/X _22643_/X _22515_/X VGND VGND VPWR VPWR _22644_/X sky130_fd_sc_hd__a22o_1
XFILLER_213_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28151_ _27701_/X _34409_/Q _28151_/S VGND VGND VPWR VPWR _28152_/A sky130_fd_sc_hd__mux2_1
X_25363_ _25363_/A VGND VGND VPWR VPWR _33153_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22575_ _33676_/Q _33612_/Q _33548_/Q _33484_/Q _22506_/X _22507_/X VGND VGND VPWR
+ VPWR _22575_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_6_9__f_CLK clkbuf_5_4_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_9__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_194_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_895 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27102_ _27102_/A VGND VGND VPWR VPWR _33963_/D sky130_fd_sc_hd__clkbuf_1
X_24314_ _22971_/X _32689_/Q _24318_/S VGND VGND VPWR VPWR _24315_/A sky130_fd_sc_hd__mux2_1
X_28082_ _34376_/Q _27189_/X _28100_/S VGND VGND VPWR VPWR _28083_/A sky130_fd_sc_hd__mux2_1
X_21526_ _21306_/X _21524_/X _21525_/X _21312_/X VGND VGND VPWR VPWR _21526_/X sky130_fd_sc_hd__a22o_1
XFILLER_194_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25294_ _25294_/A VGND VGND VPWR VPWR _33120_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27033_ input1/X VGND VGND VPWR VPWR _27033_/X sky130_fd_sc_hd__buf_4
XFILLER_108_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24245_ _32658_/Q _23487_/X _24251_/S VGND VGND VPWR VPWR _24246_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21457_ _21453_/X _21454_/X _21455_/X _21456_/X VGND VGND VPWR VPWR _21457_/X sky130_fd_sc_hd__a22o_1
X_20408_ _19453_/A _20406_/X _20407_/X _19456_/A VGND VGND VPWR VPWR _20408_/X sky130_fd_sc_hd__a22o_1
XFILLER_147_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24176_ _32625_/Q _23364_/X _24180_/S VGND VGND VPWR VPWR _24177_/A sky130_fd_sc_hd__mux2_1
X_21388_ _22447_/A VGND VGND VPWR VPWR _21388_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_150_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23127_ _22940_/X _32103_/Q _23131_/S VGND VGND VPWR VPWR _23128_/A sky130_fd_sc_hd__mux2_1
X_20339_ _33678_/Q _33614_/Q _33550_/Q _33486_/Q _20206_/X _20207_/X VGND VGND VPWR
+ VPWR _20339_/X sky130_fd_sc_hd__mux4_1
XTAP_6001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28984_ _28984_/A VGND VGND VPWR VPWR _34802_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27935_ _27935_/A VGND VGND VPWR VPWR _34306_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23058_ input51/X VGND VGND VPWR VPWR _23058_/X sky130_fd_sc_hd__buf_2
XTAP_6056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput99 _31976_/Q VGND VGND VPWR VPWR D1[18] sky130_fd_sc_hd__buf_2
XTAP_6067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22009_ _33916_/Q _33852_/Q _33788_/Q _36092_/Q _21977_/X _21978_/X VGND VGND VPWR
+ VPWR _22009_/X sky130_fd_sc_hd__mux4_1
XFILLER_248_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27866_ _27866_/A VGND VGND VPWR VPWR _34273_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29605_ _29605_/A VGND VGND VPWR VPWR _35066_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26817_ _33839_/Q _23316_/X _26825_/S VGND VGND VPWR VPWR _26818_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27797_ input46/X VGND VGND VPWR VPWR _27797_/X sky130_fd_sc_hd__clkbuf_4
XTAP_5399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17550_ _17550_/A _17550_/B _17550_/C _17550_/D VGND VGND VPWR VPWR _17551_/A sky130_fd_sc_hd__or4_1
XTAP_3942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29536_ _29536_/A VGND VGND VPWR VPWR _35033_/D sky130_fd_sc_hd__clkbuf_1
X_26748_ _26748_/A VGND VGND VPWR VPWR _33806_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16501_ _33378_/Q _33314_/Q _33250_/Q _33186_/Q _16421_/X _16422_/X VGND VGND VPWR
+ VPWR _16501_/X sky130_fd_sc_hd__mux4_1
XTAP_3986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17481_ _17834_/A VGND VGND VPWR VPWR _17481_/X sky130_fd_sc_hd__buf_4
X_29467_ _35010_/Q _29466_/X _29482_/S VGND VGND VPWR VPWR _29468_/A sky130_fd_sc_hd__mux2_1
XTAP_3997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26679_ _26679_/A VGND VGND VPWR VPWR _33773_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_225_1209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16432_ _32864_/Q _32800_/Q _32736_/Q _32672_/Q _16287_/X _16288_/X VGND VGND VPWR
+ VPWR _16432_/X sky130_fd_sc_hd__mux4_1
X_19220_ _33902_/Q _33838_/Q _33774_/Q _36078_/Q _18971_/X _18972_/X VGND VGND VPWR
+ VPWR _19220_/X sky130_fd_sc_hd__mux4_1
X_28418_ _28418_/A VGND VGND VPWR VPWR _34535_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29398_ input15/X VGND VGND VPWR VPWR _29398_/X sky130_fd_sc_hd__buf_2
XFILLER_73_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19151_ _20210_/A VGND VGND VPWR VPWR _19151_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_38_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28349_ _27794_/X _34503_/Q _28349_/S VGND VGND VPWR VPWR _28350_/A sky130_fd_sc_hd__mux2_1
X_16363_ _32094_/Q _32286_/Q _32350_/Q _35870_/Q _16221_/X _16362_/X VGND VGND VPWR
+ VPWR _16363_/X sky130_fd_sc_hd__mux4_1
XFILLER_34_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18102_ _33424_/Q _33360_/Q _33296_/Q _33232_/Q _17833_/X _17834_/X VGND VGND VPWR
+ VPWR _18102_/X sky130_fd_sc_hd__mux4_1
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19082_ _33130_/Q _36010_/Q _33002_/Q _32938_/Q _19009_/X _19010_/X VGND VGND VPWR
+ VPWR _19082_/X sky130_fd_sc_hd__mux4_1
X_31360_ _27754_/X _35898_/Q _31366_/S VGND VGND VPWR VPWR _31361_/A sky130_fd_sc_hd__mux2_1
X_16294_ _35612_/Q _34972_/Q _34332_/Q _33692_/Q _16053_/X _16055_/X VGND VGND VPWR
+ VPWR _16294_/X sky130_fd_sc_hd__mux4_1
XFILLER_199_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18033_ _34445_/Q _36173_/Q _34317_/Q _34253_/Q _17935_/X _17936_/X VGND VGND VPWR
+ VPWR _18033_/X sky130_fd_sc_hd__mux4_1
X_30311_ _35401_/Q _29488_/X _30327_/S VGND VGND VPWR VPWR _30312_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31291_ _27652_/X _35865_/Q _31303_/S VGND VGND VPWR VPWR _31292_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_1264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33030_ _36038_/CLK _33030_/D VGND VGND VPWR VPWR _33030_/Q sky130_fd_sc_hd__dfxtp_1
X_30242_ _30242_/A VGND VGND VPWR VPWR _35368_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30173_ _30200_/S VGND VGND VPWR VPWR _30192_/S sky130_fd_sc_hd__buf_4
X_19984_ _19811_/X _19982_/X _19983_/X _19816_/X VGND VGND VPWR VPWR _19984_/X sky130_fd_sc_hd__a22o_1
XFILLER_193_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18935_ _18931_/X _18934_/X _18726_/X VGND VGND VPWR VPWR _18965_/A sky130_fd_sc_hd__o21ba_1
XFILLER_80_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34981_ _35625_/CLK _34981_/D VGND VGND VPWR VPWR _34981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33932_ _36109_/CLK _33932_/D VGND VGND VPWR VPWR _33932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18866_ _33380_/Q _33316_/Q _33252_/Q _33188_/Q _18721_/X _18722_/X VGND VGND VPWR
+ VPWR _18866_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_9_CLK clkbuf_leaf_9_CLK/A VGND VGND VPWR VPWR _34921_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_6590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17817_ _35463_/Q _35399_/Q _35335_/Q _35271_/Q _17607_/X _17608_/X VGND VGND VPWR
+ VPWR _17817_/X sky130_fd_sc_hd__mux4_1
XFILLER_95_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33863_ _36159_/CLK _33863_/D VGND VGND VPWR VPWR _33863_/Q sky130_fd_sc_hd__dfxtp_1
X_18797_ _34146_/Q _34082_/Q _34018_/Q _33954_/Q _18687_/X _18688_/X VGND VGND VPWR
+ VPWR _18797_/X sky130_fd_sc_hd__mux4_1
XFILLER_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35602_ _35730_/CLK _35602_/D VGND VGND VPWR VPWR _35602_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32814_ _32911_/CLK _32814_/D VGND VGND VPWR VPWR _32814_/Q sky130_fd_sc_hd__dfxtp_1
X_17748_ _17744_/X _17747_/X _17504_/X VGND VGND VPWR VPWR _17756_/C sky130_fd_sc_hd__o21ba_1
X_33794_ _36099_/CLK _33794_/D VGND VGND VPWR VPWR _33794_/Q sky130_fd_sc_hd__dfxtp_1
X_35533_ _35663_/CLK _35533_/D VGND VGND VPWR VPWR _35533_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_913 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32745_ _32808_/CLK _32745_/D VGND VGND VPWR VPWR _32745_/Q sky130_fd_sc_hd__dfxtp_1
X_17679_ _34691_/Q _34627_/Q _34563_/Q _34499_/Q _17645_/X _17646_/X VGND VGND VPWR
+ VPWR _17679_/X sky130_fd_sc_hd__mux4_1
XFILLER_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19418_ _34419_/Q _36147_/Q _34291_/Q _34227_/Q _19176_/X _19177_/X VGND VGND VPWR
+ VPWR _19418_/X sky130_fd_sc_hd__mux4_1
X_35464_ _35466_/CLK _35464_/D VGND VGND VPWR VPWR _35464_/Q sky130_fd_sc_hd__dfxtp_1
X_20690_ _22373_/A VGND VGND VPWR VPWR _21758_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_211_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32676_ _32804_/CLK _32676_/D VGND VGND VPWR VPWR _32676_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34415_ _36144_/CLK _34415_/D VGND VGND VPWR VPWR _34415_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19349_ _19345_/X _19348_/X _19112_/X VGND VGND VPWR VPWR _19350_/D sky130_fd_sc_hd__o21ba_1
X_31627_ _31627_/A VGND VGND VPWR VPWR _36024_/D sky130_fd_sc_hd__clkbuf_1
X_35395_ _35651_/CLK _35395_/D VGND VGND VPWR VPWR _35395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22360_ _22152_/X _22358_/X _22359_/X _22157_/X VGND VGND VPWR VPWR _22360_/X sky130_fd_sc_hd__a22o_1
XFILLER_206_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34346_ _34987_/CLK _34346_/D VGND VGND VPWR VPWR _34346_/Q sky130_fd_sc_hd__dfxtp_1
X_31558_ _31558_/A VGND VGND VPWR VPWR _35991_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21311_ _33128_/Q _36008_/Q _33000_/Q _32936_/Q _21309_/X _21310_/X VGND VGND VPWR
+ VPWR _21311_/X sky130_fd_sc_hd__mux4_1
X_22291_ _33412_/Q _33348_/Q _33284_/Q _33220_/Q _22080_/X _22081_/X VGND VGND VPWR
+ VPWR _22291_/X sky130_fd_sc_hd__mux4_1
XFILLER_191_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30509_ _35495_/Q _29382_/X _30513_/S VGND VGND VPWR VPWR _30510_/A sky130_fd_sc_hd__mux2_1
X_34277_ _34405_/CLK _34277_/D VGND VGND VPWR VPWR _34277_/Q sky130_fd_sc_hd__dfxtp_1
X_31489_ _27745_/X _35959_/Q _31501_/S VGND VGND VPWR VPWR _31490_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_1034 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36016_ _36016_/CLK _36016_/D VGND VGND VPWR VPWR _36016_/Q sky130_fd_sc_hd__dfxtp_1
X_24030_ _22959_/X _32557_/Q _24042_/S VGND VGND VPWR VPWR _24031_/A sky130_fd_sc_hd__mux2_1
X_21242_ _32870_/Q _32806_/Q _32742_/Q _32678_/Q _21240_/X _21241_/X VGND VGND VPWR
+ VPWR _21242_/X sky130_fd_sc_hd__mux4_1
X_33228_ _34186_/CLK _33228_/D VGND VGND VPWR VPWR _33228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21173_ _20953_/X _21171_/X _21172_/X _20959_/X VGND VGND VPWR VPWR _21173_/X sky130_fd_sc_hd__a22o_1
X_33159_ _36038_/CLK _33159_/D VGND VGND VPWR VPWR _33159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20124_ _34439_/Q _36167_/Q _34311_/Q _34247_/Q _19882_/X _19883_/X VGND VGND VPWR
+ VPWR _20124_/X sky130_fd_sc_hd__mux4_1
XFILLER_172_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25981_ _25981_/A VGND VGND VPWR VPWR _33445_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27720_ input18/X VGND VGND VPWR VPWR _27720_/X sky130_fd_sc_hd__buf_2
X_20055_ _20051_/X _20054_/X _19818_/X VGND VGND VPWR VPWR _20056_/D sky130_fd_sc_hd__o21ba_1
X_24932_ _24932_/A VGND VGND VPWR VPWR _32960_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_246_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27651_ _27651_/A VGND VGND VPWR VPWR _34200_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24863_ _24861_/X _32938_/Q _24890_/S VGND VGND VPWR VPWR _24864_/A sky130_fd_sc_hd__mux2_1
XTAP_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26602_ _24964_/X _33739_/Q _26614_/S VGND VGND VPWR VPWR _26603_/A sky130_fd_sc_hd__mux2_1
XTAP_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23814_ _23042_/X _32392_/Q _23832_/S VGND VGND VPWR VPWR _23815_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27582_ _27582_/A VGND VGND VPWR VPWR _34170_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24794_ _23082_/X _32917_/Q _24794_/S VGND VGND VPWR VPWR _24795_/A sky130_fd_sc_hd__mux2_1
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29321_ _29321_/A VGND VGND VPWR VPWR _34962_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26533_ _24861_/X _33706_/Q _26551_/S VGND VGND VPWR VPWR _26534_/A sky130_fd_sc_hd__mux2_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23745_ _23745_/A VGND VGND VPWR VPWR _32359_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_242_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20957_ _22507_/A VGND VGND VPWR VPWR _20957_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_784 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29252_ _29252_/A VGND VGND VPWR VPWR _34929_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26464_ _33674_/Q _23463_/X _26478_/S VGND VGND VPWR VPWR _26465_/A sky130_fd_sc_hd__mux2_1
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23676_ _23042_/X _32328_/Q _23694_/S VGND VGND VPWR VPWR _23677_/A sky130_fd_sc_hd__mux2_1
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20888_ _22434_/A VGND VGND VPWR VPWR _20888_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_202_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28203_ _28203_/A VGND VGND VPWR VPWR _34433_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25415_ _24809_/X _33177_/Q _25427_/S VGND VGND VPWR VPWR _25416_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29183_ _34897_/Q _27217_/X _29183_/S VGND VGND VPWR VPWR _29184_/A sky130_fd_sc_hd__mux2_1
X_22627_ _33101_/Q _32077_/Q _35853_/Q _35789_/Q _22384_/X _22385_/X VGND VGND VPWR
+ VPWR _22627_/X sky130_fd_sc_hd__mux4_1
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26395_ _26395_/A VGND VGND VPWR VPWR _33641_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28134_ _28134_/A VGND VGND VPWR VPWR _34400_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25346_ _25346_/A VGND VGND VPWR VPWR _33145_/D sky130_fd_sc_hd__clkbuf_1
X_22558_ _35659_/Q _35019_/Q _34379_/Q _33739_/Q _22450_/X _22451_/X VGND VGND VPWR
+ VPWR _22558_/X sky130_fd_sc_hd__mux4_1
XFILLER_166_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28065_ _34368_/Q _27165_/X _28079_/S VGND VGND VPWR VPWR _28066_/A sky130_fd_sc_hd__mux2_1
X_21509_ _21400_/X _21507_/X _21508_/X _21403_/X VGND VGND VPWR VPWR _21509_/X sky130_fd_sc_hd__a22o_1
X_25277_ _25277_/A VGND VGND VPWR VPWR _33112_/D sky130_fd_sc_hd__clkbuf_1
X_22489_ _35721_/Q _32232_/Q _35593_/Q _35529_/Q _22270_/X _22271_/X VGND VGND VPWR
+ VPWR _22489_/X sky130_fd_sc_hd__mux4_1
X_27016_ _27016_/A VGND VGND VPWR VPWR _33933_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24228_ _24228_/A VGND VGND VPWR VPWR _32649_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24159_ _32617_/Q _23289_/X _24159_/S VGND VGND VPWR VPWR _24160_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28967_ _34794_/Q _27096_/X _28985_/S VGND VGND VPWR VPWR _28968_/A sky130_fd_sc_hd__mux2_1
X_16981_ _16981_/A VGND VGND VPWR VPWR _31983_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18720_ _18440_/X _18718_/X _18719_/X _18445_/X VGND VGND VPWR VPWR _18720_/X sky130_fd_sc_hd__a22o_1
XTAP_5130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27918_ _27918_/A VGND VGND VPWR VPWR _34298_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28898_ _28898_/A VGND VGND VPWR VPWR _34761_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18651_ _18447_/X _18649_/X _18650_/X _18450_/X VGND VGND VPWR VPWR _18651_/X sky130_fd_sc_hd__a22o_1
X_27849_ _27849_/A VGND VGND VPWR VPWR _34265_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17602_ _17420_/X _17600_/X _17601_/X _17424_/X VGND VGND VPWR VPWR _17602_/X sky130_fd_sc_hd__a22o_1
X_30860_ _30860_/A VGND VGND VPWR VPWR _35661_/D sky130_fd_sc_hd__clkbuf_1
X_18582_ _18578_/X _18581_/X _18315_/X VGND VGND VPWR VPWR _18612_/A sky130_fd_sc_hd__o21ba_1
XTAP_4484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29519_ _35027_/Q _29518_/X _29525_/S VGND VGND VPWR VPWR _29520_/A sky130_fd_sc_hd__mux2_1
XTAP_3783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17533_ _32895_/Q _32831_/Q _32767_/Q _32703_/Q _17346_/X _17347_/X VGND VGND VPWR
+ VPWR _17533_/X sky130_fd_sc_hd__mux4_1
XTAP_3794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30791_ _30791_/A VGND VGND VPWR VPWR _35628_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_260_CLK clkbuf_6_62__f_CLK/X VGND VGND VPWR VPWR _34177_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_44_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32530_ _35986_/CLK _32530_/D VGND VGND VPWR VPWR _32530_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17464_ _35453_/Q _35389_/Q _35325_/Q _35261_/Q _17254_/X _17255_/X VGND VGND VPWR
+ VPWR _17464_/X sky130_fd_sc_hd__mux4_1
XFILLER_232_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16415_ _16411_/X _16414_/X _16104_/X VGND VGND VPWR VPWR _16416_/D sky130_fd_sc_hd__o21ba_2
XFILLER_149_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19203_ _35437_/Q _35373_/Q _35309_/Q _35245_/Q _19201_/X _19202_/X VGND VGND VPWR
+ VPWR _19203_/X sky130_fd_sc_hd__mux4_1
XFILLER_242_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32461_ _33904_/CLK _32461_/D VGND VGND VPWR VPWR _32461_/Q sky130_fd_sc_hd__dfxtp_1
X_17395_ _17391_/X _17394_/X _17151_/X VGND VGND VPWR VPWR _17403_/C sky130_fd_sc_hd__o21ba_1
X_34200_ _34907_/CLK _34200_/D VGND VGND VPWR VPWR _34200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31412_ _27831_/X _35923_/Q _31416_/S VGND VGND VPWR VPWR _31413_/A sky130_fd_sc_hd__mux2_1
X_16346_ _33630_/Q _33566_/Q _33502_/Q _33438_/Q _16141_/X _16142_/X VGND VGND VPWR
+ VPWR _16346_/X sky130_fd_sc_hd__mux4_1
X_19134_ _33067_/Q _32043_/Q _35819_/Q _35755_/Q _19025_/X _19026_/X VGND VGND VPWR
+ VPWR _19134_/X sky130_fd_sc_hd__mux4_1
XFILLER_201_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32392_ _35978_/CLK _32392_/D VGND VGND VPWR VPWR _32392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35180_ _35180_/CLK _35180_/D VGND VGND VPWR VPWR _35180_/Q sky130_fd_sc_hd__dfxtp_1
X_34131_ _34897_/CLK _34131_/D VGND VGND VPWR VPWR _34131_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19065_ _34409_/Q _36137_/Q _34281_/Q _34217_/Q _18823_/X _18824_/X VGND VGND VPWR
+ VPWR _19065_/X sky130_fd_sc_hd__mux4_1
X_31343_ _27729_/X _35890_/Q _31345_/S VGND VGND VPWR VPWR _31344_/A sky130_fd_sc_hd__mux2_1
X_16277_ _34140_/Q _34076_/Q _34012_/Q _33948_/Q _16009_/X _16011_/X VGND VGND VPWR
+ VPWR _16277_/X sky130_fd_sc_hd__mux4_1
XFILLER_146_848 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18016_ _32653_/Q _32589_/Q _32525_/Q _35981_/Q _17982_/X _17766_/X VGND VGND VPWR
+ VPWR _18016_/X sky130_fd_sc_hd__mux4_1
X_34062_ _34192_/CLK _34062_/D VGND VGND VPWR VPWR _34062_/Q sky130_fd_sc_hd__dfxtp_1
X_31274_ _31274_/A VGND VGND VPWR VPWR _35857_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_13_0_CLK clkbuf_5_9_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_13_0_CLK/X sky130_fd_sc_hd__clkbuf_8
X_33013_ _36020_/CLK _33013_/D VGND VGND VPWR VPWR _33013_/Q sky130_fd_sc_hd__dfxtp_1
X_30225_ _35360_/Q _29360_/X _30243_/S VGND VGND VPWR VPWR _30226_/A sky130_fd_sc_hd__mux2_1
XFILLER_236_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30156_ _30156_/A VGND VGND VPWR VPWR _35327_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19967_ _32899_/Q _32835_/Q _32771_/Q _32707_/Q _19646_/X _19647_/X VGND VGND VPWR
+ VPWR _19967_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18918_ _18597_/X _18916_/X _18917_/X _18600_/X VGND VGND VPWR VPWR _18918_/X sky130_fd_sc_hd__a22o_1
X_34964_ _34964_/CLK _34964_/D VGND VGND VPWR VPWR _34964_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_5_28_0_CLK clkbuf_2_3_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_28_0_CLK/X sky130_fd_sc_hd__clkbuf_8
X_30087_ _35295_/Q _29357_/X _30087_/S VGND VGND VPWR VPWR _30088_/A sky130_fd_sc_hd__mux2_1
X_19898_ _33153_/Q _36033_/Q _33025_/Q _32961_/Q _19715_/X _19716_/X VGND VGND VPWR
+ VPWR _19898_/X sky130_fd_sc_hd__mux4_1
XFILLER_45_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33915_ _36092_/CLK _33915_/D VGND VGND VPWR VPWR _33915_/Q sky130_fd_sc_hd__dfxtp_1
X_18849_ _20261_/A VGND VGND VPWR VPWR _18849_/X sky130_fd_sc_hd__clkbuf_4
X_34895_ _34961_/CLK _34895_/D VGND VGND VPWR VPWR _34895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33846_ _33910_/CLK _33846_/D VGND VGND VPWR VPWR _33846_/Q sky130_fd_sc_hd__dfxtp_1
X_21860_ _34679_/Q _34615_/Q _34551_/Q _34487_/Q _21539_/X _21540_/X VGND VGND VPWR
+ VPWR _21860_/X sky130_fd_sc_hd__mux4_1
XFILLER_83_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_247_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20811_ _34138_/Q _34074_/Q _34010_/Q _33946_/Q _20609_/X _20611_/X VGND VGND VPWR
+ VPWR _20811_/X sky130_fd_sc_hd__mux4_1
XFILLER_42_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33777_ _36082_/CLK _33777_/D VGND VGND VPWR VPWR _33777_/Q sky130_fd_sc_hd__dfxtp_1
X_21791_ _35189_/Q _35125_/Q _35061_/Q _32242_/Q _21610_/X _21611_/X VGND VGND VPWR
+ VPWR _21791_/X sky130_fd_sc_hd__mux4_1
X_30989_ _30989_/A VGND VGND VPWR VPWR _35722_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_251_CLK clkbuf_6_63__f_CLK/X VGND VGND VPWR VPWR _34183_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_36_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23530_ _32260_/Q _23441_/X _23536_/S VGND VGND VPWR VPWR _23531_/A sky130_fd_sc_hd__mux2_1
X_35516_ _35708_/CLK _35516_/D VGND VGND VPWR VPWR _35516_/Q sky130_fd_sc_hd__dfxtp_1
X_32728_ _35990_/CLK _32728_/D VGND VGND VPWR VPWR _32728_/Q sky130_fd_sc_hd__dfxtp_1
X_20742_ _22507_/A VGND VGND VPWR VPWR _20742_/X sky130_fd_sc_hd__buf_4
XFILLER_168_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23461_ _32232_/Q _23460_/X _23485_/S VGND VGND VPWR VPWR _23462_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35447_ _36153_/CLK _35447_/D VGND VGND VPWR VPWR _35447_/Q sky130_fd_sc_hd__dfxtp_1
X_20673_ _20660_/X _20665_/X _20670_/X _20672_/X VGND VGND VPWR VPWR _20673_/X sky130_fd_sc_hd__a22o_1
X_32659_ _36051_/CLK _32659_/D VGND VGND VPWR VPWR _32659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25200_ _25200_/A VGND VGND VPWR VPWR _33076_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22412_ _22373_/X _22410_/X _22411_/X _22377_/X VGND VGND VPWR VPWR _22412_/X sky130_fd_sc_hd__a22o_1
X_26180_ _24942_/X _33540_/Q _26186_/S VGND VGND VPWR VPWR _26181_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35378_ _35828_/CLK _35378_/D VGND VGND VPWR VPWR _35378_/Q sky130_fd_sc_hd__dfxtp_1
X_23392_ _23392_/A VGND VGND VPWR VPWR _32209_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25131_ _25131_/A VGND VGND VPWR VPWR _33045_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34329_ _35610_/CLK _34329_/D VGND VGND VPWR VPWR _34329_/Q sky130_fd_sc_hd__dfxtp_1
X_22343_ _35653_/Q _35013_/Q _34373_/Q _33733_/Q _22097_/X _22098_/X VGND VGND VPWR
+ VPWR _22343_/X sky130_fd_sc_hd__mux4_1
XFILLER_136_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25062_ _24892_/X _33012_/Q _25080_/S VGND VGND VPWR VPWR _25063_/A sky130_fd_sc_hd__mux2_1
X_22274_ _21951_/X _22272_/X _22273_/X _21954_/X VGND VGND VPWR VPWR _22274_/X sky130_fd_sc_hd__a22o_1
XFILLER_117_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24013_ _22934_/X _32549_/Q _24021_/S VGND VGND VPWR VPWR _24014_/A sky130_fd_sc_hd__mux2_1
X_21225_ _21052_/X _21223_/X _21224_/X _21057_/X VGND VGND VPWR VPWR _21225_/X sky130_fd_sc_hd__a22o_1
X_29870_ _35192_/Q _29435_/X _29880_/S VGND VGND VPWR VPWR _29871_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28821_ _34725_/Q _27081_/X _28829_/S VGND VGND VPWR VPWR _28822_/A sky130_fd_sc_hd__mux2_1
XFILLER_219_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21156_ _21047_/X _21154_/X _21155_/X _21050_/X VGND VGND VPWR VPWR _21156_/X sky130_fd_sc_hd__a22o_1
XFILLER_63_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20107_ _32647_/Q _32583_/Q _32519_/Q _35975_/Q _19929_/X _20066_/X VGND VGND VPWR
+ VPWR _20107_/X sky130_fd_sc_hd__mux4_1
X_28752_ _28752_/A VGND VGND VPWR VPWR _34693_/D sky130_fd_sc_hd__clkbuf_1
X_25964_ _25964_/A VGND VGND VPWR VPWR _33437_/D sky130_fd_sc_hd__clkbuf_1
X_21087_ _34401_/Q _36129_/Q _34273_/Q _34209_/Q _20770_/X _20771_/X VGND VGND VPWR
+ VPWR _21087_/X sky130_fd_sc_hd__mux4_1
XFILLER_8_1444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20038_ _32133_/Q _32325_/Q _32389_/Q _35909_/Q _19933_/X _19721_/X VGND VGND VPWR
+ VPWR _20038_/X sky130_fd_sc_hd__mux4_1
X_27703_ _27703_/A VGND VGND VPWR VPWR _34217_/D sky130_fd_sc_hd__clkbuf_1
X_24915_ _24914_/X _32955_/Q _24921_/S VGND VGND VPWR VPWR _24916_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25895_ _24920_/X _33405_/Q _25895_/S VGND VGND VPWR VPWR _25896_/A sky130_fd_sc_hd__mux2_1
X_28683_ _28683_/A VGND VGND VPWR VPWR _34660_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27634_ _27634_/A VGND VGND VPWR VPWR _34195_/D sky130_fd_sc_hd__clkbuf_1
X_24846_ input7/X VGND VGND VPWR VPWR _24846_/X sky130_fd_sc_hd__buf_4
XFILLER_73_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27565_ _27565_/A VGND VGND VPWR VPWR _34162_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24777_ _24777_/A VGND VGND VPWR VPWR _32908_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21989_ _35707_/Q _32216_/Q _35579_/Q _35515_/Q _21917_/X _21918_/X VGND VGND VPWR
+ VPWR _21989_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_242_CLK clkbuf_6_61__f_CLK/X VGND VGND VPWR VPWR _36104_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_14_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29304_ _34954_/Q _27196_/X _29318_/S VGND VGND VPWR VPWR _29305_/A sky130_fd_sc_hd__mux2_1
X_26516_ _24837_/X _33698_/Q _26530_/S VGND VGND VPWR VPWR _26517_/A sky130_fd_sc_hd__mux2_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23728_ _23728_/A VGND VGND VPWR VPWR _32351_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27496_ _34130_/Q _27220_/X _27502_/S VGND VGND VPWR VPWR _27497_/A sky130_fd_sc_hd__mux2_1
XFILLER_202_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26447_ _33666_/Q _23435_/X _26457_/S VGND VGND VPWR VPWR _26448_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29235_ _29235_/A VGND VGND VPWR VPWR _34921_/D sky130_fd_sc_hd__clkbuf_1
X_23659_ _23018_/X _32320_/Q _23673_/S VGND VGND VPWR VPWR _23660_/A sky130_fd_sc_hd__mux2_1
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16200_ _16194_/X _16199_/X _16075_/X VGND VGND VPWR VPWR _16208_/C sky130_fd_sc_hd__o21ba_1
XFILLER_70_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29166_ _29166_/A VGND VGND VPWR VPWR _34888_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_230_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17180_ _32885_/Q _32821_/Q _32757_/Q _32693_/Q _16993_/X _16994_/X VGND VGND VPWR
+ VPWR _17180_/X sky130_fd_sc_hd__mux4_1
XFILLER_122_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26378_ _33633_/Q _23265_/X _26394_/S VGND VGND VPWR VPWR _26379_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16131_ _34647_/Q _34583_/Q _34519_/Q _34455_/Q _16079_/X _16080_/X VGND VGND VPWR
+ VPWR _16131_/X sky130_fd_sc_hd__mux4_1
X_28117_ _28117_/A VGND VGND VPWR VPWR _34392_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25329_ _25329_/A VGND VGND VPWR VPWR _33137_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29097_ _34856_/Q _27090_/X _29099_/S VGND VGND VPWR VPWR _29098_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16062_ _17850_/A VGND VGND VPWR VPWR _16062_/X sky130_fd_sc_hd__buf_6
XFILLER_143_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28048_ _34360_/Q _27140_/X _28058_/S VGND VGND VPWR VPWR _28049_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30010_ _30010_/A VGND VGND VPWR VPWR _35258_/D sky130_fd_sc_hd__clkbuf_1
X_19821_ _19821_/A VGND VGND VPWR VPWR _32446_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_190_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29999_ _35253_/Q _29426_/X _30015_/S VGND VGND VPWR VPWR _30000_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19752_ _19506_/X _19750_/X _19751_/X _19509_/X VGND VGND VPWR VPWR _19752_/X sky130_fd_sc_hd__a22o_1
X_16964_ _17799_/A VGND VGND VPWR VPWR _16964_/X sky130_fd_sc_hd__buf_4
XFILLER_110_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18703_ _35615_/Q _34975_/Q _34335_/Q _33695_/Q _18353_/X _18355_/X VGND VGND VPWR
+ VPWR _18703_/X sky130_fd_sc_hd__mux4_1
XFILLER_231_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31961_ _34148_/CLK _31961_/D VGND VGND VPWR VPWR _31961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19683_ _33147_/Q _36027_/Q _33019_/Q _32955_/Q _19362_/X _19363_/X VGND VGND VPWR
+ VPWR _19683_/X sky130_fd_sc_hd__mux4_1
XFILLER_238_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16895_ _32877_/Q _32813_/Q _32749_/Q _32685_/Q _16640_/X _16641_/X VGND VGND VPWR
+ VPWR _16895_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_481_CLK _35560_/CLK VGND VGND VPWR VPWR _34091_/CLK sky130_fd_sc_hd__clkbuf_16
X_33700_ _35177_/CLK _33700_/D VGND VGND VPWR VPWR _33700_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18634_ _33053_/Q _32029_/Q _35805_/Q _35741_/Q _18367_/X _18369_/X VGND VGND VPWR
+ VPWR _18634_/X sky130_fd_sc_hd__mux4_1
X_30912_ _35686_/Q input8/X _30918_/S VGND VGND VPWR VPWR _30913_/A sky130_fd_sc_hd__mux2_1
XFILLER_237_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34680_ _35833_/CLK _34680_/D VGND VGND VPWR VPWR _34680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31892_ _23396_/X _36150_/Q _31906_/S VGND VGND VPWR VPWR _31893_/A sky130_fd_sc_hd__mux2_1
XTAP_4292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33631_ _33821_/CLK _33631_/D VGND VGND VPWR VPWR _33631_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18565_ _18360_/X _18563_/X _18564_/X _18372_/X VGND VGND VPWR VPWR _18565_/X sky130_fd_sc_hd__a22o_1
X_30843_ _30843_/A VGND VGND VPWR VPWR _35653_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_233_CLK clkbuf_6_55__f_CLK/X VGND VGND VPWR VPWR _33934_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17516_ _17869_/A VGND VGND VPWR VPWR _17516_/X sky130_fd_sc_hd__clkbuf_4
X_33562_ _36212_/CLK _33562_/D VGND VGND VPWR VPWR _33562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18496_ _20151_/A VGND VGND VPWR VPWR _18496_/X sky130_fd_sc_hd__buf_4
X_30774_ _30774_/A VGND VGND VPWR VPWR _35620_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35301_ _35365_/CLK _35301_/D VGND VGND VPWR VPWR _35301_/Q sky130_fd_sc_hd__dfxtp_1
X_32513_ _35969_/CLK _32513_/D VGND VGND VPWR VPWR _32513_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17447_ _17961_/A VGND VGND VPWR VPWR _17447_/X sky130_fd_sc_hd__buf_8
X_33493_ _33685_/CLK _33493_/D VGND VGND VPWR VPWR _33493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35232_ _36005_/CLK _35232_/D VGND VGND VPWR VPWR _35232_/Q sky130_fd_sc_hd__dfxtp_1
X_32444_ _36075_/CLK _32444_/D VGND VGND VPWR VPWR _32444_/Q sky130_fd_sc_hd__dfxtp_1
X_17378_ _17851_/A VGND VGND VPWR VPWR _17378_/X sky130_fd_sc_hd__buf_6
XFILLER_192_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19117_ _34155_/Q _34091_/Q _34027_/Q _33963_/Q _19040_/X _19041_/X VGND VGND VPWR
+ VPWR _19117_/X sky130_fd_sc_hd__mux4_1
X_35163_ _35800_/CLK _35163_/D VGND VGND VPWR VPWR _35163_/Q sky130_fd_sc_hd__dfxtp_1
X_16329_ _16325_/X _16328_/X _16044_/X _16046_/X VGND VGND VPWR VPWR _16344_/B sky130_fd_sc_hd__o211a_1
XFILLER_174_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32375_ _35895_/CLK _32375_/D VGND VGND VPWR VPWR _32375_/Q sky130_fd_sc_hd__dfxtp_1
X_34114_ _34945_/CLK _34114_/D VGND VGND VPWR VPWR _34114_/Q sky130_fd_sc_hd__dfxtp_1
X_19048_ _32617_/Q _32553_/Q _32489_/Q _35945_/Q _18870_/X _19007_/X VGND VGND VPWR
+ VPWR _19048_/X sky130_fd_sc_hd__mux4_1
X_31326_ _31416_/S VGND VGND VPWR VPWR _31345_/S sky130_fd_sc_hd__buf_4
X_35094_ _36118_/CLK _35094_/D VGND VGND VPWR VPWR _35094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput201 _36234_/Q VGND VGND VPWR VPWR D2[52] sky130_fd_sc_hd__buf_2
XFILLER_133_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput212 _36244_/Q VGND VGND VPWR VPWR D2[62] sky130_fd_sc_hd__buf_2
X_31257_ _27801_/X _35849_/Q _31273_/S VGND VGND VPWR VPWR _31258_/A sky130_fd_sc_hd__mux2_1
Xoutput223 _32420_/Q VGND VGND VPWR VPWR D3[14] sky130_fd_sc_hd__buf_2
X_34045_ _34877_/CLK _34045_/D VGND VGND VPWR VPWR _34045_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput234 _32430_/Q VGND VGND VPWR VPWR D3[24] sky130_fd_sc_hd__buf_2
XFILLER_47_1214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput245 _32440_/Q VGND VGND VPWR VPWR D3[34] sky130_fd_sc_hd__buf_2
XFILLER_160_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput256 _32450_/Q VGND VGND VPWR VPWR D3[44] sky130_fd_sc_hd__buf_2
X_21010_ _35167_/Q _35103_/Q _35039_/Q _32159_/Q _20904_/X _20905_/X VGND VGND VPWR
+ VPWR _21010_/X sky130_fd_sc_hd__mux4_1
Xoutput267 _32460_/Q VGND VGND VPWR VPWR D3[54] sky130_fd_sc_hd__buf_2
XFILLER_86_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30208_ _35352_/Q _29336_/X _30222_/S VGND VGND VPWR VPWR _30209_/A sky130_fd_sc_hd__mux2_1
Xoutput278 _32412_/Q VGND VGND VPWR VPWR D3[6] sky130_fd_sc_hd__buf_2
X_31188_ _31188_/A VGND VGND VPWR VPWR _35816_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30139_ _30139_/A VGND VGND VPWR VPWR _35319_/D sky130_fd_sc_hd__clkbuf_1
X_35996_ _36055_/CLK _35996_/D VGND VGND VPWR VPWR _35996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34947_ _36163_/CLK _34947_/D VGND VGND VPWR VPWR _34947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22961_ _22961_/A VGND VGND VPWR VPWR _32045_/D sky130_fd_sc_hd__clkbuf_1
X_24700_ _22943_/X _32872_/Q _24702_/S VGND VGND VPWR VPWR _24701_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_472_CLK clkbuf_6_10__f_CLK/X VGND VGND VPWR VPWR _35693_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_56_846 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21912_ _21659_/X _21910_/X _21911_/X _21665_/X VGND VGND VPWR VPWR _21912_/X sky130_fd_sc_hd__a22o_1
X_25680_ _25680_/A VGND VGND VPWR VPWR _33302_/D sky130_fd_sc_hd__clkbuf_1
X_34878_ _34942_/CLK _34878_/D VGND VGND VPWR VPWR _34878_/Q sky130_fd_sc_hd__dfxtp_1
X_22892_ _22891_/X _32023_/Q _22916_/S VGND VGND VPWR VPWR _22893_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24631_ _24631_/A VGND VGND VPWR VPWR _32839_/D sky130_fd_sc_hd__clkbuf_1
X_33829_ _35622_/CLK _33829_/D VGND VGND VPWR VPWR _33829_/Q sky130_fd_sc_hd__dfxtp_1
X_21843_ _21839_/X _21842_/X _21732_/X VGND VGND VPWR VPWR _21867_/A sky130_fd_sc_hd__o21ba_1
XFILLER_82_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_224_CLK clkbuf_6_53__f_CLK/X VGND VGND VPWR VPWR _34193_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27350_ _27350_/A VGND VGND VPWR VPWR _34060_/D sky130_fd_sc_hd__clkbuf_1
X_24562_ _24562_/A VGND VGND VPWR VPWR _32806_/D sky130_fd_sc_hd__clkbuf_1
X_21774_ _21453_/X _21772_/X _21773_/X _21456_/X VGND VGND VPWR VPWR _21774_/X sky130_fd_sc_hd__a22o_1
XFILLER_70_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26301_ _26301_/A VGND VGND VPWR VPWR _33597_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23513_ _32252_/Q _23414_/X _23515_/S VGND VGND VPWR VPWR _23514_/A sky130_fd_sc_hd__mux2_1
X_20725_ _35607_/Q _34967_/Q _34327_/Q _33687_/Q _20653_/X _20655_/X VGND VGND VPWR
+ VPWR _20725_/X sky130_fd_sc_hd__mux4_1
X_27281_ _27281_/A VGND VGND VPWR VPWR _34027_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24493_ _23036_/X _32774_/Q _24495_/S VGND VGND VPWR VPWR _24494_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29020_ _29020_/A VGND VGND VPWR VPWR _34819_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26232_ _26232_/A VGND VGND VPWR VPWR _33564_/D sky130_fd_sc_hd__clkbuf_1
X_23444_ input42/X VGND VGND VPWR VPWR _23444_/X sky130_fd_sc_hd__clkbuf_8
X_20656_ _35606_/Q _34966_/Q _34326_/Q _33686_/Q _20653_/X _20655_/X VGND VGND VPWR
+ VPWR _20656_/X sky130_fd_sc_hd__mux4_1
XFILLER_196_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26163_ _24917_/X _33532_/Q _26165_/S VGND VGND VPWR VPWR _26164_/A sky130_fd_sc_hd__mux2_1
X_23375_ _32203_/Q _23316_/X _23385_/S VGND VGND VPWR VPWR _23376_/A sky130_fd_sc_hd__mux2_1
X_20587_ _22507_/A VGND VGND VPWR VPWR _20587_/X sky130_fd_sc_hd__buf_4
XFILLER_221_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25114_ _24970_/X _33037_/Q _25122_/S VGND VGND VPWR VPWR _25115_/A sky130_fd_sc_hd__mux2_1
X_22326_ _33669_/Q _33605_/Q _33541_/Q _33477_/Q _22153_/X _22154_/X VGND VGND VPWR
+ VPWR _22326_/X sky130_fd_sc_hd__mux4_1
X_26094_ _24815_/X _33499_/Q _26102_/S VGND VGND VPWR VPWR _26095_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1008 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29922_ _35217_/Q _29512_/X _29922_/S VGND VGND VPWR VPWR _29923_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25045_ _24868_/X _33004_/Q _25059_/S VGND VGND VPWR VPWR _25046_/A sky130_fd_sc_hd__mux2_1
X_22257_ _34179_/Q _34115_/Q _34051_/Q _33987_/Q _22046_/X _22047_/X VGND VGND VPWR
+ VPWR _22257_/X sky130_fd_sc_hd__mux4_1
XFILLER_2_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21208_ _32869_/Q _32805_/Q _32741_/Q _32677_/Q _20887_/X _20888_/X VGND VGND VPWR
+ VPWR _21208_/X sky130_fd_sc_hd__mux4_1
XFILLER_219_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29853_ _35184_/Q _29410_/X _29859_/S VGND VGND VPWR VPWR _29854_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_1016 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22188_ _22188_/A _22188_/B _22188_/C _22188_/D VGND VGND VPWR VPWR _22189_/A sky130_fd_sc_hd__or4_4
XFILLER_78_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28804_ _34717_/Q _27056_/X _28808_/S VGND VGND VPWR VPWR _28805_/A sky130_fd_sc_hd__mux2_1
X_21139_ _33123_/Q _36003_/Q _32995_/Q _32931_/Q _20956_/X _20957_/X VGND VGND VPWR
+ VPWR _21139_/X sky130_fd_sc_hd__mux4_1
X_29784_ _29784_/A VGND VGND VPWR VPWR _35151_/D sky130_fd_sc_hd__clkbuf_1
X_26996_ _33924_/Q _23441_/X _27002_/S VGND VGND VPWR VPWR _26997_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_219_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_219_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28735_ _28735_/A VGND VGND VPWR VPWR _34685_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25947_ _31418_/B _26352_/B VGND VGND VPWR VPWR _26080_/S sky130_fd_sc_hd__nand2_8
XFILLER_58_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_463_CLK clkbuf_6_9__f_CLK/X VGND VGND VPWR VPWR _35564_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_247_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16680_ _32871_/Q _32807_/Q _32743_/Q _32679_/Q _16640_/X _16641_/X VGND VGND VPWR
+ VPWR _16680_/X sky130_fd_sc_hd__mux4_1
X_28666_ _28666_/A VGND VGND VPWR VPWR _34652_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25878_ _25878_/A VGND VGND VPWR VPWR _33396_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27617_ _34187_/Q _27199_/X _27629_/S VGND VGND VPWR VPWR _27618_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24829_ _24829_/A VGND VGND VPWR VPWR _32927_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28597_ _28597_/A VGND VGND VPWR VPWR _34620_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_215_CLK clkbuf_6_52__f_CLK/X VGND VGND VPWR VPWR _35213_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18350_ _20100_/A VGND VGND VPWR VPWR _18350_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_215_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27548_ _34154_/Q _27096_/X _27566_/S VGND VGND VPWR VPWR _27549_/A sky130_fd_sc_hd__mux2_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17301_ _17301_/A _17301_/B _17301_/C _17301_/D VGND VGND VPWR VPWR _17302_/A sky130_fd_sc_hd__or4_4
XFILLER_187_534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27479_ _27479_/A VGND VGND VPWR VPWR _34121_/D sky130_fd_sc_hd__clkbuf_1
X_18281_ _20159_/A VGND VGND VPWR VPWR _18281_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_159_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17232_ _34934_/Q _34870_/Q _34806_/Q _34742_/Q _17160_/X _17161_/X VGND VGND VPWR
+ VPWR _17232_/X sky130_fd_sc_hd__mux4_1
X_29218_ _34913_/Q _27069_/X _29234_/S VGND VGND VPWR VPWR _29219_/A sky130_fd_sc_hd__mux2_1
XFILLER_175_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30490_ _35486_/Q _29354_/X _30492_/S VGND VGND VPWR VPWR _30491_/A sky130_fd_sc_hd__mux2_1
XFILLER_243_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17163_ _17163_/A VGND VGND VPWR VPWR _17163_/X sky130_fd_sc_hd__clkbuf_4
X_29149_ _29149_/A VGND VGND VPWR VPWR _34880_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16114_ _33879_/Q _33815_/Q _33751_/Q _36055_/Q _16112_/X _16113_/X VGND VGND VPWR
+ VPWR _16114_/X sky130_fd_sc_hd__mux4_1
X_32160_ _35297_/CLK _32160_/D VGND VGND VPWR VPWR _32160_/Q sky130_fd_sc_hd__dfxtp_1
X_17094_ _17961_/A VGND VGND VPWR VPWR _17094_/X sky130_fd_sc_hd__buf_4
XFILLER_182_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31111_ _31111_/A VGND VGND VPWR VPWR _35780_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16045_ input70/X VGND VGND VPWR VPWR _17847_/A sky130_fd_sc_hd__buf_6
X_32091_ _35860_/CLK _32091_/D VGND VGND VPWR VPWR _32091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31042_ _31042_/A VGND VGND VPWR VPWR _35747_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_237_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19804_ _20157_/A VGND VGND VPWR VPWR _19804_/X sky130_fd_sc_hd__clkbuf_4
X_35850_ _36042_/CLK _35850_/D VGND VGND VPWR VPWR _35850_/Q sky130_fd_sc_hd__dfxtp_1
X_17996_ _17709_/X _17994_/X _17995_/X _17712_/X VGND VGND VPWR VPWR _17996_/X sky130_fd_sc_hd__a22o_1
X_34801_ _35439_/CLK _34801_/D VGND VGND VPWR VPWR _34801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19735_ _19729_/X _19734_/X _19451_/X VGND VGND VPWR VPWR _19743_/C sky130_fd_sc_hd__o21ba_1
X_35781_ _35843_/CLK _35781_/D VGND VGND VPWR VPWR _35781_/Q sky130_fd_sc_hd__dfxtp_1
X_16947_ _16943_/X _16946_/X _16812_/X VGND VGND VPWR VPWR _16948_/D sky130_fd_sc_hd__o21ba_1
X_32993_ _36129_/CLK _32993_/D VGND VGND VPWR VPWR _32993_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_454_CLK clkbuf_6_14__f_CLK/X VGND VGND VPWR VPWR _36140_/CLK sky130_fd_sc_hd__clkbuf_16
X_34732_ _34924_/CLK _34732_/D VGND VGND VPWR VPWR _34732_/Q sky130_fd_sc_hd__dfxtp_1
X_31944_ _23478_/X _36175_/Q _31948_/S VGND VGND VPWR VPWR _31945_/A sky130_fd_sc_hd__mux2_1
X_19666_ _19453_/X _19662_/X _19665_/X _19456_/X VGND VGND VPWR VPWR _19666_/X sky130_fd_sc_hd__a22o_1
X_16878_ _34412_/Q _36140_/Q _34284_/Q _34220_/Q _16876_/X _16877_/X VGND VGND VPWR
+ VPWR _16878_/X sky130_fd_sc_hd__mux4_1
X_18617_ _33373_/Q _33309_/Q _33245_/Q _33181_/Q _18302_/X _18303_/X VGND VGND VPWR
+ VPWR _18617_/X sky130_fd_sc_hd__mux4_1
X_34663_ _36137_/CLK _34663_/D VGND VGND VPWR VPWR _34663_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19597_ _34424_/Q _36152_/Q _34296_/Q _34232_/Q _19529_/X _19530_/X VGND VGND VPWR
+ VPWR _19597_/X sky130_fd_sc_hd__mux4_1
X_31875_ _23305_/X _36142_/Q _31885_/S VGND VGND VPWR VPWR _31876_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_206_CLK clkbuf_6_54__f_CLK/X VGND VGND VPWR VPWR _35657_/CLK sky130_fd_sc_hd__clkbuf_16
X_33614_ _34064_/CLK _33614_/D VGND VGND VPWR VPWR _33614_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18548_ _33883_/Q _33819_/Q _33755_/Q _36059_/Q _18412_/X _18413_/X VGND VGND VPWR
+ VPWR _18548_/X sky130_fd_sc_hd__mux4_1
XFILLER_52_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30826_ _30826_/A VGND VGND VPWR VPWR _35645_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_209_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34594_ _34594_/CLK _34594_/D VGND VGND VPWR VPWR _34594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33545_ _33673_/CLK _33545_/D VGND VGND VPWR VPWR _33545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18479_ _34137_/Q _34073_/Q _34009_/Q _33945_/Q _18309_/X _18311_/X VGND VGND VPWR
+ VPWR _18479_/X sky130_fd_sc_hd__mux4_1
XFILLER_178_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30757_ _30757_/A VGND VGND VPWR VPWR _35612_/D sky130_fd_sc_hd__clkbuf_1
X_20510_ _34707_/Q _34643_/Q _34579_/Q _34515_/Q _20298_/X _20299_/X VGND VGND VPWR
+ VPWR _20510_/X sky130_fd_sc_hd__mux4_1
X_33476_ _34182_/CLK _33476_/D VGND VGND VPWR VPWR _33476_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21490_ _21486_/X _21489_/X _21379_/X VGND VGND VPWR VPWR _21514_/A sky130_fd_sc_hd__o21ba_1
XFILLER_18_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30688_ _35580_/Q _29447_/X _30690_/S VGND VGND VPWR VPWR _30689_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35215_ _35664_/CLK _35215_/D VGND VGND VPWR VPWR _35215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20441_ _19458_/A _20439_/X _20440_/X _19463_/A VGND VGND VPWR VPWR _20441_/X sky130_fd_sc_hd__a22o_1
X_32427_ _33895_/CLK _32427_/D VGND VGND VPWR VPWR _32427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36195_ _36209_/CLK _36195_/D VGND VGND VPWR VPWR _36195_/Q sky130_fd_sc_hd__dfxtp_1
X_35146_ _35210_/CLK _35146_/D VGND VGND VPWR VPWR _35146_/Q sky130_fd_sc_hd__dfxtp_1
X_23160_ _23160_/A VGND VGND VPWR VPWR _32118_/D sky130_fd_sc_hd__clkbuf_1
X_20372_ _33423_/Q _33359_/Q _33295_/Q _33231_/Q _20133_/X _20134_/X VGND VGND VPWR
+ VPWR _20372_/X sky130_fd_sc_hd__mux4_1
X_32358_ _32552_/CLK _32358_/D VGND VGND VPWR VPWR _32358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22111_ _22464_/A VGND VGND VPWR VPWR _22111_/X sky130_fd_sc_hd__clkbuf_4
XTAP_7109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31309_ _31309_/A VGND VGND VPWR VPWR _35873_/D sky130_fd_sc_hd__clkbuf_1
X_35077_ _35718_/CLK _35077_/D VGND VGND VPWR VPWR _35077_/Q sky130_fd_sc_hd__dfxtp_1
X_23091_ _23223_/S VGND VGND VPWR VPWR _23110_/S sky130_fd_sc_hd__clkbuf_8
X_32289_ _32356_/CLK _32289_/D VGND VGND VPWR VPWR _32289_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34028_ _35627_/CLK _34028_/D VGND VGND VPWR VPWR _34028_/Q sky130_fd_sc_hd__dfxtp_1
X_22042_ _22038_/X _22041_/X _21765_/X VGND VGND VPWR VPWR _22043_/D sky130_fd_sc_hd__o21ba_1
XTAP_6419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1044 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26850_ _26850_/A VGND VGND VPWR VPWR _33854_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25801_ _25801_/A VGND VGND VPWR VPWR _33360_/D sky130_fd_sc_hd__clkbuf_1
X_26781_ _33822_/Q _23255_/X _26783_/S VGND VGND VPWR VPWR _26782_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23993_ _23993_/A VGND VGND VPWR VPWR _32539_/D sky130_fd_sc_hd__clkbuf_1
X_35979_ _35980_/CLK _35979_/D VGND VGND VPWR VPWR _35979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_214_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_445_CLK clkbuf_leaf_61_CLK/A VGND VGND VPWR VPWR _32877_/CLK sky130_fd_sc_hd__clkbuf_16
X_28520_ _28520_/A VGND VGND VPWR VPWR _34583_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_229_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25732_ _25732_/A VGND VGND VPWR VPWR _33327_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22944_ _22943_/X _32040_/Q _22947_/S VGND VGND VPWR VPWR _22945_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25663_ _24976_/X _33295_/Q _25667_/S VGND VGND VPWR VPWR _25664_/A sky130_fd_sc_hd__mux2_1
XFILLER_216_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28451_ _27745_/X _34551_/Q _28463_/S VGND VGND VPWR VPWR _28452_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22875_ _20660_/X _22873_/X _22874_/X _20672_/X VGND VGND VPWR VPWR _22875_/X sky130_fd_sc_hd__a22o_1
X_24614_ _23015_/X _32831_/Q _24630_/S VGND VGND VPWR VPWR _24615_/A sky130_fd_sc_hd__mux2_1
X_27402_ _34085_/Q _27081_/X _27410_/S VGND VGND VPWR VPWR _27403_/A sky130_fd_sc_hd__mux2_1
X_28382_ _27639_/X _34518_/Q _28400_/S VGND VGND VPWR VPWR _28383_/A sky130_fd_sc_hd__mux2_1
X_21826_ _34678_/Q _34614_/Q _34550_/Q _34486_/Q _21539_/X _21540_/X VGND VGND VPWR
+ VPWR _21826_/X sky130_fd_sc_hd__mux4_1
XFILLER_93_1020 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25594_ _24874_/X _33262_/Q _25604_/S VGND VGND VPWR VPWR _25595_/A sky130_fd_sc_hd__mux2_1
XFILLER_227_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27333_ _27333_/A VGND VGND VPWR VPWR _34052_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1015 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24545_ _24545_/A VGND VGND VPWR VPWR _32798_/D sky130_fd_sc_hd__clkbuf_1
X_21757_ _21753_/X _21754_/X _21755_/X _21756_/X VGND VGND VPWR VPWR _21757_/X sky130_fd_sc_hd__a22o_1
XFILLER_200_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_994 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20708_ _33623_/Q _33559_/Q _33495_/Q _33431_/Q _20584_/X _20587_/X VGND VGND VPWR
+ VPWR _20708_/X sky130_fd_sc_hd__mux4_1
XFILLER_12_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27264_ _27264_/A VGND VGND VPWR VPWR _34019_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24476_ _24524_/S VGND VGND VPWR VPWR _24495_/S sky130_fd_sc_hd__buf_4
XFILLER_211_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21688_ _21405_/X _21686_/X _21687_/X _21410_/X VGND VGND VPWR VPWR _21688_/X sky130_fd_sc_hd__a22o_1
XFILLER_106_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26215_ _24994_/X _33557_/Q _26215_/S VGND VGND VPWR VPWR _26216_/A sky130_fd_sc_hd__mux2_1
XFILLER_221_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29003_ _29003_/A VGND VGND VPWR VPWR _34811_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_10 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23427_ _32221_/Q _23426_/X _23451_/S VGND VGND VPWR VPWR _23428_/A sky130_fd_sc_hd__mux2_1
X_27195_ _27195_/A VGND VGND VPWR VPWR _33993_/D sky130_fd_sc_hd__clkbuf_1
X_20639_ _22434_/A VGND VGND VPWR VPWR _20639_/X sky130_fd_sc_hd__buf_4
XFILLER_221_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_913 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26146_ _26215_/S VGND VGND VPWR VPWR _26165_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_4_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23358_ _23358_/A VGND VGND VPWR VPWR _32195_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22309_ _22464_/A VGND VGND VPWR VPWR _22309_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_30_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26077_ _26077_/A VGND VGND VPWR VPWR _33491_/D sky130_fd_sc_hd__clkbuf_1
X_23289_ input11/X VGND VGND VPWR VPWR _23289_/X sky130_fd_sc_hd__buf_4
XFILLER_3_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29905_ _29905_/A VGND VGND VPWR VPWR _35208_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25028_ _24843_/X _32996_/Q _25038_/S VGND VGND VPWR VPWR _25029_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17850_ _17850_/A VGND VGND VPWR VPWR _17850_/X sky130_fd_sc_hd__buf_4
X_29836_ _35176_/Q _29385_/X _29838_/S VGND VGND VPWR VPWR _29837_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16801_ _34666_/Q _34602_/Q _34538_/Q _34474_/Q _16586_/X _16587_/X VGND VGND VPWR
+ VPWR _16801_/X sky130_fd_sc_hd__mux4_1
XTAP_6997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29767_ _29767_/A VGND VGND VPWR VPWR _35143_/D sky130_fd_sc_hd__clkbuf_1
X_17781_ _35654_/Q _35014_/Q _34374_/Q _33734_/Q _17497_/X _17498_/X VGND VGND VPWR
+ VPWR _17781_/X sky130_fd_sc_hd__mux4_1
XFILLER_219_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26979_ _33916_/Q _23414_/X _26981_/S VGND VGND VPWR VPWR _26980_/A sky130_fd_sc_hd__mux2_1
XFILLER_208_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_436_CLK clkbuf_6_33__f_CLK/X VGND VGND VPWR VPWR _36143_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_208_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19520_ _35638_/Q _34998_/Q _34358_/Q _33718_/Q _19444_/X _19445_/X VGND VGND VPWR
+ VPWR _19520_/X sky130_fd_sc_hd__mux4_1
XFILLER_235_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28718_ _34677_/Q _27131_/X _28734_/S VGND VGND VPWR VPWR _28719_/A sky130_fd_sc_hd__mux2_1
X_16732_ _16447_/X _16730_/X _16731_/X _16450_/X VGND VGND VPWR VPWR _16732_/X sky130_fd_sc_hd__a22o_1
X_29698_ _29698_/A VGND VGND VPWR VPWR _35110_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_1467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19451_ _20157_/A VGND VGND VPWR VPWR _19451_/X sky130_fd_sc_hd__buf_4
X_28649_ _28649_/A VGND VGND VPWR VPWR _34645_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16663_ _16452_/X _16661_/X _16662_/X _16457_/X VGND VGND VPWR VPWR _16663_/X sky130_fd_sc_hd__a22o_1
XFILLER_74_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18402_ _18391_/X _18395_/X _18399_/X _18401_/X VGND VGND VPWR VPWR _18402_/X sky130_fd_sc_hd__a22o_1
XFILLER_90_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31660_ _27797_/X _36040_/Q _31678_/S VGND VGND VPWR VPWR _31661_/A sky130_fd_sc_hd__mux2_1
X_19382_ _19376_/X _19381_/X _19098_/X VGND VGND VPWR VPWR _19390_/C sky130_fd_sc_hd__o21ba_1
X_16594_ _16590_/X _16593_/X _16459_/X VGND VGND VPWR VPWR _16595_/D sky130_fd_sc_hd__o21ba_1
XFILLER_43_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30611_ _35543_/Q _29333_/X _30627_/S VGND VGND VPWR VPWR _30612_/A sky130_fd_sc_hd__mux2_1
X_18333_ _18363_/A VGND VGND VPWR VPWR _20074_/A sky130_fd_sc_hd__buf_8
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31591_ _31591_/A VGND VGND VPWR VPWR _36007_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33330_ _34098_/CLK _33330_/D VGND VGND VPWR VPWR _33330_/Q sky130_fd_sc_hd__dfxtp_1
X_18264_ _35669_/Q _35029_/Q _34389_/Q _33749_/Q _16112_/X _16113_/X VGND VGND VPWR
+ VPWR _18264_/X sky130_fd_sc_hd__mux4_1
X_30542_ _30542_/A VGND VGND VPWR VPWR _35510_/D sky130_fd_sc_hd__clkbuf_1
X_17215_ _32118_/Q _32310_/Q _32374_/Q _35894_/Q _16927_/X _17068_/X VGND VGND VPWR
+ VPWR _17215_/X sky130_fd_sc_hd__mux4_1
X_33261_ _36077_/CLK _33261_/D VGND VGND VPWR VPWR _33261_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18195_ _18191_/X _18194_/X _17838_/A VGND VGND VPWR VPWR _18217_/A sky130_fd_sc_hd__o21ba_1
X_30473_ _30605_/S VGND VGND VPWR VPWR _30492_/S sky130_fd_sc_hd__buf_6
XFILLER_30_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35000_ _35769_/CLK _35000_/D VGND VGND VPWR VPWR _35000_/Q sky130_fd_sc_hd__dfxtp_1
X_32212_ _35703_/CLK _32212_/D VGND VGND VPWR VPWR _32212_/Q sky130_fd_sc_hd__dfxtp_1
X_17146_ _35636_/Q _34996_/Q _34356_/Q _33716_/Q _17144_/X _17145_/X VGND VGND VPWR
+ VPWR _17146_/X sky130_fd_sc_hd__mux4_1
XFILLER_190_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33192_ _36068_/CLK _33192_/D VGND VGND VPWR VPWR _33192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32143_ _32909_/CLK _32143_/D VGND VGND VPWR VPWR _32143_/Q sky130_fd_sc_hd__dfxtp_1
X_17077_ _35442_/Q _35378_/Q _35314_/Q _35250_/Q _16901_/X _16902_/X VGND VGND VPWR
+ VPWR _17077_/X sky130_fd_sc_hd__mux4_1
XFILLER_226_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16028_ _16018_/X _16023_/X _16026_/X _16027_/X VGND VGND VPWR VPWR _16028_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32074_ _36042_/CLK _32074_/D VGND VGND VPWR VPWR _32074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31025_ _31025_/A VGND VGND VPWR VPWR _35739_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35902_ _35902_/CLK _35902_/D VGND VGND VPWR VPWR _35902_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35833_ _35833_/CLK _35833_/D VGND VGND VPWR VPWR _35833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_1211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17979_ _33932_/Q _33868_/Q _33804_/Q _36108_/Q _17730_/X _17731_/X VGND VGND VPWR
+ VPWR _17979_/X sky130_fd_sc_hd__mux4_1
XFILLER_211_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_427_CLK clkbuf_6_35__f_CLK/X VGND VGND VPWR VPWR _35829_/CLK sky130_fd_sc_hd__clkbuf_16
X_19718_ _20210_/A VGND VGND VPWR VPWR _19718_/X sky130_fd_sc_hd__clkbuf_4
X_35764_ _35764_/CLK _35764_/D VGND VGND VPWR VPWR _35764_/Q sky130_fd_sc_hd__dfxtp_1
X_32976_ _36047_/CLK _32976_/D VGND VGND VPWR VPWR _32976_/Q sky130_fd_sc_hd__dfxtp_1
X_20990_ _20740_/X _20986_/X _20989_/X _20745_/X VGND VGND VPWR VPWR _20990_/X sky130_fd_sc_hd__a22o_1
XFILLER_81_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34715_ _34911_/CLK _34715_/D VGND VGND VPWR VPWR _34715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_996 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31927_ _23450_/X _36167_/Q _31927_/S VGND VGND VPWR VPWR _31928_/A sky130_fd_sc_hd__mux2_1
X_19649_ _19367_/X _19645_/X _19648_/X _19371_/X VGND VGND VPWR VPWR _19649_/X sky130_fd_sc_hd__a22o_1
X_35695_ _35697_/CLK _35695_/D VGND VGND VPWR VPWR _35695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_246_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34646_ _34647_/CLK _34646_/D VGND VGND VPWR VPWR _34646_/Q sky130_fd_sc_hd__dfxtp_1
X_22660_ _34702_/Q _34638_/Q _34574_/Q _34510_/Q _22598_/X _22599_/X VGND VGND VPWR
+ VPWR _22660_/X sky130_fd_sc_hd__mux4_1
XFILLER_179_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31858_ _23280_/X _36134_/Q _31864_/S VGND VGND VPWR VPWR _31859_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21611_ _21611_/A VGND VGND VPWR VPWR _21611_/X sky130_fd_sc_hd__buf_4
XFILLER_209_1162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30809_ _35637_/Q input25/X _30825_/S VGND VGND VPWR VPWR _30810_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34577_ _36175_/CLK _34577_/D VGND VGND VPWR VPWR _34577_/Q sky130_fd_sc_hd__dfxtp_1
X_22591_ _35724_/Q _32235_/Q _35596_/Q _35532_/Q _22270_/X _22271_/X VGND VGND VPWR
+ VPWR _22591_/X sky130_fd_sc_hd__mux4_1
X_31789_ _31789_/A VGND VGND VPWR VPWR _36101_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24330_ _24330_/A VGND VGND VPWR VPWR _32696_/D sky130_fd_sc_hd__clkbuf_1
X_33528_ _35641_/CLK _33528_/D VGND VGND VPWR VPWR _33528_/Q sky130_fd_sc_hd__dfxtp_1
X_21542_ _35182_/Q _35118_/Q _35054_/Q _32174_/Q _21257_/X _21258_/X VGND VGND VPWR
+ VPWR _21542_/X sky130_fd_sc_hd__mux4_1
XFILLER_181_1387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24261_ _24261_/A VGND VGND VPWR VPWR _32663_/D sky130_fd_sc_hd__clkbuf_1
X_33459_ _34098_/CLK _33459_/D VGND VGND VPWR VPWR _33459_/Q sky130_fd_sc_hd__dfxtp_1
X_21473_ _34668_/Q _34604_/Q _34540_/Q _34476_/Q _21186_/X _21187_/X VGND VGND VPWR
+ VPWR _21473_/X sky130_fd_sc_hd__mux4_1
XFILLER_14_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_6_51__f_CLK clkbuf_5_25_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_51__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_26000_ _26000_/A VGND VGND VPWR VPWR _33454_/D sky130_fd_sc_hd__clkbuf_1
X_23212_ _23212_/A VGND VGND VPWR VPWR _32143_/D sky130_fd_sc_hd__clkbuf_1
X_20424_ _34960_/Q _34896_/Q _34832_/Q _34768_/Q _20166_/X _20167_/X VGND VGND VPWR
+ VPWR _20424_/X sky130_fd_sc_hd__mux4_1
XFILLER_153_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36178_ _36180_/CLK _36178_/D VGND VGND VPWR VPWR _36178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24192_ _24192_/A VGND VGND VPWR VPWR _32632_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35129_ _35191_/CLK _35129_/D VGND VGND VPWR VPWR _35129_/Q sky130_fd_sc_hd__dfxtp_1
X_23143_ _23143_/A VGND VGND VPWR VPWR _32110_/D sky130_fd_sc_hd__clkbuf_1
X_20355_ _18281_/X _20353_/X _20354_/X _18291_/X VGND VGND VPWR VPWR _20355_/X sky130_fd_sc_hd__a22o_1
XFILLER_20_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27951_ _27804_/X _34314_/Q _27965_/S VGND VGND VPWR VPWR _27952_/A sky130_fd_sc_hd__mux2_1
XTAP_6205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23074_ _23073_/X _32082_/Q _23083_/S VGND VGND VPWR VPWR _23075_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20286_ _20286_/A VGND VGND VPWR VPWR _20286_/X sky130_fd_sc_hd__buf_6
XTAP_6227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26902_ _33879_/Q _23234_/X _26918_/S VGND VGND VPWR VPWR _26903_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22025_ _22020_/X _22022_/X _22023_/X _22024_/X VGND VGND VPWR VPWR _22025_/X sky130_fd_sc_hd__a22o_1
XTAP_6249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27882_ _27882_/A VGND VGND VPWR VPWR _34281_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29621_ _35074_/Q _29466_/X _29631_/S VGND VGND VPWR VPWR _29622_/A sky130_fd_sc_hd__mux2_1
XTAP_4803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26833_ _26833_/A VGND VGND VPWR VPWR _33846_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_1480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_418_CLK clkbuf_6_33__f_CLK/X VGND VGND VPWR VPWR _35633_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29552_ _35041_/Q _29364_/X _29568_/S VGND VGND VPWR VPWR _29553_/A sky130_fd_sc_hd__mux2_1
X_23976_ _23976_/A VGND VGND VPWR VPWR _32532_/D sky130_fd_sc_hd__clkbuf_1
X_26764_ _26896_/S VGND VGND VPWR VPWR _26783_/S sky130_fd_sc_hd__buf_6
XFILLER_99_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28503_ _27822_/X _34576_/Q _28505_/S VGND VGND VPWR VPWR _28504_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_1164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25715_ _25715_/A VGND VGND VPWR VPWR _33319_/D sky130_fd_sc_hd__clkbuf_1
X_22927_ _22927_/A VGND VGND VPWR VPWR _32034_/D sky130_fd_sc_hd__clkbuf_1
X_29483_ _29483_/A VGND VGND VPWR VPWR _35015_/D sky130_fd_sc_hd__clkbuf_1
X_26695_ _33781_/Q _23393_/X _26711_/S VGND VGND VPWR VPWR _26696_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28434_ _27720_/X _34543_/Q _28442_/S VGND VGND VPWR VPWR _28435_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25646_ _24951_/X _33287_/Q _25646_/S VGND VGND VPWR VPWR _25647_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22858_ _21753_/A _22856_/X _22857_/X _21756_/A VGND VGND VPWR VPWR _22858_/X sky130_fd_sc_hd__a22o_1
XFILLER_32_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_882 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21809_ _22515_/A VGND VGND VPWR VPWR _21809_/X sky130_fd_sc_hd__buf_6
X_28365_ _28365_/A VGND VGND VPWR VPWR _34510_/D sky130_fd_sc_hd__clkbuf_1
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25577_ _24849_/X _33254_/Q _25583_/S VGND VGND VPWR VPWR _25578_/A sky130_fd_sc_hd__mux2_1
X_22789_ _33683_/Q _33619_/Q _33555_/Q _33491_/Q _22506_/X _22507_/X VGND VGND VPWR
+ VPWR _22789_/X sky130_fd_sc_hd__mux4_1
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24528_ _22879_/X _32790_/Q _24546_/S VGND VGND VPWR VPWR _24529_/A sky130_fd_sc_hd__mux2_1
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27316_ _27316_/A VGND VGND VPWR VPWR _34044_/D sky130_fd_sc_hd__clkbuf_1
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28296_ _28296_/A VGND VGND VPWR VPWR _34477_/D sky130_fd_sc_hd__clkbuf_1
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_885 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27247_ _27247_/A VGND VGND VPWR VPWR _34011_/D sky130_fd_sc_hd__clkbuf_1
X_24459_ _24459_/A VGND VGND VPWR VPWR _32757_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_902 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17000_ _35632_/Q _34992_/Q _34352_/Q _33712_/Q _16791_/X _16792_/X VGND VGND VPWR
+ VPWR _17000_/X sky130_fd_sc_hd__mux4_1
XFILLER_201_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27178_ _33988_/Q _27177_/X _27187_/S VGND VGND VPWR VPWR _27179_/A sky130_fd_sc_hd__mux2_1
XFILLER_197_1350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26129_ _26129_/A VGND VGND VPWR VPWR _33515_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18951_ _35430_/Q _35366_/Q _35302_/Q _35238_/Q _18848_/X _18849_/X VGND VGND VPWR
+ VPWR _18951_/X sky130_fd_sc_hd__mux4_1
XFILLER_141_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17902_ _17898_/X _17901_/X _17871_/X VGND VGND VPWR VPWR _17903_/D sky130_fd_sc_hd__o21ba_1
XFILLER_140_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18882_ _35428_/Q _35364_/Q _35300_/Q _35236_/Q _18848_/X _18849_/X VGND VGND VPWR
+ VPWR _18882_/X sky130_fd_sc_hd__mux4_1
XTAP_6750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17833_ _17833_/A VGND VGND VPWR VPWR _17833_/X sky130_fd_sc_hd__buf_4
XFILLER_121_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29819_ _29930_/S VGND VGND VPWR VPWR _29838_/S sky130_fd_sc_hd__buf_6
XTAP_6783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_409_CLK clkbuf_6_32__f_CLK/X VGND VGND VPWR VPWR _35697_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_187_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32830_ _32894_/CLK _32830_/D VGND VGND VPWR VPWR _32830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_952 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17764_ _17760_/X _17763_/X _17485_/X VGND VGND VPWR VPWR _17796_/A sky130_fd_sc_hd__o21ba_2
XFILLER_187_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19503_ _34166_/Q _34102_/Q _34038_/Q _33974_/Q _19393_/X _19394_/X VGND VGND VPWR
+ VPWR _19503_/X sky130_fd_sc_hd__mux4_1
XFILLER_75_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16715_ _17774_/A VGND VGND VPWR VPWR _16715_/X sky130_fd_sc_hd__clkbuf_4
X_32761_ _35895_/CLK _32761_/D VGND VGND VPWR VPWR _32761_/Q sky130_fd_sc_hd__dfxtp_1
X_17695_ _32644_/Q _32580_/Q _32516_/Q _35972_/Q _17629_/X _17413_/X VGND VGND VPWR
+ VPWR _17695_/X sky130_fd_sc_hd__mux4_1
XFILLER_74_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34500_ _34693_/CLK _34500_/D VGND VGND VPWR VPWR _34500_/Q sky130_fd_sc_hd__dfxtp_1
X_31712_ _31712_/A VGND VGND VPWR VPWR _36064_/D sky130_fd_sc_hd__clkbuf_1
X_19434_ _32628_/Q _32564_/Q _32500_/Q _35956_/Q _19223_/X _19360_/X VGND VGND VPWR
+ VPWR _19434_/X sky130_fd_sc_hd__mux4_1
XFILLER_228_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35480_ _35544_/CLK _35480_/D VGND VGND VPWR VPWR _35480_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16646_ _35686_/Q _32193_/Q _35558_/Q _35494_/Q _16611_/X _16612_/X VGND VGND VPWR
+ VPWR _16646_/X sky130_fd_sc_hd__mux4_1
XFILLER_62_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32692_ _32904_/CLK _32692_/D VGND VGND VPWR VPWR _32692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34431_ _36161_/CLK _34431_/D VGND VGND VPWR VPWR _34431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31643_ _27773_/X _36032_/Q _31657_/S VGND VGND VPWR VPWR _31644_/A sky130_fd_sc_hd__mux2_1
X_19365_ _20210_/A VGND VGND VPWR VPWR _19365_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_204_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16577_ _16361_/X _16575_/X _16576_/X _16365_/X VGND VGND VPWR VPWR _16577_/X sky130_fd_sc_hd__a22o_1
XFILLER_206_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18316_ _18297_/X _18313_/X _18315_/X VGND VGND VPWR VPWR _18406_/A sky130_fd_sc_hd__o21ba_1
XFILLER_124_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34362_ _35644_/CLK _34362_/D VGND VGND VPWR VPWR _34362_/Q sky130_fd_sc_hd__dfxtp_1
X_31574_ _31574_/A VGND VGND VPWR VPWR _35999_/D sky130_fd_sc_hd__clkbuf_1
X_19296_ _19014_/X _19292_/X _19295_/X _19018_/X VGND VGND VPWR VPWR _19296_/X sky130_fd_sc_hd__a22o_1
X_36101_ _36101_/CLK _36101_/D VGND VGND VPWR VPWR _36101_/Q sky130_fd_sc_hd__dfxtp_1
X_33313_ _33697_/CLK _33313_/D VGND VGND VPWR VPWR _33313_/Q sky130_fd_sc_hd__dfxtp_1
X_18247_ _18247_/A _18247_/B _18247_/C _18247_/D VGND VGND VPWR VPWR _18248_/A sky130_fd_sc_hd__or4_4
XFILLER_15_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30525_ _30525_/A VGND VGND VPWR VPWR _35502_/D sky130_fd_sc_hd__clkbuf_1
X_34293_ _35187_/CLK _34293_/D VGND VGND VPWR VPWR _34293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36032_ _36033_/CLK _36032_/D VGND VGND VPWR VPWR _36032_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33244_ _36188_/CLK _33244_/D VGND VGND VPWR VPWR _33244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30456_ _35470_/Q _29503_/X _30462_/S VGND VGND VPWR VPWR _30457_/A sky130_fd_sc_hd__mux2_1
X_18178_ _16001_/X _18176_/X _18177_/X _16007_/X VGND VGND VPWR VPWR _18178_/X sky130_fd_sc_hd__a22o_1
XFILLER_239_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_1412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17129_ _33396_/Q _33332_/Q _33268_/Q _33204_/Q _17127_/X _17128_/X VGND VGND VPWR
+ VPWR _17129_/X sky130_fd_sc_hd__mux4_1
X_33175_ _36054_/CLK _33175_/D VGND VGND VPWR VPWR _33175_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30387_ _35437_/Q _29401_/X _30399_/S VGND VGND VPWR VPWR _30388_/A sky130_fd_sc_hd__mux2_1
XFILLER_239_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20140_ _32648_/Q _32584_/Q _32520_/Q _35976_/Q _19929_/X _20066_/X VGND VGND VPWR
+ VPWR _20140_/X sky130_fd_sc_hd__mux4_1
XFILLER_137_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32126_ _35903_/CLK _32126_/D VGND VGND VPWR VPWR _32126_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_990 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20071_ _20071_/A VGND VGND VPWR VPWR _20071_/X sky130_fd_sc_hd__clkbuf_4
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32057_ _35835_/CLK _32057_/D VGND VGND VPWR VPWR _32057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31008_ _35732_/Q input59/X _31010_/S VGND VGND VPWR VPWR _31009_/A sky130_fd_sc_hd__mux2_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23830_ _23067_/X _32400_/Q _23832_/S VGND VGND VPWR VPWR _23831_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35816_ _35817_/CLK _35816_/D VGND VGND VPWR VPWR _35816_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35747_ _35747_/CLK _35747_/D VGND VGND VPWR VPWR _35747_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23761_ _22965_/X _32367_/Q _23769_/S VGND VGND VPWR VPWR _23762_/A sky130_fd_sc_hd__mux2_1
X_32959_ _35903_/CLK _32959_/D VGND VGND VPWR VPWR _32959_/Q sky130_fd_sc_hd__dfxtp_1
X_20973_ _22536_/A VGND VGND VPWR VPWR _20973_/X sky130_fd_sc_hd__buf_4
X_25500_ _25500_/A VGND VGND VPWR VPWR _33217_/D sky130_fd_sc_hd__clkbuf_1
X_22712_ _22708_/X _22711_/X _22446_/X _22447_/X VGND VGND VPWR VPWR _22727_/B sky130_fd_sc_hd__o211a_2
XFILLER_26_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26480_ _33682_/Q _23487_/X _26486_/S VGND VGND VPWR VPWR _26481_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23692_ _23067_/X _32336_/Q _23694_/S VGND VGND VPWR VPWR _23693_/A sky130_fd_sc_hd__mux2_1
X_35678_ _35743_/CLK _35678_/D VGND VGND VPWR VPWR _35678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25431_ _25431_/A VGND VGND VPWR VPWR _33184_/D sky130_fd_sc_hd__clkbuf_1
X_22643_ _33934_/Q _33870_/Q _33806_/Q _36110_/Q _22330_/X _22331_/X VGND VGND VPWR
+ VPWR _22643_/X sky130_fd_sc_hd__mux4_1
X_34629_ _34694_/CLK _34629_/D VGND VGND VPWR VPWR _34629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_222_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25362_ _33153_/Q _23432_/X _25374_/S VGND VGND VPWR VPWR _25363_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28150_ _28150_/A VGND VGND VPWR VPWR _34408_/D sky130_fd_sc_hd__clkbuf_1
X_22574_ _22574_/A VGND VGND VPWR VPWR _36235_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27101_ _33963_/Q _27100_/X _27125_/S VGND VGND VPWR VPWR _27102_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24313_ _24313_/A VGND VGND VPWR VPWR _32688_/D sky130_fd_sc_hd__clkbuf_1
X_28081_ _28108_/S VGND VGND VPWR VPWR _28100_/S sky130_fd_sc_hd__clkbuf_4
X_21525_ _33134_/Q _36014_/Q _33006_/Q _32942_/Q _21309_/X _21310_/X VGND VGND VPWR
+ VPWR _21525_/X sky130_fd_sc_hd__mux4_1
XFILLER_103_1108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25293_ _33120_/Q _23261_/X _25311_/S VGND VGND VPWR VPWR _25294_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27032_ _27032_/A VGND VGND VPWR VPWR _33941_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24244_ _24244_/A VGND VGND VPWR VPWR _32657_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21456_ _22515_/A VGND VGND VPWR VPWR _21456_/X sky130_fd_sc_hd__buf_4
XFILLER_5_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_946 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20407_ _33168_/Q _36048_/Q _33040_/Q _32976_/Q _18332_/X _19461_/A VGND VGND VPWR
+ VPWR _20407_/X sky130_fd_sc_hd__mux4_1
XFILLER_120_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24175_ _24175_/A VGND VGND VPWR VPWR _32624_/D sky130_fd_sc_hd__clkbuf_1
X_21387_ _22446_/A VGND VGND VPWR VPWR _21387_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_107_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_927 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23126_ _23126_/A VGND VGND VPWR VPWR _32102_/D sky130_fd_sc_hd__clkbuf_1
X_20338_ _20338_/A VGND VGND VPWR VPWR _32461_/D sky130_fd_sc_hd__clkbuf_4
X_28983_ _34802_/Q _27121_/X _28985_/S VGND VGND VPWR VPWR _28984_/A sky130_fd_sc_hd__mux2_1
XTAP_6002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27934_ _27779_/X _34306_/Q _27944_/S VGND VGND VPWR VPWR _27935_/A sky130_fd_sc_hd__mux2_1
X_23057_ _23057_/A VGND VGND VPWR VPWR _32076_/D sky130_fd_sc_hd__clkbuf_1
X_20269_ _34443_/Q _36171_/Q _34315_/Q _34251_/Q _20235_/X _20236_/X VGND VGND VPWR
+ VPWR _20269_/X sky130_fd_sc_hd__mux4_1
XTAP_6046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22008_ _33404_/Q _33340_/Q _33276_/Q _33212_/Q _21727_/X _21728_/X VGND VGND VPWR
+ VPWR _22008_/X sky130_fd_sc_hd__mux4_1
XFILLER_103_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27865_ _27677_/X _34273_/Q _27881_/S VGND VGND VPWR VPWR _27866_/A sky130_fd_sc_hd__mux2_1
XFILLER_209_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29604_ _35066_/Q _29441_/X _29610_/S VGND VGND VPWR VPWR _29605_/A sky130_fd_sc_hd__mux2_1
XTAP_5378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26816_ _26816_/A VGND VGND VPWR VPWR _33838_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27796_ _27796_/A VGND VGND VPWR VPWR _34247_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29535_ _35033_/Q _29339_/X _29547_/S VGND VGND VPWR VPWR _29536_/A sky130_fd_sc_hd__mux2_1
XTAP_3943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26747_ _33806_/Q _23475_/X _26753_/S VGND VGND VPWR VPWR _26748_/A sky130_fd_sc_hd__mux2_1
XTAP_4688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23959_ _23055_/X _32524_/Q _23969_/S VGND VGND VPWR VPWR _23960_/A sky130_fd_sc_hd__mux2_1
XTAP_3954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16500_ _17912_/A VGND VGND VPWR VPWR _16500_/X sky130_fd_sc_hd__buf_4
XFILLER_232_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17480_ _17833_/A VGND VGND VPWR VPWR _17480_/X sky130_fd_sc_hd__buf_4
X_29466_ input39/X VGND VGND VPWR VPWR _29466_/X sky130_fd_sc_hd__buf_2
XTAP_3998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26678_ _33773_/Q _23302_/X _26690_/S VGND VGND VPWR VPWR _26679_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16431_ _32096_/Q _32288_/Q _32352_/Q _35872_/Q _16221_/X _16362_/X VGND VGND VPWR
+ VPWR _16431_/X sky130_fd_sc_hd__mux4_1
X_28417_ _27695_/X _34535_/Q _28421_/S VGND VGND VPWR VPWR _28418_/A sky130_fd_sc_hd__mux2_1
X_25629_ _25629_/A VGND VGND VPWR VPWR _33278_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29397_ _29397_/A VGND VGND VPWR VPWR _34987_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19150_ _34156_/Q _34092_/Q _34028_/Q _33964_/Q _19040_/X _19041_/X VGND VGND VPWR
+ VPWR _19150_/X sky130_fd_sc_hd__mux4_1
XFILLER_34_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28348_ _28348_/A VGND VGND VPWR VPWR _34502_/D sky130_fd_sc_hd__clkbuf_1
X_16362_ _17774_/A VGND VGND VPWR VPWR _16362_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_31_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18101_ _17905_/X _18099_/X _18100_/X _17910_/X VGND VGND VPWR VPWR _18101_/X sky130_fd_sc_hd__a22o_1
XFILLER_188_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16293_ _35676_/Q _32182_/Q _35548_/Q _35484_/Q _16258_/X _16259_/X VGND VGND VPWR
+ VPWR _16293_/X sky130_fd_sc_hd__mux4_1
X_19081_ _32618_/Q _32554_/Q _32490_/Q _35946_/Q _18870_/X _19007_/X VGND VGND VPWR
+ VPWR _19081_/X sky130_fd_sc_hd__mux4_1
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28279_ _28279_/A VGND VGND VPWR VPWR _34469_/D sky130_fd_sc_hd__clkbuf_1
X_18032_ _17859_/X _18030_/X _18031_/X _17862_/X VGND VGND VPWR VPWR _18032_/X sky130_fd_sc_hd__a22o_1
X_30310_ _30310_/A VGND VGND VPWR VPWR _35400_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31290_ _31290_/A VGND VGND VPWR VPWR _35864_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30241_ _35368_/Q _29385_/X _30243_/S VGND VGND VPWR VPWR _30242_/A sky130_fd_sc_hd__mux2_1
XFILLER_236_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30172_ _30172_/A VGND VGND VPWR VPWR _35335_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19983_ _34947_/Q _34883_/Q _34819_/Q _34755_/Q _19813_/X _19814_/X VGND VGND VPWR
+ VPWR _19983_/X sky130_fd_sc_hd__mux4_1
XFILLER_140_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18934_ _18800_/X _18932_/X _18933_/X _18803_/X VGND VGND VPWR VPWR _18934_/X sky130_fd_sc_hd__a22o_1
X_34980_ _35625_/CLK _34980_/D VGND VGND VPWR VPWR _34980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33931_ _36106_/CLK _33931_/D VGND VGND VPWR VPWR _33931_/Q sky130_fd_sc_hd__dfxtp_1
X_18865_ _18793_/X _18863_/X _18864_/X _18798_/X VGND VGND VPWR VPWR _18865_/X sky130_fd_sc_hd__a22o_1
XTAP_6580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17816_ _17704_/X _17814_/X _17815_/X _17707_/X VGND VGND VPWR VPWR _17816_/X sky130_fd_sc_hd__a22o_1
XFILLER_95_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33862_ _34177_/CLK _33862_/D VGND VGND VPWR VPWR _33862_/Q sky130_fd_sc_hd__dfxtp_1
X_18796_ _33634_/Q _33570_/Q _33506_/Q _33442_/Q _18794_/X _18795_/X VGND VGND VPWR
+ VPWR _18796_/X sky130_fd_sc_hd__mux4_1
XFILLER_55_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35601_ _35729_/CLK _35601_/D VGND VGND VPWR VPWR _35601_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32813_ _32877_/CLK _32813_/D VGND VGND VPWR VPWR _32813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_236_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17747_ _17709_/X _17745_/X _17746_/X _17712_/X VGND VGND VPWR VPWR _17747_/X sky130_fd_sc_hd__a22o_1
X_33793_ _36097_/CLK _33793_/D VGND VGND VPWR VPWR _33793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_1132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35532_ _35596_/CLK _35532_/D VGND VGND VPWR VPWR _35532_/Q sky130_fd_sc_hd__dfxtp_1
X_32744_ _32808_/CLK _32744_/D VGND VGND VPWR VPWR _32744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17678_ _17674_/X _17677_/X _17504_/X VGND VGND VPWR VPWR _17686_/C sky130_fd_sc_hd__o21ba_1
XFILLER_23_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19417_ _19100_/X _19415_/X _19416_/X _19103_/X VGND VGND VPWR VPWR _19417_/X sky130_fd_sc_hd__a22o_1
X_35463_ _35463_/CLK _35463_/D VGND VGND VPWR VPWR _35463_/Q sky130_fd_sc_hd__dfxtp_1
X_16629_ _33638_/Q _33574_/Q _33510_/Q _33446_/Q _16494_/X _16495_/X VGND VGND VPWR
+ VPWR _16629_/X sky130_fd_sc_hd__mux4_1
X_32675_ _32871_/CLK _32675_/D VGND VGND VPWR VPWR _32675_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34414_ _35822_/CLK _34414_/D VGND VGND VPWR VPWR _34414_/Q sky130_fd_sc_hd__dfxtp_1
X_19348_ _19105_/X _19346_/X _19347_/X _19110_/X VGND VGND VPWR VPWR _19348_/X sky130_fd_sc_hd__a22o_1
X_31626_ _27748_/X _36024_/Q _31636_/S VGND VGND VPWR VPWR _31627_/A sky130_fd_sc_hd__mux2_1
X_35394_ _35715_/CLK _35394_/D VGND VGND VPWR VPWR _35394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34345_ _35559_/CLK _34345_/D VGND VGND VPWR VPWR _34345_/Q sky130_fd_sc_hd__dfxtp_1
X_31557_ _27646_/X _35991_/Q _31573_/S VGND VGND VPWR VPWR _31558_/A sky130_fd_sc_hd__mux2_1
XFILLER_176_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19279_ _19275_/X _19278_/X _19112_/X VGND VGND VPWR VPWR _19280_/D sky130_fd_sc_hd__o21ba_1
XFILLER_175_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21310_ _22507_/A VGND VGND VPWR VPWR _21310_/X sky130_fd_sc_hd__clkbuf_4
X_30508_ _30508_/A VGND VGND VPWR VPWR _35494_/D sky130_fd_sc_hd__clkbuf_1
X_22290_ _22152_/X _22288_/X _22289_/X _22157_/X VGND VGND VPWR VPWR _22290_/X sky130_fd_sc_hd__a22o_1
XFILLER_117_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34276_ _34405_/CLK _34276_/D VGND VGND VPWR VPWR _34276_/Q sky130_fd_sc_hd__dfxtp_1
X_31488_ _31488_/A VGND VGND VPWR VPWR _35958_/D sky130_fd_sc_hd__clkbuf_1
X_36015_ _36015_/CLK _36015_/D VGND VGND VPWR VPWR _36015_/Q sky130_fd_sc_hd__dfxtp_1
X_33227_ _33420_/CLK _33227_/D VGND VGND VPWR VPWR _33227_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21241_ _22434_/A VGND VGND VPWR VPWR _21241_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_11_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30439_ _35462_/Q _29478_/X _30441_/S VGND VGND VPWR VPWR _30440_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33158_ _36038_/CLK _33158_/D VGND VGND VPWR VPWR _33158_/Q sky130_fd_sc_hd__dfxtp_1
X_21172_ _33124_/Q _36004_/Q _32996_/Q _32932_/Q _20956_/X _20957_/X VGND VGND VPWR
+ VPWR _21172_/X sky130_fd_sc_hd__mux4_1
XFILLER_116_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20123_ _19806_/X _20121_/X _20122_/X _19809_/X VGND VGND VPWR VPWR _20123_/X sky130_fd_sc_hd__a22o_1
XFILLER_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32109_ _35951_/CLK _32109_/D VGND VGND VPWR VPWR _32109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33089_ _35646_/CLK _33089_/D VGND VGND VPWR VPWR _33089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25980_ _24846_/X _33445_/Q _25988_/S VGND VGND VPWR VPWR _25981_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20054_ _19811_/X _20052_/X _20053_/X _19816_/X VGND VGND VPWR VPWR _20054_/X sky130_fd_sc_hd__a22o_1
X_24931_ _24930_/X _32960_/Q _24952_/S VGND VGND VPWR VPWR _24932_/A sky130_fd_sc_hd__mux2_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27650_ _27649_/X _34200_/Q _27671_/S VGND VGND VPWR VPWR _27651_/A sky130_fd_sc_hd__mux2_1
X_24862_ _24995_/S VGND VGND VPWR VPWR _24890_/S sky130_fd_sc_hd__buf_4
XTAP_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_1180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26601_ _26601_/A VGND VGND VPWR VPWR _33738_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_861 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23813_ _23840_/S VGND VGND VPWR VPWR _23832_/S sky130_fd_sc_hd__buf_4
XTAP_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24793_ _24793_/A VGND VGND VPWR VPWR _32916_/D sky130_fd_sc_hd__clkbuf_1
X_27581_ _34170_/Q _27146_/X _27587_/S VGND VGND VPWR VPWR _27582_/A sky130_fd_sc_hd__mux2_1
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29320_ _34962_/Q _27220_/X _29326_/S VGND VGND VPWR VPWR _29321_/A sky130_fd_sc_hd__mux2_1
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26532_ _26622_/S VGND VGND VPWR VPWR _26551_/S sky130_fd_sc_hd__buf_4
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23744_ _22940_/X _32359_/Q _23748_/S VGND VGND VPWR VPWR _23745_/A sky130_fd_sc_hd__mux2_1
X_20956_ _22506_/A VGND VGND VPWR VPWR _20956_/X sky130_fd_sc_hd__buf_4
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_1355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29251_ _34929_/Q _27118_/X _29255_/S VGND VGND VPWR VPWR _29252_/A sky130_fd_sc_hd__mux2_1
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26463_ _26463_/A VGND VGND VPWR VPWR _33673_/D sky130_fd_sc_hd__clkbuf_1
X_23675_ _23702_/S VGND VGND VPWR VPWR _23694_/S sky130_fd_sc_hd__buf_4
X_20887_ _22433_/A VGND VGND VPWR VPWR _20887_/X sky130_fd_sc_hd__buf_4
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_1390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28202_ _27776_/X _34433_/Q _28214_/S VGND VGND VPWR VPWR _28203_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22626_ _35469_/Q _35405_/Q _35341_/Q _35277_/Q _22560_/X _22561_/X VGND VGND VPWR
+ VPWR _22626_/X sky130_fd_sc_hd__mux4_1
X_25414_ _25414_/A VGND VGND VPWR VPWR _33176_/D sky130_fd_sc_hd__clkbuf_1
X_29182_ _29182_/A VGND VGND VPWR VPWR _34896_/D sky130_fd_sc_hd__clkbuf_1
X_26394_ _33641_/Q _23289_/X _26394_/S VGND VGND VPWR VPWR _26395_/A sky130_fd_sc_hd__mux2_1
XFILLER_224_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25345_ _33145_/Q _23405_/X _25353_/S VGND VGND VPWR VPWR _25346_/A sky130_fd_sc_hd__mux2_1
X_28133_ _27673_/X _34400_/Q _28151_/S VGND VGND VPWR VPWR _28134_/A sky130_fd_sc_hd__mux2_1
X_22557_ _35723_/Q _32234_/Q _35595_/Q _35531_/Q _22270_/X _22271_/X VGND VGND VPWR
+ VPWR _22557_/X sky130_fd_sc_hd__mux4_1
XFILLER_107_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21508_ _35181_/Q _35117_/Q _35053_/Q _32173_/Q _21257_/X _21258_/X VGND VGND VPWR
+ VPWR _21508_/X sky130_fd_sc_hd__mux4_1
X_25276_ _33112_/Q _23237_/X _25290_/S VGND VGND VPWR VPWR _25277_/A sky130_fd_sc_hd__mux2_1
XFILLER_181_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28064_ _28064_/A VGND VGND VPWR VPWR _34367_/D sky130_fd_sc_hd__clkbuf_1
X_22488_ _22484_/X _22487_/X _22446_/X _22447_/X VGND VGND VPWR VPWR _22503_/B sky130_fd_sc_hd__o211a_2
XFILLER_166_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27015_ _33933_/Q _23472_/X _27023_/S VGND VGND VPWR VPWR _27016_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24227_ _32649_/Q _23460_/X _24243_/S VGND VGND VPWR VPWR _24228_/A sky130_fd_sc_hd__mux2_1
X_21439_ _21400_/X _21437_/X _21438_/X _21403_/X VGND VGND VPWR VPWR _21439_/X sky130_fd_sc_hd__a22o_1
XFILLER_123_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24158_ _24158_/A VGND VGND VPWR VPWR _32616_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23109_ _23109_/A VGND VGND VPWR VPWR _32094_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24089_ _23046_/X _32585_/Q _24105_/S VGND VGND VPWR VPWR _24090_/A sky130_fd_sc_hd__mux2_1
X_16980_ _16980_/A _16980_/B _16980_/C _16980_/D VGND VGND VPWR VPWR _16981_/A sky130_fd_sc_hd__or4_4
X_28966_ _29056_/S VGND VGND VPWR VPWR _28985_/S sky130_fd_sc_hd__buf_4
XFILLER_150_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27917_ _27754_/X _34298_/Q _27923_/S VGND VGND VPWR VPWR _27918_/A sky130_fd_sc_hd__mux2_1
XTAP_5131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28897_ _34761_/Q _27193_/X _28913_/S VGND VGND VPWR VPWR _28898_/A sky130_fd_sc_hd__mux2_1
XTAP_5142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1086 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18650_ _33886_/Q _33822_/Q _33758_/Q _36062_/Q _18618_/X _18619_/X VGND VGND VPWR
+ VPWR _18650_/X sky130_fd_sc_hd__mux4_1
XFILLER_114_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27848_ _27652_/X _34265_/Q _27860_/S VGND VGND VPWR VPWR _27849_/A sky130_fd_sc_hd__mux2_1
XTAP_5175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17601_ _32897_/Q _32833_/Q _32769_/Q _32705_/Q _17346_/X _17347_/X VGND VGND VPWR
+ VPWR _17601_/X sky130_fd_sc_hd__mux4_1
XTAP_4463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18581_ _18447_/X _18579_/X _18580_/X _18450_/X VGND VGND VPWR VPWR _18581_/X sky130_fd_sc_hd__a22o_1
XTAP_4474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27779_ input39/X VGND VGND VPWR VPWR _27779_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_149_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29518_ input58/X VGND VGND VPWR VPWR _29518_/X sky130_fd_sc_hd__buf_2
X_17532_ _32127_/Q _32319_/Q _32383_/Q _35903_/Q _17280_/X _17421_/X VGND VGND VPWR
+ VPWR _17532_/X sky130_fd_sc_hd__mux4_1
XTAP_3773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30790_ _35628_/Q input15/X _30804_/S VGND VGND VPWR VPWR _30791_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29449_ _29449_/A VGND VGND VPWR VPWR _35004_/D sky130_fd_sc_hd__clkbuf_1
X_17463_ _17351_/X _17461_/X _17462_/X _17354_/X VGND VGND VPWR VPWR _17463_/X sky130_fd_sc_hd__a22o_1
XFILLER_220_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19202_ _20261_/A VGND VGND VPWR VPWR _19202_/X sky130_fd_sc_hd__buf_4
XFILLER_60_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16414_ _16091_/X _16412_/X _16413_/X _16101_/X VGND VGND VPWR VPWR _16414_/X sky130_fd_sc_hd__a22o_1
XFILLER_149_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32460_ _33393_/CLK _32460_/D VGND VGND VPWR VPWR _32460_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17394_ _17356_/X _17392_/X _17393_/X _17359_/X VGND VGND VPWR VPWR _17394_/X sky130_fd_sc_hd__a22o_1
XFILLER_164_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31411_ _31411_/A VGND VGND VPWR VPWR _35922_/D sky130_fd_sc_hd__clkbuf_1
X_19133_ _35435_/Q _35371_/Q _35307_/Q _35243_/Q _18848_/X _18849_/X VGND VGND VPWR
+ VPWR _19133_/X sky130_fd_sc_hd__mux4_1
X_16345_ _16345_/A VGND VGND VPWR VPWR _31965_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32391_ _35976_/CLK _32391_/D VGND VGND VPWR VPWR _32391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34130_ _34897_/CLK _34130_/D VGND VGND VPWR VPWR _34130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19064_ _18747_/X _19062_/X _19063_/X _18750_/X VGND VGND VPWR VPWR _19064_/X sky130_fd_sc_hd__a22o_1
X_31342_ _31342_/A VGND VGND VPWR VPWR _35889_/D sky130_fd_sc_hd__clkbuf_1
X_16276_ _33628_/Q _33564_/Q _33500_/Q _33436_/Q _16141_/X _16142_/X VGND VGND VPWR
+ VPWR _16276_/X sky130_fd_sc_hd__mux4_1
XFILLER_201_1051 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18015_ _18011_/X _18014_/X _17838_/X VGND VGND VPWR VPWR _18037_/A sky130_fd_sc_hd__o21ba_1
XFILLER_172_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34061_ _34193_/CLK _34061_/D VGND VGND VPWR VPWR _34061_/Q sky130_fd_sc_hd__dfxtp_1
X_31273_ _27825_/X _35857_/Q _31273_/S VGND VGND VPWR VPWR _31274_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33012_ _36020_/CLK _33012_/D VGND VGND VPWR VPWR _33012_/Q sky130_fd_sc_hd__dfxtp_1
X_30224_ _30335_/S VGND VGND VPWR VPWR _30243_/S sky130_fd_sc_hd__buf_4
XFILLER_172_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_908 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19966_ _32131_/Q _32323_/Q _32387_/Q _35907_/Q _19933_/X _19721_/X VGND VGND VPWR
+ VPWR _19966_/X sky130_fd_sc_hd__mux4_1
X_30155_ _35327_/Q _29457_/X _30171_/S VGND VGND VPWR VPWR _30156_/A sky130_fd_sc_hd__mux2_1
XFILLER_234_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18917_ _33061_/Q _32037_/Q _35813_/Q _35749_/Q _18672_/X _18673_/X VGND VGND VPWR
+ VPWR _18917_/X sky130_fd_sc_hd__mux4_1
X_34963_ _34963_/CLK _34963_/D VGND VGND VPWR VPWR _34963_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19897_ _32641_/Q _32577_/Q _32513_/Q _35969_/Q _19576_/X _19713_/X VGND VGND VPWR
+ VPWR _19897_/X sky130_fd_sc_hd__mux4_1
X_30086_ _30086_/A VGND VGND VPWR VPWR _35294_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_790 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33914_ _33914_/CLK _33914_/D VGND VGND VPWR VPWR _33914_/Q sky130_fd_sc_hd__dfxtp_1
X_18848_ _20260_/A VGND VGND VPWR VPWR _18848_/X sky130_fd_sc_hd__buf_4
X_34894_ _34961_/CLK _34894_/D VGND VGND VPWR VPWR _34894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33845_ _34100_/CLK _33845_/D VGND VGND VPWR VPWR _33845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18779_ _18592_/X _18777_/X _18778_/X _18595_/X VGND VGND VPWR VPWR _18779_/X sky130_fd_sc_hd__a22o_1
X_20810_ _33626_/Q _33562_/Q _33498_/Q _33434_/Q _20741_/X _20742_/X VGND VGND VPWR
+ VPWR _20810_/X sky130_fd_sc_hd__mux4_1
XFILLER_36_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33776_ _36080_/CLK _33776_/D VGND VGND VPWR VPWR _33776_/Q sky130_fd_sc_hd__dfxtp_1
X_21790_ _34677_/Q _34613_/Q _34549_/Q _34485_/Q _21539_/X _21540_/X VGND VGND VPWR
+ VPWR _21790_/X sky130_fd_sc_hd__mux4_1
X_30988_ _35722_/Q input48/X _31002_/S VGND VGND VPWR VPWR _30989_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32727_ _35863_/CLK _32727_/D VGND VGND VPWR VPWR _32727_/Q sky130_fd_sc_hd__dfxtp_1
X_20741_ _22506_/A VGND VGND VPWR VPWR _20741_/X sky130_fd_sc_hd__buf_6
X_35515_ _35709_/CLK _35515_/D VGND VGND VPWR VPWR _35515_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23460_ input47/X VGND VGND VPWR VPWR _23460_/X sky130_fd_sc_hd__buf_6
X_35446_ _35446_/CLK _35446_/D VGND VGND VPWR VPWR _35446_/Q sky130_fd_sc_hd__dfxtp_1
X_20672_ _22469_/A VGND VGND VPWR VPWR _20672_/X sky130_fd_sc_hd__buf_4
X_32658_ _35986_/CLK _32658_/D VGND VGND VPWR VPWR _32658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22411_ _32903_/Q _32839_/Q _32775_/Q _32711_/Q _22299_/X _22300_/X VGND VGND VPWR
+ VPWR _22411_/X sky130_fd_sc_hd__mux4_1
XFILLER_195_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31609_ _27723_/X _36016_/Q _31615_/S VGND VGND VPWR VPWR _31610_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35377_ _35377_/CLK _35377_/D VGND VGND VPWR VPWR _35377_/Q sky130_fd_sc_hd__dfxtp_1
X_23391_ _32209_/Q _23381_/X _23424_/S VGND VGND VPWR VPWR _23392_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32589_ _32655_/CLK _32589_/D VGND VGND VPWR VPWR _32589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25130_ _24994_/X _33045_/Q _25130_/S VGND VGND VPWR VPWR _25131_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34328_ _35609_/CLK _34328_/D VGND VGND VPWR VPWR _34328_/Q sky130_fd_sc_hd__dfxtp_1
X_22342_ _35717_/Q _32227_/Q _35589_/Q _35525_/Q _22270_/X _22271_/X VGND VGND VPWR
+ VPWR _22342_/X sky130_fd_sc_hd__mux4_1
XFILLER_148_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_1209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25061_ _25130_/S VGND VGND VPWR VPWR _25080_/S sky130_fd_sc_hd__buf_4
X_34259_ _34963_/CLK _34259_/D VGND VGND VPWR VPWR _34259_/Q sky130_fd_sc_hd__dfxtp_1
X_22273_ _35651_/Q _35011_/Q _34371_/Q _33731_/Q _22097_/X _22098_/X VGND VGND VPWR
+ VPWR _22273_/X sky130_fd_sc_hd__mux4_1
X_24012_ _24012_/A VGND VGND VPWR VPWR _32548_/D sky130_fd_sc_hd__clkbuf_1
X_21224_ _34917_/Q _34853_/Q _34789_/Q _34725_/Q _21054_/X _21055_/X VGND VGND VPWR
+ VPWR _21224_/X sky130_fd_sc_hd__mux4_1
XFILLER_219_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28820_ _28820_/A VGND VGND VPWR VPWR _34724_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21155_ _35171_/Q _35107_/Q _35043_/Q _32163_/Q _20904_/X _20905_/X VGND VGND VPWR
+ VPWR _21155_/X sky130_fd_sc_hd__mux4_1
XFILLER_144_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20106_ _20102_/X _20105_/X _19785_/X VGND VGND VPWR VPWR _20128_/A sky130_fd_sc_hd__o21ba_2
XFILLER_132_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28751_ _34693_/Q _27180_/X _28755_/S VGND VGND VPWR VPWR _28752_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25963_ _24821_/X _33437_/Q _25967_/S VGND VGND VPWR VPWR _25964_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21086_ _21047_/X _21084_/X _21085_/X _21050_/X VGND VGND VPWR VPWR _21086_/X sky130_fd_sc_hd__a22o_1
XFILLER_8_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27702_ _27701_/X _34217_/Q _27702_/S VGND VGND VPWR VPWR _27703_/A sky130_fd_sc_hd__mux2_1
X_20037_ _19712_/X _20035_/X _20036_/X _19718_/X VGND VGND VPWR VPWR _20037_/X sky130_fd_sc_hd__a22o_1
XFILLER_8_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24914_ input31/X VGND VGND VPWR VPWR _24914_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_247_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28682_ _34660_/Q _27078_/X _28692_/S VGND VGND VPWR VPWR _28683_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25894_ _25894_/A VGND VGND VPWR VPWR _33404_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27633_ _34195_/Q _27223_/X _27637_/S VGND VGND VPWR VPWR _27634_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24845_ _24845_/A VGND VGND VPWR VPWR _32932_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27564_ _34162_/Q _27121_/X _27566_/S VGND VGND VPWR VPWR _27565_/A sky130_fd_sc_hd__mux2_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24776_ _23055_/X _32908_/Q _24786_/S VGND VGND VPWR VPWR _24777_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21988_ _21984_/X _21987_/X _21740_/X _21741_/X VGND VGND VPWR VPWR _22003_/B sky130_fd_sc_hd__o211a_1
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29303_ _29303_/A VGND VGND VPWR VPWR _34953_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_226_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26515_ _26515_/A VGND VGND VPWR VPWR _33697_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20939_ _20678_/X _20937_/X _20938_/X _20688_/X VGND VGND VPWR VPWR _20939_/X sky130_fd_sc_hd__a22o_1
X_23727_ _22915_/X _32351_/Q _23727_/S VGND VGND VPWR VPWR _23728_/A sky130_fd_sc_hd__mux2_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27495_ _27495_/A VGND VGND VPWR VPWR _34129_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29234_ _34921_/Q _27093_/X _29234_/S VGND VGND VPWR VPWR _29235_/A sky130_fd_sc_hd__mux2_1
X_26446_ _26446_/A VGND VGND VPWR VPWR _33665_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23658_ _23658_/A VGND VGND VPWR VPWR _32319_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22609_ _33677_/Q _33613_/Q _33549_/Q _33485_/Q _22506_/X _22507_/X VGND VGND VPWR
+ VPWR _22609_/X sky130_fd_sc_hd__mux4_1
X_29165_ _34888_/Q _27189_/X _29183_/S VGND VGND VPWR VPWR _29166_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23589_ _22915_/X _32287_/Q _23589_/S VGND VGND VPWR VPWR _23590_/A sky130_fd_sc_hd__mux2_1
X_26377_ _26377_/A VGND VGND VPWR VPWR _33632_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28116_ _27649_/X _34392_/Q _28130_/S VGND VGND VPWR VPWR _28117_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16130_ _16126_/X _16129_/X _16075_/X VGND VGND VPWR VPWR _16138_/C sky130_fd_sc_hd__o21ba_1
XFILLER_167_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_1336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25328_ _33137_/Q _23364_/X _25332_/S VGND VGND VPWR VPWR _25329_/A sky130_fd_sc_hd__mux2_1
X_29096_ _29096_/A VGND VGND VPWR VPWR _34855_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16061_ _16061_/A VGND VGND VPWR VPWR _17850_/A sky130_fd_sc_hd__buf_12
X_28047_ _28047_/A VGND VGND VPWR VPWR _34359_/D sky130_fd_sc_hd__clkbuf_1
X_25259_ _33105_/Q _23484_/X _25259_/S VGND VGND VPWR VPWR _25260_/A sky130_fd_sc_hd__mux2_1
XFILLER_237_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19820_ _19820_/A _19820_/B _19820_/C _19820_/D VGND VGND VPWR VPWR _19821_/A sky130_fd_sc_hd__or4_4
XFILLER_97_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29998_ _29998_/A VGND VGND VPWR VPWR _35252_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19751_ _33917_/Q _33853_/Q _33789_/Q _36093_/Q _19677_/X _19678_/X VGND VGND VPWR
+ VPWR _19751_/X sky130_fd_sc_hd__mux4_1
X_28949_ _28949_/A VGND VGND VPWR VPWR _34785_/D sky130_fd_sc_hd__clkbuf_1
X_16963_ _16959_/X _16962_/X _16787_/X _16788_/X VGND VGND VPWR VPWR _16980_/B sky130_fd_sc_hd__o211a_1
XFILLER_238_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18702_ _35679_/Q _32185_/Q _35551_/Q _35487_/Q _18558_/X _18559_/X VGND VGND VPWR
+ VPWR _18702_/X sky130_fd_sc_hd__mux4_1
XFILLER_49_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_6_28__f_CLK clkbuf_5_14_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_28__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_42_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31960_ _34148_/CLK _31960_/D VGND VGND VPWR VPWR _31960_/Q sky130_fd_sc_hd__dfxtp_1
X_19682_ _32635_/Q _32571_/Q _32507_/Q _35963_/Q _19576_/X _19360_/X VGND VGND VPWR
+ VPWR _19682_/X sky130_fd_sc_hd__mux4_1
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16894_ _32109_/Q _32301_/Q _32365_/Q _35885_/Q _16574_/X _16715_/X VGND VGND VPWR
+ VPWR _16894_/X sky130_fd_sc_hd__mux4_1
XFILLER_237_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18633_ _35421_/Q _35357_/Q _35293_/Q _35229_/Q _18495_/X _18496_/X VGND VGND VPWR
+ VPWR _18633_/X sky130_fd_sc_hd__mux4_1
X_30911_ _30911_/A VGND VGND VPWR VPWR _35685_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31891_ _31891_/A VGND VGND VPWR VPWR _36149_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33630_ _36191_/CLK _33630_/D VGND VGND VPWR VPWR _33630_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30842_ _35653_/Q input42/X _30846_/S VGND VGND VPWR VPWR _30843_/A sky130_fd_sc_hd__mux2_1
X_18564_ _33051_/Q _32027_/Q _35803_/Q _35739_/Q _18367_/X _18369_/X VGND VGND VPWR
+ VPWR _18564_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17515_ _34942_/Q _34878_/Q _34814_/Q _34750_/Q _17513_/X _17514_/X VGND VGND VPWR
+ VPWR _17515_/X sky130_fd_sc_hd__mux4_1
XTAP_3592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33561_ _34009_/CLK _33561_/D VGND VGND VPWR VPWR _33561_/Q sky130_fd_sc_hd__dfxtp_1
X_18495_ _20150_/A VGND VGND VPWR VPWR _18495_/X sky130_fd_sc_hd__buf_6
X_30773_ _35620_/Q input6/X _30783_/S VGND VGND VPWR VPWR _30774_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35300_ _35817_/CLK _35300_/D VGND VGND VPWR VPWR _35300_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32512_ _35969_/CLK _32512_/D VGND VGND VPWR VPWR _32512_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17446_ _17960_/A VGND VGND VPWR VPWR _17446_/X sky130_fd_sc_hd__buf_8
X_33492_ _33685_/CLK _33492_/D VGND VGND VPWR VPWR _33492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35231_ _35743_/CLK _35231_/D VGND VGND VPWR VPWR _35231_/Q sky130_fd_sc_hd__dfxtp_1
X_32443_ _33895_/CLK _32443_/D VGND VGND VPWR VPWR _32443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17377_ _17850_/A VGND VGND VPWR VPWR _17377_/X sky130_fd_sc_hd__buf_8
XFILLER_207_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_1184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19116_ _33643_/Q _33579_/Q _33515_/Q _33451_/Q _18794_/X _18795_/X VGND VGND VPWR
+ VPWR _19116_/X sky130_fd_sc_hd__mux4_1
X_35162_ _35162_/CLK _35162_/D VGND VGND VPWR VPWR _35162_/Q sky130_fd_sc_hd__dfxtp_1
X_16328_ _16030_/X _16326_/X _16327_/X _16041_/X VGND VGND VPWR VPWR _16328_/X sky130_fd_sc_hd__a22o_1
XFILLER_229_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32374_ _32887_/CLK _32374_/D VGND VGND VPWR VPWR _32374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34113_ _34177_/CLK _34113_/D VGND VGND VPWR VPWR _34113_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19047_ _19043_/X _19046_/X _18726_/X VGND VGND VPWR VPWR _19069_/A sky130_fd_sc_hd__o21ba_1
XFILLER_51_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31325_ _31325_/A VGND VGND VPWR VPWR _35881_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35093_ _35865_/CLK _35093_/D VGND VGND VPWR VPWR _35093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16259_ _17800_/A VGND VGND VPWR VPWR _16259_/X sky130_fd_sc_hd__buf_4
XFILLER_145_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput202 _36235_/Q VGND VGND VPWR VPWR D2[53] sky130_fd_sc_hd__buf_2
Xoutput213 _36245_/Q VGND VGND VPWR VPWR D2[63] sky130_fd_sc_hd__buf_2
XFILLER_245_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34044_ _34172_/CLK _34044_/D VGND VGND VPWR VPWR _34044_/Q sky130_fd_sc_hd__dfxtp_1
X_31256_ _31256_/A VGND VGND VPWR VPWR _35848_/D sky130_fd_sc_hd__clkbuf_1
Xoutput224 _32421_/Q VGND VGND VPWR VPWR D3[15] sky130_fd_sc_hd__buf_2
XFILLER_173_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput235 _32431_/Q VGND VGND VPWR VPWR D3[25] sky130_fd_sc_hd__buf_2
XFILLER_245_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput246 _32441_/Q VGND VGND VPWR VPWR D3[35] sky130_fd_sc_hd__buf_2
XFILLER_47_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30207_ _30207_/A VGND VGND VPWR VPWR _35351_/D sky130_fd_sc_hd__clkbuf_1
Xoutput257 _32451_/Q VGND VGND VPWR VPWR D3[45] sky130_fd_sc_hd__buf_2
XFILLER_47_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput268 _32461_/Q VGND VGND VPWR VPWR D3[55] sky130_fd_sc_hd__buf_2
XFILLER_173_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput279 _32413_/Q VGND VGND VPWR VPWR D3[7] sky130_fd_sc_hd__buf_2
X_31187_ _27698_/X _35816_/Q _31189_/S VGND VGND VPWR VPWR _31188_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30138_ _35319_/Q _29432_/X _30150_/S VGND VGND VPWR VPWR _30139_/A sky130_fd_sc_hd__mux2_1
X_19949_ _19806_/X _19947_/X _19948_/X _19809_/X VGND VGND VPWR VPWR _19949_/X sky130_fd_sc_hd__a22o_1
XFILLER_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35995_ _35995_/CLK _35995_/D VGND VGND VPWR VPWR _35995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22960_ _22959_/X _32045_/Q _22978_/S VGND VGND VPWR VPWR _22961_/A sky130_fd_sc_hd__mux2_1
X_30069_ _35286_/Q _29328_/X _30087_/S VGND VGND VPWR VPWR _30070_/A sky130_fd_sc_hd__mux2_1
X_34946_ _36163_/CLK _34946_/D VGND VGND VPWR VPWR _34946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21911_ _33145_/Q _36025_/Q _33017_/Q _32953_/Q _21662_/X _21663_/X VGND VGND VPWR
+ VPWR _21911_/X sky130_fd_sc_hd__mux4_1
XFILLER_228_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22891_ input12/X VGND VGND VPWR VPWR _22891_/X sky130_fd_sc_hd__buf_2
XFILLER_28_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34877_ _34877_/CLK _34877_/D VGND VGND VPWR VPWR _34877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24630_ _23039_/X _32839_/Q _24630_/S VGND VGND VPWR VPWR _24631_/A sky130_fd_sc_hd__mux2_1
X_21842_ _21806_/X _21840_/X _21841_/X _21809_/X VGND VGND VPWR VPWR _21842_/X sky130_fd_sc_hd__a22o_1
XFILLER_243_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33828_ _33828_/CLK _33828_/D VGND VGND VPWR VPWR _33828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24561_ _22937_/X _32806_/Q _24567_/S VGND VGND VPWR VPWR _24562_/A sky130_fd_sc_hd__mux2_1
X_33759_ _35551_/CLK _33759_/D VGND VGND VPWR VPWR _33759_/Q sky130_fd_sc_hd__dfxtp_1
X_21773_ _33909_/Q _33845_/Q _33781_/Q _36085_/Q _21624_/X _21625_/X VGND VGND VPWR
+ VPWR _21773_/X sky130_fd_sc_hd__mux4_1
XFILLER_208_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26300_ _24920_/X _33597_/Q _26300_/S VGND VGND VPWR VPWR _26301_/A sky130_fd_sc_hd__mux2_1
X_20724_ _35671_/Q _32177_/Q _35543_/Q _35479_/Q _20649_/X _20650_/X VGND VGND VPWR
+ VPWR _20724_/X sky130_fd_sc_hd__mux4_1
XFILLER_184_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23512_ _23512_/A VGND VGND VPWR VPWR _32251_/D sky130_fd_sc_hd__clkbuf_1
X_24492_ _24492_/A VGND VGND VPWR VPWR _32773_/D sky130_fd_sc_hd__clkbuf_1
X_27280_ _34027_/Q _27100_/X _27296_/S VGND VGND VPWR VPWR _27281_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23443_ _23443_/A VGND VGND VPWR VPWR _32226_/D sky130_fd_sc_hd__clkbuf_1
X_26231_ _24818_/X _33564_/Q _26237_/S VGND VGND VPWR VPWR _26232_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20655_ _22599_/A VGND VGND VPWR VPWR _20655_/X sky130_fd_sc_hd__buf_4
XFILLER_23_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35429_ _35817_/CLK _35429_/D VGND VGND VPWR VPWR _35429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26162_ _26162_/A VGND VGND VPWR VPWR _33531_/D sky130_fd_sc_hd__clkbuf_1
X_23374_ _23374_/A VGND VGND VPWR VPWR _32202_/D sky130_fd_sc_hd__clkbuf_1
X_20586_ _20663_/A VGND VGND VPWR VPWR _22507_/A sky130_fd_sc_hd__buf_12
XFILLER_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22325_ _22325_/A VGND VGND VPWR VPWR _36228_/D sky130_fd_sc_hd__clkbuf_1
X_25113_ _25113_/A VGND VGND VPWR VPWR _33036_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26093_ _26093_/A VGND VGND VPWR VPWR _33498_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29921_ _29921_/A VGND VGND VPWR VPWR _35216_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25044_ _25044_/A VGND VGND VPWR VPWR _33003_/D sky130_fd_sc_hd__clkbuf_1
X_22256_ _33667_/Q _33603_/Q _33539_/Q _33475_/Q _22153_/X _22154_/X VGND VGND VPWR
+ VPWR _22256_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21207_ _32101_/Q _32293_/Q _32357_/Q _35877_/Q _21174_/X _20962_/X VGND VGND VPWR
+ VPWR _21207_/X sky130_fd_sc_hd__mux4_1
X_29852_ _29852_/A VGND VGND VPWR VPWR _35183_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_160_CLK clkbuf_6_31__f_CLK/X VGND VGND VPWR VPWR _36177_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_191_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22187_ _22181_/X _22186_/X _22118_/X VGND VGND VPWR VPWR _22188_/D sky130_fd_sc_hd__o21ba_1
XFILLER_2_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28803_ _28803_/A VGND VGND VPWR VPWR _34716_/D sky130_fd_sc_hd__clkbuf_1
X_21138_ _32611_/Q _32547_/Q _32483_/Q _35939_/Q _20817_/X _20954_/X VGND VGND VPWR
+ VPWR _21138_/X sky130_fd_sc_hd__mux4_1
X_29783_ _35151_/Q _29506_/X _29787_/S VGND VGND VPWR VPWR _29784_/A sky130_fd_sc_hd__mux2_1
X_26995_ _26995_/A VGND VGND VPWR VPWR _33923_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28734_ _34685_/Q _27155_/X _28734_/S VGND VGND VPWR VPWR _28735_/A sky130_fd_sc_hd__mux2_1
X_25946_ _25946_/A VGND VGND VPWR VPWR _33429_/D sky130_fd_sc_hd__clkbuf_1
X_21069_ _21065_/X _21068_/X _21026_/X VGND VGND VPWR VPWR _21091_/A sky130_fd_sc_hd__o21ba_1
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28665_ _34652_/Q _27053_/X _28671_/S VGND VGND VPWR VPWR _28666_/A sky130_fd_sc_hd__mux2_1
XFILLER_207_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25877_ _24892_/X _33396_/Q _25895_/S VGND VGND VPWR VPWR _25878_/A sky130_fd_sc_hd__mux2_1
XFILLER_206_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_246_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27616_ _27616_/A VGND VGND VPWR VPWR _34186_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_185_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24828_ _24827_/X _32927_/Q _24828_/S VGND VGND VPWR VPWR _24829_/A sky130_fd_sc_hd__mux2_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28596_ _27760_/X _34620_/Q _28598_/S VGND VGND VPWR VPWR _28597_/A sky130_fd_sc_hd__mux2_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_12_0_CLK clkbuf_5_9_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_12_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27547_ _27637_/S VGND VGND VPWR VPWR _27566_/S sky130_fd_sc_hd__buf_4
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24759_ _23030_/X _32900_/Q _24765_/S VGND VGND VPWR VPWR _24760_/A sky130_fd_sc_hd__mux2_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17300_ _17296_/X _17299_/X _17165_/X VGND VGND VPWR VPWR _17301_/D sky130_fd_sc_hd__o21ba_1
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18280_ _20065_/A VGND VGND VPWR VPWR _20159_/A sky130_fd_sc_hd__buf_12
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27478_ _34121_/Q _27193_/X _27494_/S VGND VGND VPWR VPWR _27479_/A sky130_fd_sc_hd__mux2_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29217_ _29217_/A VGND VGND VPWR VPWR _34912_/D sky130_fd_sc_hd__clkbuf_1
X_17231_ _34422_/Q _36150_/Q _34294_/Q _34230_/Q _17229_/X _17230_/X VGND VGND VPWR
+ VPWR _17231_/X sky130_fd_sc_hd__mux4_1
X_26429_ _26429_/A VGND VGND VPWR VPWR _33657_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_204_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_27_0_CLK clkbuf_2_3_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_27_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_11_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29148_ _34880_/Q _27165_/X _29162_/S VGND VGND VPWR VPWR _29149_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17162_ _34932_/Q _34868_/Q _34804_/Q _34740_/Q _17160_/X _17161_/X VGND VGND VPWR
+ VPWR _17162_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16113_ _17851_/A VGND VGND VPWR VPWR _16113_/X sky130_fd_sc_hd__buf_4
X_29079_ _29079_/A VGND VGND VPWR VPWR _34847_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17093_ _17960_/A VGND VGND VPWR VPWR _17093_/X sky130_fd_sc_hd__buf_4
XFILLER_10_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31110_ _35780_/Q input41/X _31116_/S VGND VGND VPWR VPWR _31111_/A sky130_fd_sc_hd__mux2_1
X_16044_ _17846_/A VGND VGND VPWR VPWR _16044_/X sky130_fd_sc_hd__buf_4
X_32090_ _35995_/CLK _32090_/D VGND VGND VPWR VPWR _32090_/Q sky130_fd_sc_hd__dfxtp_1
X_31041_ _35747_/Q input5/X _31053_/S VGND VGND VPWR VPWR _31042_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_151_CLK clkbuf_6_29__f_CLK/X VGND VGND VPWR VPWR _34964_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_9_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19803_ _19656_/X _19801_/X _19802_/X _19659_/X VGND VGND VPWR VPWR _19803_/X sky130_fd_sc_hd__a22o_1
XFILLER_215_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17995_ _33100_/Q _32076_/Q _35852_/Q _35788_/Q _17784_/X _17785_/X VGND VGND VPWR
+ VPWR _17995_/X sky130_fd_sc_hd__mux4_1
XFILLER_111_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_950 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34800_ _35439_/CLK _34800_/D VGND VGND VPWR VPWR _34800_/Q sky130_fd_sc_hd__dfxtp_1
X_16946_ _16805_/X _16944_/X _16945_/X _16810_/X VGND VGND VPWR VPWR _16946_/X sky130_fd_sc_hd__a22o_1
X_19734_ _19656_/X _19730_/X _19733_/X _19659_/X VGND VGND VPWR VPWR _19734_/X sky130_fd_sc_hd__a22o_1
X_35780_ _36038_/CLK _35780_/D VGND VGND VPWR VPWR _35780_/Q sky130_fd_sc_hd__dfxtp_1
X_32992_ _36129_/CLK _32992_/D VGND VGND VPWR VPWR _32992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31943_ _31943_/A VGND VGND VPWR VPWR _36174_/D sky130_fd_sc_hd__clkbuf_1
X_34731_ _34924_/CLK _34731_/D VGND VGND VPWR VPWR _34731_/Q sky130_fd_sc_hd__dfxtp_1
X_19665_ _35194_/Q _35130_/Q _35066_/Q _32250_/Q _19663_/X _19664_/X VGND VGND VPWR
+ VPWR _19665_/X sky130_fd_sc_hd__mux4_1
XFILLER_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16877_ _16877_/A VGND VGND VPWR VPWR _16877_/X sky130_fd_sc_hd__buf_4
X_18616_ _18440_/X _18614_/X _18615_/X _18445_/X VGND VGND VPWR VPWR _18616_/X sky130_fd_sc_hd__a22o_1
XTAP_4090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34662_ _35618_/CLK _34662_/D VGND VGND VPWR VPWR _34662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19596_ _19453_/X _19594_/X _19595_/X _19456_/X VGND VGND VPWR VPWR _19596_/X sky130_fd_sc_hd__a22o_1
X_31874_ _31874_/A VGND VGND VPWR VPWR _36141_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_225_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33613_ _34193_/CLK _33613_/D VGND VGND VPWR VPWR _33613_/Q sky130_fd_sc_hd__dfxtp_1
X_18547_ _33371_/Q _33307_/Q _33243_/Q _33179_/Q _18302_/X _18303_/X VGND VGND VPWR
+ VPWR _18547_/X sky130_fd_sc_hd__mux4_1
X_30825_ _35645_/Q input33/X _30825_/S VGND VGND VPWR VPWR _30826_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34593_ _34593_/CLK _34593_/D VGND VGND VPWR VPWR _34593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33544_ _33673_/CLK _33544_/D VGND VGND VPWR VPWR _33544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18478_ _33625_/Q _33561_/Q _33497_/Q _33433_/Q _18441_/X _18442_/X VGND VGND VPWR
+ VPWR _18478_/X sky130_fd_sc_hd__mux4_1
X_30756_ _35612_/Q input61/X _30762_/S VGND VGND VPWR VPWR _30757_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17429_ _17351_/X _17427_/X _17428_/X _17354_/X VGND VGND VPWR VPWR _17429_/X sky130_fd_sc_hd__a22o_1
X_33475_ _34180_/CLK _33475_/D VGND VGND VPWR VPWR _33475_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30687_ _30687_/A VGND VGND VPWR VPWR _35579_/D sky130_fd_sc_hd__clkbuf_1
X_35214_ _35731_/CLK _35214_/D VGND VGND VPWR VPWR _35214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20440_ _32913_/Q _32849_/Q _32785_/Q _32721_/Q _18284_/X _18287_/X VGND VGND VPWR
+ VPWR _20440_/X sky130_fd_sc_hd__mux4_1
XFILLER_14_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32426_ _33895_/CLK _32426_/D VGND VGND VPWR VPWR _32426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36194_ _36209_/CLK _36194_/D VGND VGND VPWR VPWR _36194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35145_ _35210_/CLK _35145_/D VGND VGND VPWR VPWR _35145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20371_ _20205_/X _20369_/X _20370_/X _20210_/X VGND VGND VPWR VPWR _20371_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32357_ _35945_/CLK _32357_/D VGND VGND VPWR VPWR _32357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_390_CLK clkbuf_6_40__f_CLK/X VGND VGND VPWR VPWR _36087_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_162_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22110_ _22106_/X _22107_/X _22108_/X _22109_/X VGND VGND VPWR VPWR _22110_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31308_ _27677_/X _35873_/Q _31324_/S VGND VGND VPWR VPWR _31309_/A sky130_fd_sc_hd__mux2_1
X_35076_ _35717_/CLK _35076_/D VGND VGND VPWR VPWR _35076_/Q sky130_fd_sc_hd__dfxtp_1
X_23090_ _31418_/A _28110_/A VGND VGND VPWR VPWR _23223_/S sky130_fd_sc_hd__nand2_8
X_32288_ _35875_/CLK _32288_/D VGND VGND VPWR VPWR _32288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34027_ _35627_/CLK _34027_/D VGND VGND VPWR VPWR _34027_/Q sky130_fd_sc_hd__dfxtp_1
X_22041_ _21758_/X _22039_/X _22040_/X _21763_/X VGND VGND VPWR VPWR _22041_/X sky130_fd_sc_hd__a22o_1
XTAP_6409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_142_CLK clkbuf_6_28__f_CLK/X VGND VGND VPWR VPWR _35863_/CLK sky130_fd_sc_hd__clkbuf_16
X_31239_ _31239_/A VGND VGND VPWR VPWR _35840_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25800_ _24979_/X _33360_/Q _25802_/S VGND VGND VPWR VPWR _25801_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26780_ _26780_/A VGND VGND VPWR VPWR _33821_/D sky130_fd_sc_hd__clkbuf_1
X_23992_ _22903_/X _32539_/Q _24000_/S VGND VGND VPWR VPWR _23993_/A sky130_fd_sc_hd__mux2_1
X_35978_ _35978_/CLK _35978_/D VGND VGND VPWR VPWR _35978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_217_904 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25731_ _24877_/X _33327_/Q _25739_/S VGND VGND VPWR VPWR _25732_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_6_11__f_CLK clkbuf_5_5_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_11__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_25_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34929_ _35633_/CLK _34929_/D VGND VGND VPWR VPWR _34929_/Q sky130_fd_sc_hd__dfxtp_1
X_22943_ input10/X VGND VGND VPWR VPWR _22943_/X sky130_fd_sc_hd__buf_2
XFILLER_229_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28450_ _28450_/A VGND VGND VPWR VPWR _34550_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25662_ _25662_/A VGND VGND VPWR VPWR _33294_/D sky130_fd_sc_hd__clkbuf_1
X_22874_ _34965_/Q _34901_/Q _34837_/Q _34773_/Q _20683_/X _20685_/X VGND VGND VPWR
+ VPWR _22874_/X sky130_fd_sc_hd__mux4_1
XFILLER_55_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27401_ _27401_/A VGND VGND VPWR VPWR _34084_/D sky130_fd_sc_hd__clkbuf_1
X_24613_ _24613_/A VGND VGND VPWR VPWR _32830_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_227_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28381_ _28513_/S VGND VGND VPWR VPWR _28400_/S sky130_fd_sc_hd__clkbuf_8
X_21825_ _21821_/X _21824_/X _21751_/X VGND VGND VPWR VPWR _21835_/C sky130_fd_sc_hd__o21ba_1
X_25593_ _25593_/A VGND VGND VPWR VPWR _33261_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_1032 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27332_ _34052_/Q _27177_/X _27338_/S VGND VGND VPWR VPWR _27333_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24544_ _22912_/X _32798_/Q _24546_/S VGND VGND VPWR VPWR _24545_/A sky130_fd_sc_hd__mux2_1
X_21756_ _21756_/A VGND VGND VPWR VPWR _21756_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_169_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20707_ _20707_/A VGND VGND VPWR VPWR _36182_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_169_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27263_ _34019_/Q _27075_/X _27275_/S VGND VGND VPWR VPWR _27264_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24475_ _24475_/A VGND VGND VPWR VPWR _32765_/D sky130_fd_sc_hd__clkbuf_1
X_21687_ _34930_/Q _34866_/Q _34802_/Q _34738_/Q _21407_/X _21408_/X VGND VGND VPWR
+ VPWR _21687_/X sky130_fd_sc_hd__mux4_1
XFILLER_11_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29002_ _34811_/Q _27149_/X _29006_/S VGND VGND VPWR VPWR _29003_/A sky130_fd_sc_hd__mux2_1
X_26214_ _26214_/A VGND VGND VPWR VPWR _33556_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20638_ _20663_/A VGND VGND VPWR VPWR _22434_/A sky130_fd_sc_hd__buf_12
XFILLER_149_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23426_ input36/X VGND VGND VPWR VPWR _23426_/X sky130_fd_sc_hd__buf_4
X_27194_ _33993_/Q _27193_/X _27218_/S VGND VGND VPWR VPWR _27195_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23357_ _32195_/Q _23286_/X _23359_/S VGND VGND VPWR VPWR _23358_/A sky130_fd_sc_hd__mux2_1
X_26145_ _26145_/A VGND VGND VPWR VPWR _33523_/D sky130_fd_sc_hd__clkbuf_1
X_20569_ _20565_/X _20568_/X _20157_/A VGND VGND VPWR VPWR _20577_/C sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_381_CLK clkbuf_6_42__f_CLK/X VGND VGND VPWR VPWR _36093_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_165_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22308_ _22304_/X _22305_/X _22306_/X _22307_/X VGND VGND VPWR VPWR _22308_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26076_ _24988_/X _33491_/Q _26080_/S VGND VGND VPWR VPWR _26077_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23288_ _23288_/A VGND VGND VPWR VPWR _32168_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29904_ _35208_/Q _29484_/X _29922_/S VGND VGND VPWR VPWR _29905_/A sky130_fd_sc_hd__mux2_1
X_22239_ _35650_/Q _35010_/Q _34370_/Q _33730_/Q _22097_/X _22098_/X VGND VGND VPWR
+ VPWR _22239_/X sky130_fd_sc_hd__mux4_1
X_25027_ _25027_/A VGND VGND VPWR VPWR _32995_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_133_CLK clkbuf_6_23__f_CLK/X VGND VGND VPWR VPWR _34647_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_6910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29835_ _29835_/A VGND VGND VPWR VPWR _35175_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16800_ _17153_/A VGND VGND VPWR VPWR _16800_/X sky130_fd_sc_hd__clkbuf_4
XTAP_6987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29766_ _35143_/Q _29481_/X _29766_/S VGND VGND VPWR VPWR _29767_/A sky130_fd_sc_hd__mux2_1
X_17780_ _35718_/Q _32228_/Q _35590_/Q _35526_/Q _17670_/X _17671_/X VGND VGND VPWR
+ VPWR _17780_/X sky130_fd_sc_hd__mux4_1
XFILLER_121_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26978_ _26978_/A VGND VGND VPWR VPWR _33915_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16731_ _35176_/Q _35112_/Q _35048_/Q _32168_/Q _16657_/X _16658_/X VGND VGND VPWR
+ VPWR _16731_/X sky130_fd_sc_hd__mux4_1
X_28717_ _28717_/A VGND VGND VPWR VPWR _34676_/D sky130_fd_sc_hd__clkbuf_1
X_25929_ _24970_/X _33421_/Q _25937_/S VGND VGND VPWR VPWR _25930_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29697_ _35110_/Q _29379_/X _29703_/S VGND VGND VPWR VPWR _29698_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19450_ _19303_/X _19448_/X _19449_/X _19306_/X VGND VGND VPWR VPWR _19450_/X sky130_fd_sc_hd__a22o_1
X_28648_ _27837_/X _34645_/Q _28648_/S VGND VGND VPWR VPWR _28649_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16662_ _34918_/Q _34854_/Q _34790_/Q _34726_/Q _16454_/X _16455_/X VGND VGND VPWR
+ VPWR _16662_/X sky130_fd_sc_hd__mux4_1
XFILLER_235_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18401_ _19463_/A VGND VGND VPWR VPWR _18401_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_61_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19381_ _19303_/X _19377_/X _19380_/X _19306_/X VGND VGND VPWR VPWR _19381_/X sky130_fd_sc_hd__a22o_1
XFILLER_90_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_222_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16593_ _16452_/X _16591_/X _16592_/X _16457_/X VGND VGND VPWR VPWR _16593_/X sky130_fd_sc_hd__a22o_1
X_28579_ _28648_/S VGND VGND VPWR VPWR _28598_/S sky130_fd_sc_hd__buf_4
XFILLER_90_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30610_ _30610_/A VGND VGND VPWR VPWR _35542_/D sky130_fd_sc_hd__clkbuf_1
X_18332_ _20286_/A VGND VGND VPWR VPWR _18332_/X sky130_fd_sc_hd__buf_6
XFILLER_37_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31590_ _27695_/X _36007_/Q _31594_/S VGND VGND VPWR VPWR _31591_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18263_ _35733_/Q _32245_/Q _35605_/Q _35541_/Q _15993_/X _15995_/X VGND VGND VPWR
+ VPWR _18263_/X sky130_fd_sc_hd__mux4_1
X_30541_ _35510_/Q _29429_/X _30555_/S VGND VGND VPWR VPWR _30542_/A sky130_fd_sc_hd__mux2_1
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17214_ _17059_/X _17212_/X _17213_/X _17065_/X VGND VGND VPWR VPWR _17214_/X sky130_fd_sc_hd__a22o_1
X_33260_ _36076_/CLK _33260_/D VGND VGND VPWR VPWR _33260_/Q sky130_fd_sc_hd__dfxtp_1
X_18194_ _17912_/X _18192_/X _18193_/X _17915_/X VGND VGND VPWR VPWR _18194_/X sky130_fd_sc_hd__a22o_1
X_30472_ _30472_/A _30877_/A VGND VGND VPWR VPWR _30605_/S sky130_fd_sc_hd__nor2_8
XFILLER_200_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32211_ _35703_/CLK _32211_/D VGND VGND VPWR VPWR _32211_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17145_ _17999_/A VGND VGND VPWR VPWR _17145_/X sky130_fd_sc_hd__buf_4
X_33191_ _36072_/CLK _33191_/D VGND VGND VPWR VPWR _33191_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_372_CLK clkbuf_6_43__f_CLK/X VGND VGND VPWR VPWR _36154_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_200_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32142_ _35921_/CLK _32142_/D VGND VGND VPWR VPWR _32142_/Q sky130_fd_sc_hd__dfxtp_1
X_17076_ _16998_/X _17074_/X _17075_/X _17001_/X VGND VGND VPWR VPWR _17076_/X sky130_fd_sc_hd__a22o_1
XFILLER_155_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16027_ _17910_/A VGND VGND VPWR VPWR _16027_/X sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_124_CLK clkbuf_6_21__f_CLK/X VGND VGND VPWR VPWR _36242_/CLK sky130_fd_sc_hd__clkbuf_16
X_32073_ _33160_/CLK _32073_/D VGND VGND VPWR VPWR _32073_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_671 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31024_ _35739_/Q input56/X _31032_/S VGND VGND VPWR VPWR _31025_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35901_ _35962_/CLK _35901_/D VGND VGND VPWR VPWR _35901_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35832_ _35833_/CLK _35832_/D VGND VGND VPWR VPWR _35832_/Q sky130_fd_sc_hd__dfxtp_1
X_17978_ _33420_/Q _33356_/Q _33292_/Q _33228_/Q _17833_/X _17834_/X VGND VGND VPWR
+ VPWR _17978_/X sky130_fd_sc_hd__mux4_1
XFILLER_211_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16929_ _32878_/Q _32814_/Q _32750_/Q _32686_/Q _16640_/X _16641_/X VGND VGND VPWR
+ VPWR _16929_/X sky130_fd_sc_hd__mux4_1
X_19717_ _33148_/Q _36028_/Q _33020_/Q _32956_/Q _19715_/X _19716_/X VGND VGND VPWR
+ VPWR _19717_/X sky130_fd_sc_hd__mux4_1
X_32975_ _36045_/CLK _32975_/D VGND VGND VPWR VPWR _32975_/Q sky130_fd_sc_hd__dfxtp_1
X_35763_ _36147_/CLK _35763_/D VGND VGND VPWR VPWR _35763_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34714_ _36245_/CLK _34714_/D VGND VGND VPWR VPWR _34714_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31926_ _31926_/A VGND VGND VPWR VPWR _36166_/D sky130_fd_sc_hd__clkbuf_1
X_19648_ _32890_/Q _32826_/Q _32762_/Q _32698_/Q _19646_/X _19647_/X VGND VGND VPWR
+ VPWR _19648_/X sky130_fd_sc_hd__mux4_1
X_35694_ _35694_/CLK _35694_/D VGND VGND VPWR VPWR _35694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34645_ _36117_/CLK _34645_/D VGND VGND VPWR VPWR _34645_/Q sky130_fd_sc_hd__dfxtp_1
X_31857_ _31857_/A VGND VGND VPWR VPWR _36133_/D sky130_fd_sc_hd__clkbuf_1
X_19579_ _19359_/X _19577_/X _19578_/X _19365_/X VGND VGND VPWR VPWR _19579_/X sky130_fd_sc_hd__a22o_1
XFILLER_197_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_1190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21610_ _22316_/A VGND VGND VPWR VPWR _21610_/X sky130_fd_sc_hd__buf_4
X_30808_ _30808_/A VGND VGND VPWR VPWR _35636_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22590_ _22585_/X _22589_/X _22446_/X _22447_/X VGND VGND VPWR VPWR _22607_/B sky130_fd_sc_hd__o211a_2
XFILLER_55_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34576_ _36177_/CLK _34576_/D VGND VGND VPWR VPWR _34576_/Q sky130_fd_sc_hd__dfxtp_1
X_31788_ _36101_/Q input42/X _31792_/S VGND VGND VPWR VPWR _31789_/A sky130_fd_sc_hd__mux2_1
XFILLER_209_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_244_1076 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21541_ _34670_/Q _34606_/Q _34542_/Q _34478_/Q _21539_/X _21540_/X VGND VGND VPWR
+ VPWR _21541_/X sky130_fd_sc_hd__mux4_1
X_30739_ _30739_/A VGND VGND VPWR VPWR _35604_/D sky130_fd_sc_hd__clkbuf_1
X_33527_ _33850_/CLK _33527_/D VGND VGND VPWR VPWR _33527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24260_ _22891_/X _32663_/Q _24276_/S VGND VGND VPWR VPWR _24261_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33458_ _34098_/CLK _33458_/D VGND VGND VPWR VPWR _33458_/Q sky130_fd_sc_hd__dfxtp_1
X_21472_ _21468_/X _21471_/X _21398_/X VGND VGND VPWR VPWR _21482_/C sky130_fd_sc_hd__o21ba_1
XFILLER_193_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23211_ _23064_/X _32143_/Q _23215_/S VGND VGND VPWR VPWR _23212_/A sky130_fd_sc_hd__mux2_1
X_20423_ _34448_/Q _36176_/Q _34320_/Q _34256_/Q _20235_/X _20236_/X VGND VGND VPWR
+ VPWR _20423_/X sky130_fd_sc_hd__mux4_1
X_32409_ _34151_/CLK _32409_/D VGND VGND VPWR VPWR _32409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24191_ _32632_/Q _23402_/X _24201_/S VGND VGND VPWR VPWR _24192_/A sky130_fd_sc_hd__mux2_1
X_36177_ _36177_/CLK _36177_/D VGND VGND VPWR VPWR _36177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33389_ _36079_/CLK _33389_/D VGND VGND VPWR VPWR _33389_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_363_CLK clkbuf_6_44__f_CLK/X VGND VGND VPWR VPWR _35193_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_147_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23142_ _22962_/X _32110_/Q _23152_/S VGND VGND VPWR VPWR _23143_/A sky130_fd_sc_hd__mux2_1
X_20354_ _35662_/Q _35022_/Q _34382_/Q _33742_/Q _20150_/X _20151_/X VGND VGND VPWR
+ VPWR _20354_/X sky130_fd_sc_hd__mux4_1
X_35128_ _35192_/CLK _35128_/D VGND VGND VPWR VPWR _35128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27950_ _27950_/A VGND VGND VPWR VPWR _34313_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_115_CLK clkbuf_6_20__f_CLK/X VGND VGND VPWR VPWR _35610_/CLK sky130_fd_sc_hd__clkbuf_16
X_23073_ input57/X VGND VGND VPWR VPWR _23073_/X sky130_fd_sc_hd__buf_2
X_35059_ _36146_/CLK _35059_/D VGND VGND VPWR VPWR _35059_/Q sky130_fd_sc_hd__dfxtp_1
X_20285_ _20065_/X _20283_/X _20284_/X _20071_/X VGND VGND VPWR VPWR _20285_/X sky130_fd_sc_hd__a22o_1
XTAP_6206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26901_ _26901_/A VGND VGND VPWR VPWR _33878_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22024_ _22515_/A VGND VGND VPWR VPWR _22024_/X sky130_fd_sc_hd__clkbuf_4
XTAP_6239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27881_ _27701_/X _34281_/Q _27881_/S VGND VGND VPWR VPWR _27882_/A sky130_fd_sc_hd__mux2_1
XTAP_5516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29620_ _29620_/A VGND VGND VPWR VPWR _35073_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_216_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26832_ _33846_/Q _23396_/X _26846_/S VGND VGND VPWR VPWR _26833_/A sky130_fd_sc_hd__mux2_1
XTAP_5549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29551_ _29551_/A VGND VGND VPWR VPWR _35040_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26763_ _30202_/A _31688_/B VGND VGND VPWR VPWR _26896_/S sky130_fd_sc_hd__nor2_8
XTAP_4859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23975_ _23079_/X _32532_/Q _23977_/S VGND VGND VPWR VPWR _23976_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_1015 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28502_ _28502_/A VGND VGND VPWR VPWR _34575_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25714_ _24852_/X _33319_/Q _25718_/S VGND VGND VPWR VPWR _25715_/A sky130_fd_sc_hd__mux2_1
X_29482_ _35015_/Q _29481_/X _29482_/S VGND VGND VPWR VPWR _29483_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22926_ _22925_/X _32034_/Q _22947_/S VGND VGND VPWR VPWR _22927_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26694_ _26694_/A VGND VGND VPWR VPWR _33780_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28433_ _28433_/A VGND VGND VPWR VPWR _34542_/D sky130_fd_sc_hd__clkbuf_1
X_25645_ _25645_/A VGND VGND VPWR VPWR _33286_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22857_ _33173_/Q _36053_/Q _33045_/Q _32981_/Q _20632_/X _21761_/A VGND VGND VPWR
+ VPWR _22857_/X sky130_fd_sc_hd__mux4_1
XFILLER_231_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28364_ _27816_/X _34510_/Q _28370_/S VGND VGND VPWR VPWR _28365_/A sky130_fd_sc_hd__mux2_1
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21808_ _33910_/Q _33846_/Q _33782_/Q _36086_/Q _21624_/X _21625_/X VGND VGND VPWR
+ VPWR _21808_/X sky130_fd_sc_hd__mux4_1
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25576_ _25576_/A VGND VGND VPWR VPWR _33253_/D sky130_fd_sc_hd__clkbuf_1
X_22788_ _22788_/A VGND VGND VPWR VPWR _36242_/D sky130_fd_sc_hd__clkbuf_1
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27315_ _34044_/Q _27152_/X _27317_/S VGND VGND VPWR VPWR _27316_/A sky130_fd_sc_hd__mux2_1
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24527_ _24659_/S VGND VGND VPWR VPWR _24546_/S sky130_fd_sc_hd__buf_6
XFILLER_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28295_ _27714_/X _34477_/Q _28307_/S VGND VGND VPWR VPWR _28296_/A sky130_fd_sc_hd__mux2_1
X_21739_ _21667_/X _21737_/X _21738_/X _21671_/X VGND VGND VPWR VPWR _21739_/X sky130_fd_sc_hd__a22o_1
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27246_ _34011_/Q _27050_/X _27254_/S VGND VGND VPWR VPWR _27247_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24458_ _22984_/X _32757_/Q _24474_/S VGND VGND VPWR VPWR _24459_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23409_ _32215_/Q _23408_/X _23418_/S VGND VGND VPWR VPWR _23410_/A sky130_fd_sc_hd__mux2_1
X_27177_ input41/X VGND VGND VPWR VPWR _27177_/X sky130_fd_sc_hd__buf_4
XFILLER_126_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_354_CLK clkbuf_6_46__f_CLK/X VGND VGND VPWR VPWR _35581_/CLK sky130_fd_sc_hd__clkbuf_16
X_24389_ _23082_/X _32725_/Q _24389_/S VGND VGND VPWR VPWR _24390_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26128_ _24865_/X _33515_/Q _26144_/S VGND VGND VPWR VPWR _26129_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26059_ _26059_/A VGND VGND VPWR VPWR _33482_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_106_CLK clkbuf_leaf_81_CLK/A VGND VGND VPWR VPWR _36059_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_140_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18950_ _20164_/A VGND VGND VPWR VPWR _18950_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_79_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17901_ _17864_/X _17899_/X _17900_/X _17869_/X VGND VGND VPWR VPWR _17901_/X sky130_fd_sc_hd__a22o_1
XFILLER_3_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18881_ _18592_/X _18879_/X _18880_/X _18595_/X VGND VGND VPWR VPWR _18881_/X sky130_fd_sc_hd__a22o_1
XTAP_6740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17832_ _17552_/X _17830_/X _17831_/X _17557_/X VGND VGND VPWR VPWR _17832_/X sky130_fd_sc_hd__a22o_1
XTAP_6773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29818_ _29818_/A VGND VGND VPWR VPWR _35167_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17763_ _17559_/X _17761_/X _17762_/X _17562_/X VGND VGND VPWR VPWR _17763_/X sky130_fd_sc_hd__a22o_1
XFILLER_43_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29749_ _29749_/A VGND VGND VPWR VPWR _35134_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19502_ _33654_/Q _33590_/Q _33526_/Q _33462_/Q _19500_/X _19501_/X VGND VGND VPWR
+ VPWR _19502_/X sky130_fd_sc_hd__mux4_1
X_16714_ _17912_/A VGND VGND VPWR VPWR _16714_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_35_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32760_ _32887_/CLK _32760_/D VGND VGND VPWR VPWR _32760_/Q sky130_fd_sc_hd__dfxtp_1
X_17694_ _17690_/X _17693_/X _17485_/X VGND VGND VPWR VPWR _17724_/A sky130_fd_sc_hd__o21ba_1
XFILLER_19_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_778 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19433_ _19426_/X _19431_/X _19432_/X VGND VGND VPWR VPWR _19467_/A sky130_fd_sc_hd__o21ba_1
X_31711_ _36064_/Q input2/X _31729_/S VGND VGND VPWR VPWR _31712_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16645_ _17859_/A VGND VGND VPWR VPWR _16645_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_78_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32691_ _32906_/CLK _32691_/D VGND VGND VPWR VPWR _32691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34430_ _36103_/CLK _34430_/D VGND VGND VPWR VPWR _34430_/Q sky130_fd_sc_hd__dfxtp_1
X_31642_ _31642_/A VGND VGND VPWR VPWR _36031_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19364_ _33138_/Q _36018_/Q _33010_/Q _32946_/Q _19362_/X _19363_/X VGND VGND VPWR
+ VPWR _19364_/X sky130_fd_sc_hd__mux4_1
X_16576_ _32868_/Q _32804_/Q _32740_/Q _32676_/Q _16287_/X _16288_/X VGND VGND VPWR
+ VPWR _16576_/X sky130_fd_sc_hd__mux4_1
XFILLER_76_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18315_ _20138_/A VGND VGND VPWR VPWR _18315_/X sky130_fd_sc_hd__buf_4
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34361_ _35769_/CLK _34361_/D VGND VGND VPWR VPWR _34361_/Q sky130_fd_sc_hd__dfxtp_1
X_31573_ _27670_/X _35999_/Q _31573_/S VGND VGND VPWR VPWR _31574_/A sky130_fd_sc_hd__mux2_1
X_19295_ _32880_/Q _32816_/Q _32752_/Q _32688_/Q _19293_/X _19294_/X VGND VGND VPWR
+ VPWR _19295_/X sky130_fd_sc_hd__mux4_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_1249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36100_ _36100_/CLK _36100_/D VGND VGND VPWR VPWR _36100_/Q sky130_fd_sc_hd__dfxtp_1
X_33312_ _36066_/CLK _33312_/D VGND VGND VPWR VPWR _33312_/Q sky130_fd_sc_hd__dfxtp_1
X_18246_ _18242_/X _18245_/X _17871_/A VGND VGND VPWR VPWR _18247_/D sky130_fd_sc_hd__o21ba_1
X_30524_ _35502_/Q _29404_/X _30534_/S VGND VGND VPWR VPWR _30525_/A sky130_fd_sc_hd__mux2_1
X_34292_ _34612_/CLK _34292_/D VGND VGND VPWR VPWR _34292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33243_ _35547_/CLK _33243_/D VGND VGND VPWR VPWR _33243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36031_ _36031_/CLK _36031_/D VGND VGND VPWR VPWR _36031_/Q sky130_fd_sc_hd__dfxtp_1
X_30455_ _30455_/A VGND VGND VPWR VPWR _35469_/D sky130_fd_sc_hd__clkbuf_1
X_18177_ _33106_/Q _32082_/Q _35858_/Q _35794_/Q _16079_/X _16080_/X VGND VGND VPWR
+ VPWR _18177_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_345_CLK clkbuf_6_47__f_CLK/X VGND VGND VPWR VPWR _35965_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_129_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_1277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17128_ _17834_/A VGND VGND VPWR VPWR _17128_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_237_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33174_ _35804_/CLK _33174_/D VGND VGND VPWR VPWR _33174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30386_ _30386_/A VGND VGND VPWR VPWR _35436_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_239_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32125_ _32895_/CLK _32125_/D VGND VGND VPWR VPWR _32125_/Q sky130_fd_sc_hd__dfxtp_1
X_17059_ _17905_/A VGND VGND VPWR VPWR _17059_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_239_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20070_ _33158_/Q _36038_/Q _33030_/Q _32966_/Q _20068_/X _20069_/X VGND VGND VPWR
+ VPWR _20070_/X sky130_fd_sc_hd__mux4_1
XFILLER_131_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32056_ _35768_/CLK _32056_/D VGND VGND VPWR VPWR _32056_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31007_ _31007_/A VGND VGND VPWR VPWR _35731_/D sky130_fd_sc_hd__clkbuf_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35815_ _35943_/CLK _35815_/D VGND VGND VPWR VPWR _35815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20972_ _22535_/A VGND VGND VPWR VPWR _20972_/X sky130_fd_sc_hd__buf_6
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35746_ _35812_/CLK _35746_/D VGND VGND VPWR VPWR _35746_/Q sky130_fd_sc_hd__dfxtp_1
X_23760_ _23760_/A VGND VGND VPWR VPWR _32366_/D sky130_fd_sc_hd__clkbuf_1
X_32958_ _35839_/CLK _32958_/D VGND VGND VPWR VPWR _32958_/Q sky130_fd_sc_hd__dfxtp_1
X_22711_ _21758_/A _22709_/X _22710_/X _21763_/A VGND VGND VPWR VPWR _22711_/X sky130_fd_sc_hd__a22o_1
X_31909_ _23420_/X _36158_/Q _31927_/S VGND VGND VPWR VPWR _31910_/A sky130_fd_sc_hd__mux2_1
XFILLER_226_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35677_ _35677_/CLK _35677_/D VGND VGND VPWR VPWR _35677_/Q sky130_fd_sc_hd__dfxtp_1
X_23691_ _23691_/A VGND VGND VPWR VPWR _32335_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32889_ _32889_/CLK _32889_/D VGND VGND VPWR VPWR _32889_/Q sky130_fd_sc_hd__dfxtp_1
X_25430_ _24830_/X _33184_/Q _25448_/S VGND VGND VPWR VPWR _25431_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22642_ _33422_/Q _33358_/Q _33294_/Q _33230_/Q _22433_/X _22434_/X VGND VGND VPWR
+ VPWR _22642_/X sky130_fd_sc_hd__mux4_1
X_34628_ _36164_/CLK _34628_/D VGND VGND VPWR VPWR _34628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_1130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_910 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22573_ _22573_/A _22573_/B _22573_/C _22573_/D VGND VGND VPWR VPWR _22574_/A sky130_fd_sc_hd__or4_4
X_25361_ _25361_/A VGND VGND VPWR VPWR _33152_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34559_ _35071_/CLK _34559_/D VGND VGND VPWR VPWR _34559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_1046 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27100_ input14/X VGND VGND VPWR VPWR _27100_/X sky130_fd_sc_hd__buf_2
X_24312_ _22968_/X _32688_/Q _24318_/S VGND VGND VPWR VPWR _24313_/A sky130_fd_sc_hd__mux2_1
X_28080_ _28080_/A VGND VGND VPWR VPWR _34375_/D sky130_fd_sc_hd__clkbuf_1
X_21524_ _32622_/Q _32558_/Q _32494_/Q _35950_/Q _21523_/X _21307_/X VGND VGND VPWR
+ VPWR _21524_/X sky130_fd_sc_hd__mux4_1
X_25292_ _25403_/S VGND VGND VPWR VPWR _25311_/S sky130_fd_sc_hd__buf_4
XFILLER_210_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27031_ _33941_/Q _23498_/X _27031_/S VGND VGND VPWR VPWR _27032_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_903 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36229_ _36229_/CLK _36229_/D VGND VGND VPWR VPWR _36229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24243_ _32657_/Q _23484_/X _24243_/S VGND VGND VPWR VPWR _24244_/A sky130_fd_sc_hd__mux2_1
X_21455_ _33900_/Q _33836_/Q _33772_/Q _36076_/Q _21271_/X _21272_/X VGND VGND VPWR
+ VPWR _21455_/X sky130_fd_sc_hd__mux4_1
XFILLER_215_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_336_CLK clkbuf_6_44__f_CLK/X VGND VGND VPWR VPWR _36027_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_135_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20406_ _32656_/Q _32592_/Q _32528_/Q _35984_/Q _20282_/X _19177_/A VGND VGND VPWR
+ VPWR _20406_/X sky130_fd_sc_hd__mux4_1
XFILLER_147_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24174_ _32624_/Q _23340_/X _24180_/S VGND VGND VPWR VPWR _24175_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21386_ _21314_/X _21384_/X _21385_/X _21318_/X VGND VGND VPWR VPWR _21386_/X sky130_fd_sc_hd__a22o_1
XFILLER_200_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20337_ _20337_/A _20337_/B _20337_/C _20337_/D VGND VGND VPWR VPWR _20338_/A sky130_fd_sc_hd__or4_1
X_23125_ _22937_/X _32102_/Q _23131_/S VGND VGND VPWR VPWR _23126_/A sky130_fd_sc_hd__mux2_1
X_28982_ _28982_/A VGND VGND VPWR VPWR _34801_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27933_ _27933_/A VGND VGND VPWR VPWR _34305_/D sky130_fd_sc_hd__clkbuf_1
X_23056_ _23055_/X _32076_/Q _23071_/S VGND VGND VPWR VPWR _23057_/A sky130_fd_sc_hd__mux2_1
X_20268_ _20159_/X _20266_/X _20267_/X _20162_/X VGND VGND VPWR VPWR _20268_/X sky130_fd_sc_hd__a22o_1
XTAP_6025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22007_ _21799_/X _22005_/X _22006_/X _21804_/X VGND VGND VPWR VPWR _22007_/X sky130_fd_sc_hd__a22o_1
XTAP_6069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27864_ _27864_/A VGND VGND VPWR VPWR _34272_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20199_ _34441_/Q _36169_/Q _34313_/Q _34249_/Q _19882_/X _19883_/X VGND VGND VPWR
+ VPWR _20199_/X sky130_fd_sc_hd__mux4_1
XTAP_4601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26815_ _33838_/Q _23305_/X _26825_/S VGND VGND VPWR VPWR _26816_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_1020 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29603_ _29603_/A VGND VGND VPWR VPWR _35065_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27795_ _27794_/X _34247_/Q _27795_/S VGND VGND VPWR VPWR _27796_/A sky130_fd_sc_hd__mux2_1
XTAP_4645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29534_ _29534_/A VGND VGND VPWR VPWR _35032_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26746_ _26746_/A VGND VGND VPWR VPWR _33805_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_217_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23958_ _23958_/A VGND VGND VPWR VPWR _32523_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29465_ _29465_/A VGND VGND VPWR VPWR _35009_/D sky130_fd_sc_hd__clkbuf_1
X_22909_ input62/X VGND VGND VPWR VPWR _22909_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26677_ _26677_/A VGND VGND VPWR VPWR _33772_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23889_ _23889_/A VGND VGND VPWR VPWR _32490_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_189_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16430_ _16353_/X _16428_/X _16429_/X _16359_/X VGND VGND VPWR VPWR _16430_/X sky130_fd_sc_hd__a22o_1
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28416_ _28416_/A VGND VGND VPWR VPWR _34534_/D sky130_fd_sc_hd__clkbuf_1
X_25628_ _24923_/X _33278_/Q _25646_/S VGND VGND VPWR VPWR _25629_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29396_ _34987_/Q _29395_/X _29420_/S VGND VGND VPWR VPWR _29397_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28347_ _27791_/X _34502_/Q _28349_/S VGND VGND VPWR VPWR _28348_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16361_ _17912_/A VGND VGND VPWR VPWR _16361_/X sky130_fd_sc_hd__clkbuf_4
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25559_ _25559_/A VGND VGND VPWR VPWR _33245_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18100_ _34192_/Q _34128_/Q _34064_/Q _34000_/Q _17799_/X _17800_/X VGND VGND VPWR
+ VPWR _18100_/X sky130_fd_sc_hd__mux4_1
XFILLER_164_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19080_ _19073_/X _19078_/X _19079_/X VGND VGND VPWR VPWR _19114_/A sky130_fd_sc_hd__o21ba_1
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16292_ _17859_/A VGND VGND VPWR VPWR _16292_/X sky130_fd_sc_hd__buf_4
XFILLER_13_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28278_ _27689_/X _34469_/Q _28286_/S VGND VGND VPWR VPWR _28279_/A sky130_fd_sc_hd__mux2_1
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18031_ _35213_/Q _35149_/Q _35085_/Q _32269_/Q _17716_/X _17717_/X VGND VGND VPWR
+ VPWR _18031_/X sky130_fd_sc_hd__mux4_1
XFILLER_199_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27229_ input60/X VGND VGND VPWR VPWR _27229_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_172_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_327_CLK clkbuf_6_39__f_CLK/X VGND VGND VPWR VPWR _35895_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_138_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30240_ _30240_/A VGND VGND VPWR VPWR _35367_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30171_ _35335_/Q _29481_/X _30171_/S VGND VGND VPWR VPWR _30172_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19982_ _34435_/Q _36163_/Q _34307_/Q _34243_/Q _19882_/X _19883_/X VGND VGND VPWR
+ VPWR _19982_/X sky130_fd_sc_hd__mux4_1
XFILLER_141_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18933_ _33894_/Q _33830_/Q _33766_/Q _36070_/Q _18618_/X _18619_/X VGND VGND VPWR
+ VPWR _18933_/X sky130_fd_sc_hd__mux4_1
XFILLER_45_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33930_ _36105_/CLK _33930_/D VGND VGND VPWR VPWR _33930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_1365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18864_ _34148_/Q _34084_/Q _34020_/Q _33956_/Q _18687_/X _18688_/X VGND VGND VPWR
+ VPWR _18864_/X sky130_fd_sc_hd__mux4_1
XFILLER_95_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17815_ _35655_/Q _35015_/Q _34375_/Q _33735_/Q _17497_/X _17498_/X VGND VGND VPWR
+ VPWR _17815_/X sky130_fd_sc_hd__mux4_1
X_33861_ _34177_/CLK _33861_/D VGND VGND VPWR VPWR _33861_/Q sky130_fd_sc_hd__dfxtp_1
X_18795_ _20207_/A VGND VGND VPWR VPWR _18795_/X sky130_fd_sc_hd__buf_4
XFILLER_39_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35600_ _35729_/CLK _35600_/D VGND VGND VPWR VPWR _35600_/Q sky130_fd_sc_hd__dfxtp_1
X_17746_ _33093_/Q _32069_/Q _35845_/Q _35781_/Q _17431_/X _17432_/X VGND VGND VPWR
+ VPWR _17746_/X sky130_fd_sc_hd__mux4_1
X_32812_ _32914_/CLK _32812_/D VGND VGND VPWR VPWR _32812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_242_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33792_ _36096_/CLK _33792_/D VGND VGND VPWR VPWR _33792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_247_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35531_ _35596_/CLK _35531_/D VGND VGND VPWR VPWR _35531_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17677_ _17356_/X _17675_/X _17676_/X _17359_/X VGND VGND VPWR VPWR _17677_/X sky130_fd_sc_hd__a22o_1
X_32743_ _32871_/CLK _32743_/D VGND VGND VPWR VPWR _32743_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16628_ _16628_/A VGND VGND VPWR VPWR _31973_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19416_ _35187_/Q _35123_/Q _35059_/Q _32220_/Q _19310_/X _19311_/X VGND VGND VPWR
+ VPWR _19416_/X sky130_fd_sc_hd__mux4_1
X_35462_ _35463_/CLK _35462_/D VGND VGND VPWR VPWR _35462_/Q sky130_fd_sc_hd__dfxtp_1
X_32674_ _35871_/CLK _32674_/D VGND VGND VPWR VPWR _32674_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34413_ _34413_/CLK _34413_/D VGND VGND VPWR VPWR _34413_/Q sky130_fd_sc_hd__dfxtp_1
X_31625_ _31625_/A VGND VGND VPWR VPWR _36023_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_245_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19347_ _34929_/Q _34865_/Q _34801_/Q _34737_/Q _19107_/X _19108_/X VGND VGND VPWR
+ VPWR _19347_/X sky130_fd_sc_hd__mux4_1
X_16559_ _16452_/X _16557_/X _16558_/X _16457_/X VGND VGND VPWR VPWR _16559_/X sky130_fd_sc_hd__a22o_1
XFILLER_206_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35393_ _35458_/CLK _35393_/D VGND VGND VPWR VPWR _35393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31556_ _31556_/A VGND VGND VPWR VPWR _35990_/D sky130_fd_sc_hd__clkbuf_1
X_34344_ _35559_/CLK _34344_/D VGND VGND VPWR VPWR _34344_/Q sky130_fd_sc_hd__dfxtp_1
X_19278_ _19105_/X _19276_/X _19277_/X _19110_/X VGND VGND VPWR VPWR _19278_/X sky130_fd_sc_hd__a22o_1
XFILLER_104_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18229_ _32148_/Q _32340_/Q _32404_/Q _35924_/Q _17986_/X _17011_/A VGND VGND VPWR
+ VPWR _18229_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30507_ _35494_/Q _29379_/X _30513_/S VGND VGND VPWR VPWR _30508_/A sky130_fd_sc_hd__mux2_1
XFILLER_175_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_318_CLK clkbuf_6_37__f_CLK/X VGND VGND VPWR VPWR _32907_/CLK sky130_fd_sc_hd__clkbuf_16
X_34275_ _34405_/CLK _34275_/D VGND VGND VPWR VPWR _34275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31487_ _27742_/X _35958_/Q _31501_/S VGND VGND VPWR VPWR _31488_/A sky130_fd_sc_hd__mux2_1
X_33226_ _33673_/CLK _33226_/D VGND VGND VPWR VPWR _33226_/Q sky130_fd_sc_hd__dfxtp_1
X_21240_ _22433_/A VGND VGND VPWR VPWR _21240_/X sky130_fd_sc_hd__buf_4
X_36014_ _36015_/CLK _36014_/D VGND VGND VPWR VPWR _36014_/Q sky130_fd_sc_hd__dfxtp_1
X_30438_ _30438_/A VGND VGND VPWR VPWR _35461_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33157_ _36037_/CLK _33157_/D VGND VGND VPWR VPWR _33157_/Q sky130_fd_sc_hd__dfxtp_1
X_21171_ _32612_/Q _32548_/Q _32484_/Q _35940_/Q _21170_/X _20954_/X VGND VGND VPWR
+ VPWR _21171_/X sky130_fd_sc_hd__mux4_1
X_30369_ _30369_/A VGND VGND VPWR VPWR _35428_/D sky130_fd_sc_hd__clkbuf_1
X_20122_ _35207_/Q _35143_/Q _35079_/Q _32263_/Q _20016_/X _20017_/X VGND VGND VPWR
+ VPWR _20122_/X sky130_fd_sc_hd__mux4_1
X_32108_ _35949_/CLK _32108_/D VGND VGND VPWR VPWR _32108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33088_ _35713_/CLK _33088_/D VGND VGND VPWR VPWR _33088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20053_ _34949_/Q _34885_/Q _34821_/Q _34757_/Q _19813_/X _19814_/X VGND VGND VPWR
+ VPWR _20053_/X sky130_fd_sc_hd__mux4_1
X_24930_ input37/X VGND VGND VPWR VPWR _24930_/X sky130_fd_sc_hd__clkbuf_4
X_32039_ _35943_/CLK _32039_/D VGND VGND VPWR VPWR _32039_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24861_ input13/X VGND VGND VPWR VPWR _24861_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_100_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26600_ _24961_/X _33738_/Q _26614_/S VGND VGND VPWR VPWR _26601_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23812_ _23812_/A VGND VGND VPWR VPWR _32391_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27580_ _27580_/A VGND VGND VPWR VPWR _34169_/D sky130_fd_sc_hd__clkbuf_1
X_24792_ _23079_/X _32916_/Q _24794_/S VGND VGND VPWR VPWR _24793_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26531_ _26531_/A VGND VGND VPWR VPWR _33705_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35729_ _35729_/CLK _35729_/D VGND VGND VPWR VPWR _35729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23743_ _23743_/A VGND VGND VPWR VPWR _32358_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_214_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20955_ _32606_/Q _32542_/Q _32478_/Q _35934_/Q _20817_/X _20954_/X VGND VGND VPWR
+ VPWR _20955_/X sky130_fd_sc_hd__mux4_1
XFILLER_27_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29250_ _29250_/A VGND VGND VPWR VPWR _34928_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26462_ _33673_/Q _23460_/X _26478_/S VGND VGND VPWR VPWR _26463_/A sky130_fd_sc_hd__mux2_1
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23674_ _23674_/A VGND VGND VPWR VPWR _32327_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20886_ _32092_/Q _32284_/Q _32348_/Q _35868_/Q _20821_/X _22467_/A VGND VGND VPWR
+ VPWR _20886_/X sky130_fd_sc_hd__mux4_1
XFILLER_214_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28201_ _28201_/A VGND VGND VPWR VPWR _34432_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25413_ _24806_/X _33176_/Q _25427_/S VGND VGND VPWR VPWR _25414_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29181_ _34896_/Q _27214_/X _29183_/S VGND VGND VPWR VPWR _29182_/A sky130_fd_sc_hd__mux2_1
X_22625_ _22304_/X _22623_/X _22624_/X _22307_/X VGND VGND VPWR VPWR _22625_/X sky130_fd_sc_hd__a22o_1
XFILLER_167_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26393_ _26393_/A VGND VGND VPWR VPWR _33640_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28132_ _28243_/S VGND VGND VPWR VPWR _28151_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_195_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25344_ _25344_/A VGND VGND VPWR VPWR _33144_/D sky130_fd_sc_hd__clkbuf_1
X_22556_ _22552_/X _22555_/X _22446_/X _22447_/X VGND VGND VPWR VPWR _22573_/B sky130_fd_sc_hd__o211a_2
XFILLER_166_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28063_ _34367_/Q _27162_/X _28079_/S VGND VGND VPWR VPWR _28064_/A sky130_fd_sc_hd__mux2_1
X_21507_ _34669_/Q _34605_/Q _34541_/Q _34477_/Q _21186_/X _21187_/X VGND VGND VPWR
+ VPWR _21507_/X sky130_fd_sc_hd__mux4_1
X_25275_ _25275_/A VGND VGND VPWR VPWR _33111_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_309_CLK clkbuf_6_50__f_CLK/X VGND VGND VPWR VPWR _35973_/CLK sky130_fd_sc_hd__clkbuf_16
X_22487_ _22373_/X _22485_/X _22486_/X _22377_/X VGND VGND VPWR VPWR _22487_/X sky130_fd_sc_hd__a22o_1
XFILLER_182_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27014_ _27014_/A VGND VGND VPWR VPWR _33932_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24226_ _24226_/A VGND VGND VPWR VPWR _32648_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21438_ _35179_/Q _35115_/Q _35051_/Q _32171_/Q _21257_/X _21258_/X VGND VGND VPWR
+ VPWR _21438_/X sky130_fd_sc_hd__mux4_1
XFILLER_181_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21369_ _21369_/A _21369_/B _21369_/C _21369_/D VGND VGND VPWR VPWR _21370_/A sky130_fd_sc_hd__or4_4
X_24157_ _32616_/Q _23286_/X _24159_/S VGND VGND VPWR VPWR _24158_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23108_ _22912_/X _32094_/Q _23110_/S VGND VGND VPWR VPWR _23109_/A sky130_fd_sc_hd__mux2_1
X_24088_ _24088_/A VGND VGND VPWR VPWR _32584_/D sky130_fd_sc_hd__clkbuf_1
X_28965_ _28965_/A VGND VGND VPWR VPWR _34793_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23039_ input44/X VGND VGND VPWR VPWR _23039_/X sky130_fd_sc_hd__buf_2
X_27916_ _27916_/A VGND VGND VPWR VPWR _34297_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28896_ _28896_/A VGND VGND VPWR VPWR _34760_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27847_ _27847_/A VGND VGND VPWR VPWR _34264_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17600_ _32129_/Q _32321_/Q _32385_/Q _35905_/Q _17280_/X _17421_/X VGND VGND VPWR
+ VPWR _17600_/X sky130_fd_sc_hd__mux4_1
XFILLER_114_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_218_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18580_ _33884_/Q _33820_/Q _33756_/Q _36060_/Q _18412_/X _18413_/X VGND VGND VPWR
+ VPWR _18580_/X sky130_fd_sc_hd__mux4_1
XTAP_4464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27778_ _27778_/A VGND VGND VPWR VPWR _34241_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17531_ _17412_/X _17529_/X _17530_/X _17418_/X VGND VGND VPWR VPWR _17531_/X sky130_fd_sc_hd__a22o_1
X_26729_ _26729_/A VGND VGND VPWR VPWR _33797_/D sky130_fd_sc_hd__clkbuf_1
X_29517_ _29517_/A VGND VGND VPWR VPWR _35026_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17462_ _35645_/Q _35005_/Q _34365_/Q _33725_/Q _17144_/X _17145_/X VGND VGND VPWR
+ VPWR _17462_/X sky130_fd_sc_hd__mux4_1
X_29448_ _35004_/Q _29447_/X _29451_/S VGND VGND VPWR VPWR _29449_/A sky130_fd_sc_hd__mux2_1
XFILLER_229_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16413_ _34911_/Q _34847_/Q _34783_/Q _34719_/Q _16096_/X _16098_/X VGND VGND VPWR
+ VPWR _16413_/X sky130_fd_sc_hd__mux4_1
X_19201_ _20260_/A VGND VGND VPWR VPWR _19201_/X sky130_fd_sc_hd__buf_4
XFILLER_177_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29379_ input8/X VGND VGND VPWR VPWR _29379_/X sky130_fd_sc_hd__buf_2
X_17393_ _33083_/Q _32059_/Q _35835_/Q _35771_/Q _17078_/X _17079_/X VGND VGND VPWR
+ VPWR _17393_/X sky130_fd_sc_hd__mux4_1
XFILLER_13_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31410_ _27828_/X _35922_/Q _31416_/S VGND VGND VPWR VPWR _31411_/A sky130_fd_sc_hd__mux2_1
X_19132_ _18945_/X _19130_/X _19131_/X _18948_/X VGND VGND VPWR VPWR _19132_/X sky130_fd_sc_hd__a22o_1
XFILLER_157_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16344_ _16344_/A _16344_/B _16344_/C _16344_/D VGND VGND VPWR VPWR _16345_/A sky130_fd_sc_hd__or4_4
XFILLER_73_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32390_ _35976_/CLK _32390_/D VGND VGND VPWR VPWR _32390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_242_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19063_ _35177_/Q _35113_/Q _35049_/Q _32169_/Q _18957_/X _18958_/X VGND VGND VPWR
+ VPWR _19063_/X sky130_fd_sc_hd__mux4_1
X_31341_ _27726_/X _35889_/Q _31345_/S VGND VGND VPWR VPWR _31342_/A sky130_fd_sc_hd__mux2_1
X_16275_ _16275_/A VGND VGND VPWR VPWR _31963_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_173_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_1361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18014_ _17912_/X _18012_/X _18013_/X _17915_/X VGND VGND VPWR VPWR _18014_/X sky130_fd_sc_hd__a22o_1
X_34060_ _34188_/CLK _34060_/D VGND VGND VPWR VPWR _34060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31272_ _31272_/A VGND VGND VPWR VPWR _35856_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33011_ _36019_/CLK _33011_/D VGND VGND VPWR VPWR _33011_/Q sky130_fd_sc_hd__dfxtp_1
X_30223_ _30223_/A VGND VGND VPWR VPWR _35359_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30154_ _30154_/A VGND VGND VPWR VPWR _35326_/D sky130_fd_sc_hd__clkbuf_1
X_19965_ _19712_/X _19963_/X _19964_/X _19718_/X VGND VGND VPWR VPWR _19965_/X sky130_fd_sc_hd__a22o_1
XFILLER_45_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18916_ _35429_/Q _35365_/Q _35301_/Q _35237_/Q _18848_/X _18849_/X VGND VGND VPWR
+ VPWR _18916_/X sky130_fd_sc_hd__mux4_1
XTAP_7090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34962_ _34964_/CLK _34962_/D VGND VGND VPWR VPWR _34962_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30085_ _35294_/Q _29354_/X _30087_/S VGND VGND VPWR VPWR _30086_/A sky130_fd_sc_hd__mux2_1
X_19896_ _19892_/X _19895_/X _19785_/X VGND VGND VPWR VPWR _19920_/A sky130_fd_sc_hd__o21ba_1
X_33913_ _33913_/CLK _33913_/D VGND VGND VPWR VPWR _33913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18847_ _18592_/X _18845_/X _18846_/X _18595_/X VGND VGND VPWR VPWR _18847_/X sky130_fd_sc_hd__a22o_1
X_34893_ _34957_/CLK _34893_/D VGND VGND VPWR VPWR _34893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_243_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33844_ _34100_/CLK _33844_/D VGND VGND VPWR VPWR _33844_/Q sky130_fd_sc_hd__dfxtp_1
X_18778_ _35617_/Q _34977_/Q _34337_/Q _33697_/Q _18738_/X _18739_/X VGND VGND VPWR
+ VPWR _18778_/X sky130_fd_sc_hd__mux4_2
XFILLER_94_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17729_ _33413_/Q _33349_/Q _33285_/Q _33221_/Q _17480_/X _17481_/X VGND VGND VPWR
+ VPWR _17729_/X sky130_fd_sc_hd__mux4_1
XFILLER_82_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30987_ _30987_/A VGND VGND VPWR VPWR _35721_/D sky130_fd_sc_hd__clkbuf_1
X_33775_ _36079_/CLK _33775_/D VGND VGND VPWR VPWR _33775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_242_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35514_ _35581_/CLK _35514_/D VGND VGND VPWR VPWR _35514_/Q sky130_fd_sc_hd__dfxtp_1
X_32726_ _32856_/CLK _32726_/D VGND VGND VPWR VPWR _32726_/Q sky130_fd_sc_hd__dfxtp_1
X_20740_ _22459_/A VGND VGND VPWR VPWR _20740_/X sky130_fd_sc_hd__buf_4
XFILLER_35_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20671_ _22377_/A VGND VGND VPWR VPWR _22469_/A sky130_fd_sc_hd__buf_12
X_35445_ _35446_/CLK _35445_/D VGND VGND VPWR VPWR _35445_/Q sky130_fd_sc_hd__dfxtp_1
X_32657_ _36049_/CLK _32657_/D VGND VGND VPWR VPWR _32657_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_95_CLK clkbuf_leaf_96_CLK/A VGND VGND VPWR VPWR _36188_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_143_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22410_ _32135_/Q _32327_/Q _32391_/Q _35911_/Q _22233_/X _22374_/X VGND VGND VPWR
+ VPWR _22410_/X sky130_fd_sc_hd__mux4_1
XFILLER_32_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31608_ _31608_/A VGND VGND VPWR VPWR _36015_/D sky130_fd_sc_hd__clkbuf_1
X_32588_ _35980_/CLK _32588_/D VGND VGND VPWR VPWR _32588_/Q sky130_fd_sc_hd__dfxtp_1
X_23390_ _23390_/A VGND VGND VPWR VPWR _32208_/D sky130_fd_sc_hd__clkbuf_1
X_35376_ _35634_/CLK _35376_/D VGND VGND VPWR VPWR _35376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34327_ _35674_/CLK _34327_/D VGND VGND VPWR VPWR _34327_/Q sky130_fd_sc_hd__dfxtp_1
X_22341_ _22337_/X _22340_/X _22093_/X _22094_/X VGND VGND VPWR VPWR _22356_/B sky130_fd_sc_hd__o211a_1
XFILLER_136_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31539_ _27819_/X _35983_/Q _31543_/S VGND VGND VPWR VPWR _31540_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22272_ _35715_/Q _32225_/Q _35587_/Q _35523_/Q _22270_/X _22271_/X VGND VGND VPWR
+ VPWR _22272_/X sky130_fd_sc_hd__mux4_1
XFILLER_163_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25060_ _25060_/A VGND VGND VPWR VPWR _33011_/D sky130_fd_sc_hd__clkbuf_1
X_34258_ _34964_/CLK _34258_/D VGND VGND VPWR VPWR _34258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21223_ _34405_/Q _36133_/Q _34277_/Q _34213_/Q _21123_/X _21124_/X VGND VGND VPWR
+ VPWR _21223_/X sky130_fd_sc_hd__mux4_1
XFILLER_89_1081 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24011_ _22931_/X _32548_/Q _24021_/S VGND VGND VPWR VPWR _24012_/A sky130_fd_sc_hd__mux2_1
X_33209_ _36090_/CLK _33209_/D VGND VGND VPWR VPWR _33209_/Q sky130_fd_sc_hd__dfxtp_1
X_34189_ _34193_/CLK _34189_/D VGND VGND VPWR VPWR _34189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21154_ _34659_/Q _34595_/Q _34531_/Q _34467_/Q _20833_/X _20834_/X VGND VGND VPWR
+ VPWR _21154_/X sky130_fd_sc_hd__mux4_1
XFILLER_104_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20105_ _19859_/X _20103_/X _20104_/X _19862_/X VGND VGND VPWR VPWR _20105_/X sky130_fd_sc_hd__a22o_1
XFILLER_120_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28750_ _28750_/A VGND VGND VPWR VPWR _34692_/D sky130_fd_sc_hd__clkbuf_1
X_25962_ _25962_/A VGND VGND VPWR VPWR _33436_/D sky130_fd_sc_hd__clkbuf_1
X_21085_ _35169_/Q _35105_/Q _35041_/Q _32161_/Q _20904_/X _20905_/X VGND VGND VPWR
+ VPWR _21085_/X sky130_fd_sc_hd__mux4_1
XFILLER_150_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27701_ input11/X VGND VGND VPWR VPWR _27701_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_189_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20036_ _33157_/Q _36037_/Q _33029_/Q _32965_/Q _19715_/X _19716_/X VGND VGND VPWR
+ VPWR _20036_/X sky130_fd_sc_hd__mux4_1
XFILLER_28_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24913_ _24913_/A VGND VGND VPWR VPWR _32954_/D sky130_fd_sc_hd__clkbuf_1
X_28681_ _28681_/A VGND VGND VPWR VPWR _34659_/D sky130_fd_sc_hd__clkbuf_1
X_25893_ _24917_/X _33404_/Q _25895_/S VGND VGND VPWR VPWR _25894_/A sky130_fd_sc_hd__mux2_1
XTAP_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27632_ _27632_/A VGND VGND VPWR VPWR _34194_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24844_ _24843_/X _32932_/Q _24859_/S VGND VGND VPWR VPWR _24845_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27563_ _27563_/A VGND VGND VPWR VPWR _34161_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24775_ _24775_/A VGND VGND VPWR VPWR _32907_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_233_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21987_ _21667_/X _21985_/X _21986_/X _21671_/X VGND VGND VPWR VPWR _21987_/X sky130_fd_sc_hd__a22o_1
X_29302_ _34953_/Q _27193_/X _29318_/S VGND VGND VPWR VPWR _29303_/A sky130_fd_sc_hd__mux2_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26514_ _24834_/X _33697_/Q _26530_/S VGND VGND VPWR VPWR _26515_/A sky130_fd_sc_hd__mux2_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23726_ _23726_/A VGND VGND VPWR VPWR _32350_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27494_ _34129_/Q _27217_/X _27494_/S VGND VGND VPWR VPWR _27495_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20938_ _35165_/Q _35101_/Q _35037_/Q _32157_/Q _20904_/X _20905_/X VGND VGND VPWR
+ VPWR _20938_/X sky130_fd_sc_hd__mux4_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_22 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29233_ _29233_/A VGND VGND VPWR VPWR _34920_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26445_ _33665_/Q _23432_/X _26457_/S VGND VGND VPWR VPWR _26446_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_1186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23657_ _23015_/X _32319_/Q _23673_/S VGND VGND VPWR VPWR _23658_/A sky130_fd_sc_hd__mux2_1
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20869_ _20678_/X _20867_/X _20868_/X _20688_/X VGND VGND VPWR VPWR _20869_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_86_CLK clkbuf_leaf_88_CLK/A VGND VGND VPWR VPWR _35807_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_39_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29164_ _29191_/S VGND VGND VPWR VPWR _29183_/S sky130_fd_sc_hd__buf_4
X_22608_ _22608_/A VGND VGND VPWR VPWR _36236_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26376_ _33632_/Q _23261_/X _26394_/S VGND VGND VPWR VPWR _26377_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23588_ _23588_/A VGND VGND VPWR VPWR _32286_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28115_ _28115_/A VGND VGND VPWR VPWR _34391_/D sky130_fd_sc_hd__clkbuf_1
X_25327_ _25327_/A VGND VGND VPWR VPWR _33136_/D sky130_fd_sc_hd__clkbuf_1
X_22539_ _22464_/X _22537_/X _22538_/X _22469_/X VGND VGND VPWR VPWR _22539_/X sky130_fd_sc_hd__a22o_1
XFILLER_182_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29095_ _34855_/Q _27087_/X _29099_/S VGND VGND VPWR VPWR _29096_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16060_ _17864_/A VGND VGND VPWR VPWR _16060_/X sky130_fd_sc_hd__buf_4
X_28046_ _34359_/Q _27137_/X _28058_/S VGND VGND VPWR VPWR _28047_/A sky130_fd_sc_hd__mux2_1
X_25258_ _25258_/A VGND VGND VPWR VPWR _33104_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24209_ _24209_/A VGND VGND VPWR VPWR _32640_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25189_ _25189_/A VGND VGND VPWR VPWR _33071_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_1165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29997_ _35252_/Q _29422_/X _30015_/S VGND VGND VPWR VPWR _29998_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19750_ _33405_/Q _33341_/Q _33277_/Q _33213_/Q _19427_/X _19428_/X VGND VGND VPWR
+ VPWR _19750_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28948_ _34785_/Q _27069_/X _28964_/S VGND VGND VPWR VPWR _28949_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16962_ _16714_/X _16960_/X _16961_/X _16718_/X VGND VGND VPWR VPWR _16962_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_10_CLK clkbuf_leaf_9_CLK/A VGND VGND VPWR VPWR _35618_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_81_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18701_ _18697_/X _18700_/X _18344_/X _18346_/X VGND VGND VPWR VPWR _18716_/B sky130_fd_sc_hd__o211a_1
XFILLER_133_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19681_ _19675_/X _19680_/X _19432_/X VGND VGND VPWR VPWR _19703_/A sky130_fd_sc_hd__o21ba_1
X_16893_ _16706_/X _16891_/X _16892_/X _16712_/X VGND VGND VPWR VPWR _16893_/X sky130_fd_sc_hd__a22o_1
XFILLER_237_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28879_ _28879_/A VGND VGND VPWR VPWR _34752_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18632_ _18592_/X _18630_/X _18631_/X _18595_/X VGND VGND VPWR VPWR _18632_/X sky130_fd_sc_hd__a22o_1
XFILLER_37_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30910_ _35685_/Q input7/X _30918_/S VGND VGND VPWR VPWR _30911_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31890_ _23393_/X _36149_/Q _31906_/S VGND VGND VPWR VPWR _31891_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30841_ _30841_/A VGND VGND VPWR VPWR _35652_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18563_ _35419_/Q _35355_/Q _35291_/Q _35227_/Q _18495_/X _18496_/X VGND VGND VPWR
+ VPWR _18563_/X sky130_fd_sc_hd__mux4_1
XTAP_3560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_1272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17514_ _17867_/A VGND VGND VPWR VPWR _17514_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18494_ _18348_/X _18492_/X _18493_/X _18358_/X VGND VGND VPWR VPWR _18494_/X sky130_fd_sc_hd__a22o_1
X_33560_ _34331_/CLK _33560_/D VGND VGND VPWR VPWR _33560_/Q sky130_fd_sc_hd__dfxtp_1
X_30772_ _30772_/A VGND VGND VPWR VPWR _35619_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32511_ _32575_/CLK _32511_/D VGND VGND VPWR VPWR _32511_/Q sky130_fd_sc_hd__dfxtp_1
X_17445_ _33661_/Q _33597_/Q _33533_/Q _33469_/Q _17200_/X _17201_/X VGND VGND VPWR
+ VPWR _17445_/X sky130_fd_sc_hd__mux4_1
XFILLER_32_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33491_ _34897_/CLK _33491_/D VGND VGND VPWR VPWR _33491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_77_CLK clkbuf_leaf_77_CLK/A VGND VGND VPWR VPWR _35995_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_242_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35230_ _35743_/CLK _35230_/D VGND VGND VPWR VPWR _35230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32442_ _33895_/CLK _32442_/D VGND VGND VPWR VPWR _32442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17376_ _33403_/Q _33339_/Q _33275_/Q _33211_/Q _17127_/X _17128_/X VGND VGND VPWR
+ VPWR _17376_/X sky130_fd_sc_hd__mux4_1
XFILLER_203_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16327_ _32861_/Q _32797_/Q _32733_/Q _32669_/Q _16287_/X _16288_/X VGND VGND VPWR
+ VPWR _16327_/X sky130_fd_sc_hd__mux4_1
X_19115_ _19115_/A VGND VGND VPWR VPWR _32426_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_242_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35161_ _35799_/CLK _35161_/D VGND VGND VPWR VPWR _35161_/Q sky130_fd_sc_hd__dfxtp_1
X_32373_ _32885_/CLK _32373_/D VGND VGND VPWR VPWR _32373_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34112_ _36159_/CLK _34112_/D VGND VGND VPWR VPWR _34112_/Q sky130_fd_sc_hd__dfxtp_1
X_19046_ _18800_/X _19044_/X _19045_/X _18803_/X VGND VGND VPWR VPWR _19046_/X sky130_fd_sc_hd__a22o_1
X_31324_ _27701_/X _35881_/Q _31324_/S VGND VGND VPWR VPWR _31325_/A sky130_fd_sc_hd__mux2_1
X_35092_ _35221_/CLK _35092_/D VGND VGND VPWR VPWR _35092_/Q sky130_fd_sc_hd__dfxtp_1
X_16258_ _17799_/A VGND VGND VPWR VPWR _16258_/X sky130_fd_sc_hd__buf_6
XFILLER_220_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput203 _36236_/Q VGND VGND VPWR VPWR D2[54] sky130_fd_sc_hd__buf_2
X_31255_ _27797_/X _35848_/Q _31273_/S VGND VGND VPWR VPWR _31256_/A sky130_fd_sc_hd__mux2_1
X_34043_ _35448_/CLK _34043_/D VGND VGND VPWR VPWR _34043_/Q sky130_fd_sc_hd__dfxtp_1
X_16189_ _32857_/Q _32793_/Q _32729_/Q _32665_/Q _16037_/X _16039_/X VGND VGND VPWR
+ VPWR _16189_/X sky130_fd_sc_hd__mux4_1
Xoutput214 _36188_/Q VGND VGND VPWR VPWR D2[6] sky130_fd_sc_hd__buf_2
XFILLER_245_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput225 _32422_/Q VGND VGND VPWR VPWR D3[16] sky130_fd_sc_hd__buf_2
Xoutput236 _32432_/Q VGND VGND VPWR VPWR D3[26] sky130_fd_sc_hd__buf_2
X_30206_ _35351_/Q _29333_/X _30222_/S VGND VGND VPWR VPWR _30207_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput247 _32442_/Q VGND VGND VPWR VPWR D3[36] sky130_fd_sc_hd__buf_2
XFILLER_177_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput258 _32452_/Q VGND VGND VPWR VPWR D3[46] sky130_fd_sc_hd__buf_2
XFILLER_138_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31186_ _31186_/A VGND VGND VPWR VPWR _35815_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput269 _32462_/Q VGND VGND VPWR VPWR D3[56] sky130_fd_sc_hd__buf_2
XFILLER_142_886 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30137_ _30137_/A VGND VGND VPWR VPWR _35318_/D sky130_fd_sc_hd__clkbuf_1
X_19948_ _35202_/Q _35138_/Q _35074_/Q _32258_/Q _19663_/X _19664_/X VGND VGND VPWR
+ VPWR _19948_/X sky130_fd_sc_hd__mux4_1
X_35994_ _35994_/CLK _35994_/D VGND VGND VPWR VPWR _35994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34945_ _34945_/CLK _34945_/D VGND VGND VPWR VPWR _34945_/Q sky130_fd_sc_hd__dfxtp_1
X_30068_ _30200_/S VGND VGND VPWR VPWR _30087_/S sky130_fd_sc_hd__buf_6
X_19879_ _34688_/Q _34624_/Q _34560_/Q _34496_/Q _19592_/X _19593_/X VGND VGND VPWR
+ VPWR _19879_/X sky130_fd_sc_hd__mux4_1
XFILLER_210_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21910_ _32633_/Q _32569_/Q _32505_/Q _35961_/Q _21876_/X _21660_/X VGND VGND VPWR
+ VPWR _21910_/X sky130_fd_sc_hd__mux4_1
X_22890_ _22890_/A VGND VGND VPWR VPWR _32022_/D sky130_fd_sc_hd__clkbuf_1
X_34876_ _34941_/CLK _34876_/D VGND VGND VPWR VPWR _34876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33827_ _33827_/CLK _33827_/D VGND VGND VPWR VPWR _33827_/Q sky130_fd_sc_hd__dfxtp_1
X_21841_ _33911_/Q _33847_/Q _33783_/Q _36087_/Q _21624_/X _21625_/X VGND VGND VPWR
+ VPWR _21841_/X sky130_fd_sc_hd__mux4_1
XFILLER_43_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24560_ _24560_/A VGND VGND VPWR VPWR _32805_/D sky130_fd_sc_hd__clkbuf_1
X_33758_ _36207_/CLK _33758_/D VGND VGND VPWR VPWR _33758_/Q sky130_fd_sc_hd__dfxtp_1
X_21772_ _33397_/Q _33333_/Q _33269_/Q _33205_/Q _21727_/X _21728_/X VGND VGND VPWR
+ VPWR _21772_/X sky130_fd_sc_hd__mux4_1
XFILLER_212_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23511_ _32251_/Q _23411_/X _23515_/S VGND VGND VPWR VPWR _23512_/A sky130_fd_sc_hd__mux2_1
X_20723_ _20719_/X _20722_/X _20644_/X _20646_/X VGND VGND VPWR VPWR _20738_/B sky130_fd_sc_hd__o211a_1
X_32709_ _32903_/CLK _32709_/D VGND VGND VPWR VPWR _32709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24491_ _23033_/X _32773_/Q _24495_/S VGND VGND VPWR VPWR _24492_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33689_ _35610_/CLK _33689_/D VGND VGND VPWR VPWR _33689_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_68_CLK clkbuf_leaf_73_CLK/A VGND VGND VPWR VPWR _32869_/CLK sky130_fd_sc_hd__clkbuf_16
X_26230_ _26230_/A VGND VGND VPWR VPWR _33563_/D sky130_fd_sc_hd__clkbuf_1
X_23442_ _32226_/Q _23441_/X _23451_/S VGND VGND VPWR VPWR _23443_/A sky130_fd_sc_hd__mux2_1
X_35428_ _35753_/CLK _35428_/D VGND VGND VPWR VPWR _35428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20654_ _22366_/A VGND VGND VPWR VPWR _22599_/A sky130_fd_sc_hd__buf_12
XFILLER_23_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26161_ _24914_/X _33531_/Q _26165_/S VGND VGND VPWR VPWR _26162_/A sky130_fd_sc_hd__mux2_1
X_20585_ input72/X VGND VGND VPWR VPWR _20663_/A sky130_fd_sc_hd__buf_6
X_35359_ _35677_/CLK _35359_/D VGND VGND VPWR VPWR _35359_/Q sky130_fd_sc_hd__dfxtp_1
X_23373_ _32202_/Q _23305_/X _23385_/S VGND VGND VPWR VPWR _23374_/A sky130_fd_sc_hd__mux2_1
X_25112_ _24967_/X _33036_/Q _25122_/S VGND VGND VPWR VPWR _25113_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22324_ _22324_/A _22324_/B _22324_/C _22324_/D VGND VGND VPWR VPWR _22325_/A sky130_fd_sc_hd__or4_4
XFILLER_109_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26092_ _24812_/X _33498_/Q _26102_/S VGND VGND VPWR VPWR _26093_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_6_34__f_CLK clkbuf_5_17_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_34__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_30_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29920_ _35216_/Q _29509_/X _29922_/S VGND VGND VPWR VPWR _29921_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25043_ _24865_/X _33003_/Q _25059_/S VGND VGND VPWR VPWR _25044_/A sky130_fd_sc_hd__mux2_1
X_22255_ _22255_/A VGND VGND VPWR VPWR _36226_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_219_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21206_ _20953_/X _21204_/X _21205_/X _20959_/X VGND VGND VPWR VPWR _21206_/X sky130_fd_sc_hd__a22o_1
X_22186_ _22111_/X _22184_/X _22185_/X _22116_/X VGND VGND VPWR VPWR _22186_/X sky130_fd_sc_hd__a22o_1
XFILLER_156_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29851_ _35183_/Q _29407_/X _29859_/S VGND VGND VPWR VPWR _29852_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28802_ _34716_/Q _27053_/X _28808_/S VGND VGND VPWR VPWR _28803_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21137_ _21133_/X _21136_/X _21026_/X VGND VGND VPWR VPWR _21161_/A sky130_fd_sc_hd__o21ba_1
X_29782_ _29782_/A VGND VGND VPWR VPWR _35150_/D sky130_fd_sc_hd__clkbuf_1
X_26994_ _33923_/Q _23438_/X _27002_/S VGND VGND VPWR VPWR _26995_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25945_ _24994_/X _33429_/Q _25945_/S VGND VGND VPWR VPWR _25946_/A sky130_fd_sc_hd__mux2_1
X_21068_ _20747_/X _21066_/X _21067_/X _20750_/X VGND VGND VPWR VPWR _21068_/X sky130_fd_sc_hd__a22o_1
X_28733_ _28733_/A VGND VGND VPWR VPWR _34684_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20019_ _19806_/X _20015_/X _20018_/X _19809_/X VGND VGND VPWR VPWR _20019_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28664_ _28664_/A VGND VGND VPWR VPWR _34651_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25876_ _25945_/S VGND VGND VPWR VPWR _25895_/S sky130_fd_sc_hd__buf_4
XFILLER_101_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_246_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27615_ _34186_/Q _27196_/X _27629_/S VGND VGND VPWR VPWR _27616_/A sky130_fd_sc_hd__mux2_1
X_24827_ input64/X VGND VGND VPWR VPWR _24827_/X sky130_fd_sc_hd__buf_2
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28595_ _28595_/A VGND VGND VPWR VPWR _34619_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27546_ _27546_/A VGND VGND VPWR VPWR _34153_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24758_ _24758_/A VGND VGND VPWR VPWR _32899_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23709_ _22879_/X _32342_/Q _23727_/S VGND VGND VPWR VPWR _23710_/A sky130_fd_sc_hd__mux2_1
XFILLER_199_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27477_ _27477_/A VGND VGND VPWR VPWR _34120_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24689_ _24689_/A VGND VGND VPWR VPWR _32866_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_59_CLK clkbuf_leaf_61_CLK/A VGND VGND VPWR VPWR _32875_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_30_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _17936_/A VGND VGND VPWR VPWR _17230_/X sky130_fd_sc_hd__buf_6
XFILLER_187_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26428_ _33657_/Q _23405_/X _26436_/S VGND VGND VPWR VPWR _26429_/A sky130_fd_sc_hd__mux2_1
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29216_ _34912_/Q _27065_/X _29234_/S VGND VGND VPWR VPWR _29217_/A sky130_fd_sc_hd__mux2_1
XFILLER_187_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29147_ _29147_/A VGND VGND VPWR VPWR _34879_/D sky130_fd_sc_hd__clkbuf_1
X_17161_ _17161_/A VGND VGND VPWR VPWR _17161_/X sky130_fd_sc_hd__buf_4
X_26359_ _33624_/Q _23237_/X _26373_/S VGND VGND VPWR VPWR _26360_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16112_ _17850_/A VGND VGND VPWR VPWR _16112_/X sky130_fd_sc_hd__buf_6
X_29078_ _34847_/Q _27062_/X _29078_/S VGND VGND VPWR VPWR _29079_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17092_ _33651_/Q _33587_/Q _33523_/Q _33459_/Q _16847_/X _16848_/X VGND VGND VPWR
+ VPWR _17092_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16043_ input69/X VGND VGND VPWR VPWR _17846_/A sky130_fd_sc_hd__buf_6
XFILLER_129_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28029_ _34351_/Q _27112_/X _28037_/S VGND VGND VPWR VPWR _28030_/A sky130_fd_sc_hd__mux2_1
X_31040_ _31040_/A VGND VGND VPWR VPWR _35746_/D sky130_fd_sc_hd__clkbuf_1
X_19802_ _33086_/Q _32062_/Q _35838_/Q _35774_/Q _19731_/X _19732_/X VGND VGND VPWR
+ VPWR _19802_/X sky130_fd_sc_hd__mux4_1
XFILLER_170_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17994_ _35468_/Q _35404_/Q _35340_/Q _35276_/Q _17960_/X _17961_/X VGND VGND VPWR
+ VPWR _17994_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19733_ _33084_/Q _32060_/Q _35836_/Q _35772_/Q _19731_/X _19732_/X VGND VGND VPWR
+ VPWR _19733_/X sky130_fd_sc_hd__mux4_1
X_16945_ _34926_/Q _34862_/Q _34798_/Q _34734_/Q _16807_/X _16808_/X VGND VGND VPWR
+ VPWR _16945_/X sky130_fd_sc_hd__mux4_1
X_32991_ _35807_/CLK _32991_/D VGND VGND VPWR VPWR _32991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34730_ _35692_/CLK _34730_/D VGND VGND VPWR VPWR _34730_/Q sky130_fd_sc_hd__dfxtp_1
X_31942_ _23475_/X _36174_/Q _31948_/S VGND VGND VPWR VPWR _31943_/A sky130_fd_sc_hd__mux2_1
X_19664_ _20017_/A VGND VGND VPWR VPWR _19664_/X sky130_fd_sc_hd__buf_6
XFILLER_225_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16876_ _17716_/A VGND VGND VPWR VPWR _16876_/X sky130_fd_sc_hd__buf_4
XFILLER_64_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18615_ _34141_/Q _34077_/Q _34013_/Q _33949_/Q _18309_/X _18311_/X VGND VGND VPWR
+ VPWR _18615_/X sky130_fd_sc_hd__mux4_1
XFILLER_65_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34661_ _34913_/CLK _34661_/D VGND VGND VPWR VPWR _34661_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19595_ _35192_/Q _35128_/Q _35064_/Q _32248_/Q _19310_/X _19311_/X VGND VGND VPWR
+ VPWR _19595_/X sky130_fd_sc_hd__mux4_1
X_31873_ _23302_/X _36141_/Q _31885_/S VGND VGND VPWR VPWR _31874_/A sky130_fd_sc_hd__mux2_1
XFILLER_206_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33612_ _34188_/CLK _33612_/D VGND VGND VPWR VPWR _33612_/Q sky130_fd_sc_hd__dfxtp_1
X_18546_ _18440_/X _18544_/X _18545_/X _18445_/X VGND VGND VPWR VPWR _18546_/X sky130_fd_sc_hd__a22o_1
XFILLER_46_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30824_ _30824_/A VGND VGND VPWR VPWR _35644_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_209_1323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34592_ _34594_/CLK _34592_/D VGND VGND VPWR VPWR _34592_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33543_ _34185_/CLK _33543_/D VGND VGND VPWR VPWR _33543_/Q sky130_fd_sc_hd__dfxtp_1
X_18477_ _18477_/A VGND VGND VPWR VPWR _32408_/D sky130_fd_sc_hd__clkbuf_4
X_30755_ _30755_/A VGND VGND VPWR VPWR _35611_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17428_ _35644_/Q _35004_/Q _34364_/Q _33724_/Q _17144_/X _17145_/X VGND VGND VPWR
+ VPWR _17428_/X sky130_fd_sc_hd__mux4_1
X_33474_ _34942_/CLK _33474_/D VGND VGND VPWR VPWR _33474_/Q sky130_fd_sc_hd__dfxtp_1
X_30686_ _35579_/Q _29444_/X _30690_/S VGND VGND VPWR VPWR _30687_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35213_ _35213_/CLK _35213_/D VGND VGND VPWR VPWR _35213_/Q sky130_fd_sc_hd__dfxtp_1
X_32425_ _33897_/CLK _32425_/D VGND VGND VPWR VPWR _32425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36193_ _36202_/CLK _36193_/D VGND VGND VPWR VPWR _36193_/Q sky130_fd_sc_hd__dfxtp_1
X_17359_ _17869_/A VGND VGND VPWR VPWR _17359_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_179_1422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20370_ _34191_/Q _34127_/Q _34063_/Q _33999_/Q _20099_/X _20100_/X VGND VGND VPWR
+ VPWR _20370_/X sky130_fd_sc_hd__mux4_1
X_35144_ _36169_/CLK _35144_/D VGND VGND VPWR VPWR _35144_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32356_ _32356_/CLK _32356_/D VGND VGND VPWR VPWR _32356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31307_ _31307_/A VGND VGND VPWR VPWR _35872_/D sky130_fd_sc_hd__clkbuf_1
X_19029_ _19023_/X _19028_/X _18745_/X VGND VGND VPWR VPWR _19037_/C sky130_fd_sc_hd__o21ba_1
X_35075_ _35717_/CLK _35075_/D VGND VGND VPWR VPWR _35075_/Q sky130_fd_sc_hd__dfxtp_1
X_32287_ _35870_/CLK _32287_/D VGND VGND VPWR VPWR _32287_/Q sky130_fd_sc_hd__dfxtp_1
X_22040_ _34940_/Q _34876_/Q _34812_/Q _34748_/Q _21760_/X _21761_/X VGND VGND VPWR
+ VPWR _22040_/X sky130_fd_sc_hd__mux4_1
XFILLER_161_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31238_ _27773_/X _35840_/Q _31252_/S VGND VGND VPWR VPWR _31239_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34026_ _35627_/CLK _34026_/D VGND VGND VPWR VPWR _34026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31169_ _31169_/A VGND VGND VPWR VPWR _35807_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_940 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_878 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23991_ _23991_/A VGND VGND VPWR VPWR _32538_/D sky130_fd_sc_hd__clkbuf_1
X_35977_ _35980_/CLK _35977_/D VGND VGND VPWR VPWR _35977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25730_ _25730_/A VGND VGND VPWR VPWR _33326_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_217_916 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34928_ _35439_/CLK _34928_/D VGND VGND VPWR VPWR _34928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22942_ _22942_/A VGND VGND VPWR VPWR _32039_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25661_ _24973_/X _33294_/Q _25667_/S VGND VGND VPWR VPWR _25662_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22873_ _34453_/Q _36181_/Q _34325_/Q _34261_/Q _20667_/X _20669_/X VGND VGND VPWR
+ VPWR _22873_/X sky130_fd_sc_hd__mux4_1
X_34859_ _34924_/CLK _34859_/D VGND VGND VPWR VPWR _34859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27400_ _34084_/Q _27078_/X _27410_/S VGND VGND VPWR VPWR _27401_/A sky130_fd_sc_hd__mux2_1
XFILLER_243_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24612_ _23011_/X _32830_/Q _24630_/S VGND VGND VPWR VPWR _24613_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28380_ _28380_/A _31823_/B VGND VGND VPWR VPWR _28513_/S sky130_fd_sc_hd__nand2_8
X_21824_ _21603_/X _21822_/X _21823_/X _21606_/X VGND VGND VPWR VPWR _21824_/X sky130_fd_sc_hd__a22o_1
XFILLER_55_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25592_ _24871_/X _33261_/Q _25604_/S VGND VGND VPWR VPWR _25593_/A sky130_fd_sc_hd__mux2_1
XFILLER_231_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27331_ _27331_/A VGND VGND VPWR VPWR _34051_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24543_ _24543_/A VGND VGND VPWR VPWR _32797_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21755_ _35188_/Q _35124_/Q _35060_/Q _32231_/Q _21610_/X _21611_/X VGND VGND VPWR
+ VPWR _21755_/X sky130_fd_sc_hd__mux4_1
XFILLER_245_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20706_ _20706_/A _20706_/B _20706_/C _20706_/D VGND VGND VPWR VPWR _20707_/A sky130_fd_sc_hd__or4_2
X_27262_ _27262_/A VGND VGND VPWR VPWR _34018_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24474_ _23008_/X _32765_/Q _24474_/S VGND VGND VPWR VPWR _24475_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21686_ _34418_/Q _36146_/Q _34290_/Q _34226_/Q _21476_/X _21477_/X VGND VGND VPWR
+ VPWR _21686_/X sky130_fd_sc_hd__mux4_1
XFILLER_123_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29001_ _29001_/A VGND VGND VPWR VPWR _34810_/D sky130_fd_sc_hd__clkbuf_1
X_26213_ _24991_/X _33556_/Q _26215_/S VGND VGND VPWR VPWR _26214_/A sky130_fd_sc_hd__mux2_1
X_23425_ _23425_/A VGND VGND VPWR VPWR _32220_/D sky130_fd_sc_hd__clkbuf_1
X_20637_ _22433_/A VGND VGND VPWR VPWR _20637_/X sky130_fd_sc_hd__clkbuf_8
X_27193_ input47/X VGND VGND VPWR VPWR _27193_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_32_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26144_ _24889_/X _33523_/Q _26144_/S VGND VGND VPWR VPWR _26145_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23356_ _23356_/A VGND VGND VPWR VPWR _32194_/D sky130_fd_sc_hd__clkbuf_1
X_20568_ _18301_/X _20566_/X _20567_/X _18307_/X VGND VGND VPWR VPWR _20568_/X sky130_fd_sc_hd__a22o_1
XFILLER_180_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22307_ _22462_/A VGND VGND VPWR VPWR _22307_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_165_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26075_ _26075_/A VGND VGND VPWR VPWR _33490_/D sky130_fd_sc_hd__clkbuf_1
X_23287_ _32168_/Q _23286_/X _23290_/S VGND VGND VPWR VPWR _23288_/A sky130_fd_sc_hd__mux2_1
X_20499_ _32147_/Q _32339_/Q _32403_/Q _35923_/Q _20286_/X _19311_/A VGND VGND VPWR
+ VPWR _20499_/X sky130_fd_sc_hd__mux4_1
X_29903_ _29930_/S VGND VGND VPWR VPWR _29922_/S sky130_fd_sc_hd__buf_4
X_25026_ _24840_/X _32995_/Q _25038_/S VGND VGND VPWR VPWR _25027_/A sky130_fd_sc_hd__mux2_1
X_22238_ _35714_/Q _32224_/Q _35586_/Q _35522_/Q _21917_/X _21918_/X VGND VGND VPWR
+ VPWR _22238_/X sky130_fd_sc_hd__mux4_1
XFILLER_105_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29834_ _35175_/Q _29382_/X _29838_/S VGND VGND VPWR VPWR _29835_/A sky130_fd_sc_hd__mux2_1
XTAP_6944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22169_ _32896_/Q _32832_/Q _32768_/Q _32704_/Q _21946_/X _21947_/X VGND VGND VPWR
+ VPWR _22169_/X sky130_fd_sc_hd__mux4_1
XFILLER_65_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29765_ _29765_/A VGND VGND VPWR VPWR _35142_/D sky130_fd_sc_hd__clkbuf_1
X_26977_ _33915_/Q _23411_/X _26981_/S VGND VGND VPWR VPWR _26978_/A sky130_fd_sc_hd__mux2_1
XTAP_6999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28716_ _34676_/Q _27127_/X _28734_/S VGND VGND VPWR VPWR _28717_/A sky130_fd_sc_hd__mux2_1
X_16730_ _34664_/Q _34600_/Q _34536_/Q _34472_/Q _16586_/X _16587_/X VGND VGND VPWR
+ VPWR _16730_/X sky130_fd_sc_hd__mux4_1
X_25928_ _25928_/A VGND VGND VPWR VPWR _33420_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29696_ _29696_/A VGND VGND VPWR VPWR _35109_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_235_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16661_ _34406_/Q _36134_/Q _34278_/Q _34214_/Q _16523_/X _16524_/X VGND VGND VPWR
+ VPWR _16661_/X sky130_fd_sc_hd__mux4_1
X_28647_ _28647_/A VGND VGND VPWR VPWR _34644_/D sky130_fd_sc_hd__clkbuf_1
X_25859_ _25859_/A VGND VGND VPWR VPWR _33387_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18400_ _20077_/A VGND VGND VPWR VPWR _19463_/A sky130_fd_sc_hd__buf_12
XFILLER_210_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16592_ _34916_/Q _34852_/Q _34788_/Q _34724_/Q _16454_/X _16455_/X VGND VGND VPWR
+ VPWR _16592_/X sky130_fd_sc_hd__mux4_1
X_19380_ _33074_/Q _32050_/Q _35826_/Q _35762_/Q _19378_/X _19379_/X VGND VGND VPWR
+ VPWR _19380_/X sky130_fd_sc_hd__mux4_1
XFILLER_15_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28578_ _28578_/A VGND VGND VPWR VPWR _34611_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_234_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18331_ _18361_/A VGND VGND VPWR VPWR _20286_/A sky130_fd_sc_hd__buf_6
XFILLER_61_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27529_ _34145_/Q _27069_/X _27545_/S VGND VGND VPWR VPWR _27530_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18262_ _18258_/X _18261_/X _17846_/A _17847_/A VGND VGND VPWR VPWR _18277_/B sky130_fd_sc_hd__o211a_1
X_30540_ _30540_/A VGND VGND VPWR VPWR _35509_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17213_ _33142_/Q _36022_/Q _33014_/Q _32950_/Q _17062_/X _17063_/X VGND VGND VPWR
+ VPWR _17213_/X sky130_fd_sc_hd__mux4_1
X_18193_ _33939_/Q _33875_/Q _33811_/Q _36115_/Q _16062_/X _16064_/X VGND VGND VPWR
+ VPWR _18193_/X sky130_fd_sc_hd__mux4_1
XFILLER_202_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30471_ _30471_/A VGND VGND VPWR VPWR _35477_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32210_ _35701_/CLK _32210_/D VGND VGND VPWR VPWR _32210_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17144_ _17998_/A VGND VGND VPWR VPWR _17144_/X sky130_fd_sc_hd__buf_6
X_33190_ _33697_/CLK _33190_/D VGND VGND VPWR VPWR _33190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32141_ _35980_/CLK _32141_/D VGND VGND VPWR VPWR _32141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17075_ _35634_/Q _34994_/Q _34354_/Q _33714_/Q _16791_/X _16792_/X VGND VGND VPWR
+ VPWR _17075_/X sky130_fd_sc_hd__mux4_1
XFILLER_226_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16026_ _33110_/Q _35990_/Q _32982_/Q _32918_/Q _16024_/X _16025_/X VGND VGND VPWR
+ VPWR _16026_/X sky130_fd_sc_hd__mux4_1
X_32072_ _33160_/CLK _32072_/D VGND VGND VPWR VPWR _32072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31023_ _31023_/A VGND VGND VPWR VPWR _35738_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35900_ _35964_/CLK _35900_/D VGND VGND VPWR VPWR _35900_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35831_ _36151_/CLK _35831_/D VGND VGND VPWR VPWR _35831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17977_ _17905_/X _17975_/X _17976_/X _17910_/X VGND VGND VPWR VPWR _17977_/X sky130_fd_sc_hd__a22o_1
XFILLER_85_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19716_ _20074_/A VGND VGND VPWR VPWR _19716_/X sky130_fd_sc_hd__buf_4
X_35762_ _36146_/CLK _35762_/D VGND VGND VPWR VPWR _35762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16928_ _32110_/Q _32302_/Q _32366_/Q _35886_/Q _16927_/X _16715_/X VGND VGND VPWR
+ VPWR _16928_/X sky130_fd_sc_hd__mux4_1
X_32974_ _35853_/CLK _32974_/D VGND VGND VPWR VPWR _32974_/Q sky130_fd_sc_hd__dfxtp_1
X_34713_ _34911_/CLK _34713_/D VGND VGND VPWR VPWR _34713_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31925_ _23447_/X _36166_/Q _31927_/S VGND VGND VPWR VPWR _31926_/A sky130_fd_sc_hd__mux2_1
X_19647_ _20134_/A VGND VGND VPWR VPWR _19647_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_1_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35693_ _35693_/CLK _35693_/D VGND VGND VPWR VPWR _35693_/Q sky130_fd_sc_hd__dfxtp_1
X_16859_ _32620_/Q _32556_/Q _32492_/Q _35948_/Q _16570_/X _16707_/X VGND VGND VPWR
+ VPWR _16859_/X sky130_fd_sc_hd__mux4_1
XFILLER_92_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34644_ _34708_/CLK _34644_/D VGND VGND VPWR VPWR _34644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31856_ _23277_/X _36133_/Q _31864_/S VGND VGND VPWR VPWR _31857_/A sky130_fd_sc_hd__mux2_1
X_19578_ _33144_/Q _36024_/Q _33016_/Q _32952_/Q _19362_/X _19363_/X VGND VGND VPWR
+ VPWR _19578_/X sky130_fd_sc_hd__mux4_1
XFILLER_168_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18529_ _35418_/Q _35354_/Q _35290_/Q _35226_/Q _18495_/X _18496_/X VGND VGND VPWR
+ VPWR _18529_/X sky130_fd_sc_hd__mux4_1
X_30807_ _35636_/Q input24/X _30825_/S VGND VGND VPWR VPWR _30808_/A sky130_fd_sc_hd__mux2_1
XFILLER_244_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34575_ _34705_/CLK _34575_/D VGND VGND VPWR VPWR _34575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31787_ _31787_/A VGND VGND VPWR VPWR _36100_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33526_ _34166_/CLK _33526_/D VGND VGND VPWR VPWR _33526_/Q sky130_fd_sc_hd__dfxtp_1
X_21540_ _22599_/A VGND VGND VPWR VPWR _21540_/X sky130_fd_sc_hd__clkbuf_4
X_30738_ _35604_/Q _29521_/X _30740_/S VGND VGND VPWR VPWR _30739_/A sky130_fd_sc_hd__mux2_1
XFILLER_244_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36245_ _36245_/CLK _36245_/D VGND VGND VPWR VPWR _36245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33457_ _33904_/CLK _33457_/D VGND VGND VPWR VPWR _33457_/Q sky130_fd_sc_hd__dfxtp_1
X_21471_ _21250_/X _21469_/X _21470_/X _21253_/X VGND VGND VPWR VPWR _21471_/X sky130_fd_sc_hd__a22o_1
XFILLER_194_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30669_ _35571_/Q _29419_/X _30669_/S VGND VGND VPWR VPWR _30670_/A sky130_fd_sc_hd__mux2_1
X_23210_ _23210_/A VGND VGND VPWR VPWR _32142_/D sky130_fd_sc_hd__clkbuf_1
X_20422_ _20159_/X _20420_/X _20421_/X _20162_/X VGND VGND VPWR VPWR _20422_/X sky130_fd_sc_hd__a22o_1
XFILLER_147_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32408_ _34151_/CLK _32408_/D VGND VGND VPWR VPWR _32408_/Q sky130_fd_sc_hd__dfxtp_1
X_36176_ _36176_/CLK _36176_/D VGND VGND VPWR VPWR _36176_/Q sky130_fd_sc_hd__dfxtp_1
X_24190_ _24190_/A VGND VGND VPWR VPWR _32631_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33388_ _36076_/CLK _33388_/D VGND VGND VPWR VPWR _33388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35127_ _35191_/CLK _35127_/D VGND VGND VPWR VPWR _35127_/Q sky130_fd_sc_hd__dfxtp_1
X_23141_ _23141_/A VGND VGND VPWR VPWR _32109_/D sky130_fd_sc_hd__clkbuf_1
X_20353_ _35726_/Q _32237_/Q _35598_/Q _35534_/Q _18293_/X _18295_/X VGND VGND VPWR
+ VPWR _20353_/X sky130_fd_sc_hd__mux4_1
X_32339_ _35986_/CLK _32339_/D VGND VGND VPWR VPWR _32339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23072_ _23072_/A VGND VGND VPWR VPWR _32081_/D sky130_fd_sc_hd__clkbuf_1
X_20284_ _33164_/Q _36044_/Q _33036_/Q _32972_/Q _20068_/X _20069_/X VGND VGND VPWR
+ VPWR _20284_/X sky130_fd_sc_hd__mux4_1
X_35058_ _35828_/CLK _35058_/D VGND VGND VPWR VPWR _35058_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_11_0_CLK clkbuf_5_9_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_11_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XTAP_6218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34009_ _34009_/CLK _34009_/D VGND VGND VPWR VPWR _34009_/Q sky130_fd_sc_hd__dfxtp_1
X_26900_ _33878_/Q _23225_/X _26918_/S VGND VGND VPWR VPWR _26901_/A sky130_fd_sc_hd__mux2_1
X_22023_ _32892_/Q _32828_/Q _32764_/Q _32700_/Q _21946_/X _21947_/X VGND VGND VPWR
+ VPWR _22023_/X sky130_fd_sc_hd__mux4_1
XTAP_6229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27880_ _27880_/A VGND VGND VPWR VPWR _34280_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26831_ _26831_/A VGND VGND VPWR VPWR _33845_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26762_ _26762_/A VGND VGND VPWR VPWR _33813_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29550_ _35040_/Q _29360_/X _29568_/S VGND VGND VPWR VPWR _29551_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_5_26_0_CLK clkbuf_2_3_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_26_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XTAP_4849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23974_ _23974_/A VGND VGND VPWR VPWR _32531_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28501_ _27819_/X _34575_/Q _28505_/S VGND VGND VPWR VPWR _28502_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25713_ _25713_/A VGND VGND VPWR VPWR _33318_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22925_ input4/X VGND VGND VPWR VPWR _22925_/X sky130_fd_sc_hd__clkbuf_4
X_29481_ input44/X VGND VGND VPWR VPWR _29481_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_21_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26693_ _33780_/Q _23387_/X _26711_/S VGND VGND VPWR VPWR _26694_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25644_ _24948_/X _33286_/Q _25646_/S VGND VGND VPWR VPWR _25645_/A sky130_fd_sc_hd__mux2_1
X_28432_ _27717_/X _34542_/Q _28442_/S VGND VGND VPWR VPWR _28433_/A sky130_fd_sc_hd__mux2_1
XFILLER_189_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22856_ _32661_/Q _32597_/Q _32533_/Q _35989_/Q _22582_/X _21477_/A VGND VGND VPWR
+ VPWR _22856_/X sky130_fd_sc_hd__mux4_1
XFILLER_244_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28363_ _28363_/A VGND VGND VPWR VPWR _34509_/D sky130_fd_sc_hd__clkbuf_1
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21807_ _33398_/Q _33334_/Q _33270_/Q _33206_/Q _21727_/X _21728_/X VGND VGND VPWR
+ VPWR _21807_/X sky130_fd_sc_hd__mux4_1
XFILLER_73_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25575_ _24846_/X _33253_/Q _25583_/S VGND VGND VPWR VPWR _25576_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22787_ _22787_/A _22787_/B _22787_/C _22787_/D VGND VGND VPWR VPWR _22788_/A sky130_fd_sc_hd__or4_4
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27314_ _27314_/A VGND VGND VPWR VPWR _34043_/D sky130_fd_sc_hd__clkbuf_1
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24526_ _31823_/A _31553_/B VGND VGND VPWR VPWR _24659_/S sky130_fd_sc_hd__nand2_8
XFILLER_213_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28294_ _28294_/A VGND VGND VPWR VPWR _34476_/D sky130_fd_sc_hd__clkbuf_1
X_21738_ _32884_/Q _32820_/Q _32756_/Q _32692_/Q _21593_/X _21594_/X VGND VGND VPWR
+ VPWR _21738_/X sky130_fd_sc_hd__mux4_1
XFILLER_213_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27245_ _27245_/A VGND VGND VPWR VPWR _34010_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24457_ _24457_/A VGND VGND VPWR VPWR _32756_/D sky130_fd_sc_hd__clkbuf_1
X_21669_ _32114_/Q _32306_/Q _32370_/Q _35890_/Q _21527_/X _21668_/X VGND VGND VPWR
+ VPWR _21669_/X sky130_fd_sc_hd__mux4_1
XFILLER_201_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23408_ input30/X VGND VGND VPWR VPWR _23408_/X sky130_fd_sc_hd__buf_4
X_27176_ _27176_/A VGND VGND VPWR VPWR _33987_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24388_ _24388_/A VGND VGND VPWR VPWR _32724_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26127_ _26127_/A VGND VGND VPWR VPWR _33514_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23339_ _23339_/A VGND VGND VPWR VPWR _32186_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26058_ _24961_/X _33482_/Q _26072_/S VGND VGND VPWR VPWR _26059_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17900_ _34953_/Q _34889_/Q _34825_/Q _34761_/Q _17866_/X _17867_/X VGND VGND VPWR
+ VPWR _17900_/X sky130_fd_sc_hd__mux4_1
XFILLER_180_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25009_ _24815_/X _32987_/Q _25017_/S VGND VGND VPWR VPWR _25010_/A sky130_fd_sc_hd__mux2_1
X_18880_ _35620_/Q _34980_/Q _34340_/Q _33700_/Q _18738_/X _18739_/X VGND VGND VPWR
+ VPWR _18880_/X sky130_fd_sc_hd__mux4_1
XTAP_6730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17831_ _34184_/Q _34120_/Q _34056_/Q _33992_/Q _17799_/X _17800_/X VGND VGND VPWR
+ VPWR _17831_/X sky130_fd_sc_hd__mux4_1
XFILLER_239_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29817_ _35167_/Q _29357_/X _29817_/S VGND VGND VPWR VPWR _29818_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17762_ _33926_/Q _33862_/Q _33798_/Q _36102_/Q _17730_/X _17731_/X VGND VGND VPWR
+ VPWR _17762_/X sky130_fd_sc_hd__mux4_1
X_29748_ _35134_/Q _29453_/X _29766_/S VGND VGND VPWR VPWR _29749_/A sky130_fd_sc_hd__mux2_1
XFILLER_187_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_1244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19501_ _20207_/A VGND VGND VPWR VPWR _19501_/X sky130_fd_sc_hd__buf_4
XFILLER_169_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_762 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16713_ _16706_/X _16708_/X _16711_/X _16712_/X VGND VGND VPWR VPWR _16713_/X sky130_fd_sc_hd__a22o_1
X_29679_ _29679_/A VGND VGND VPWR VPWR _35101_/D sky130_fd_sc_hd__clkbuf_1
X_17693_ _17559_/X _17691_/X _17692_/X _17562_/X VGND VGND VPWR VPWR _17693_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_290_CLK clkbuf_6_56__f_CLK/X VGND VGND VPWR VPWR _36033_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_34_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19432_ _20138_/A VGND VGND VPWR VPWR _19432_/X sky130_fd_sc_hd__buf_2
X_31710_ _31821_/S VGND VGND VPWR VPWR _31729_/S sky130_fd_sc_hd__buf_4
X_16644_ _16638_/X _16643_/X _16434_/X _16435_/X VGND VGND VPWR VPWR _16665_/B sky130_fd_sc_hd__o211a_1
X_32690_ _32818_/CLK _32690_/D VGND VGND VPWR VPWR _32690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_216_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31641_ _27770_/X _36031_/Q _31657_/S VGND VGND VPWR VPWR _31642_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19363_ _20074_/A VGND VGND VPWR VPWR _19363_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_245_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16575_ _32100_/Q _32292_/Q _32356_/Q _35876_/Q _16574_/X _16362_/X VGND VGND VPWR
+ VPWR _16575_/X sky130_fd_sc_hd__mux4_1
XFILLER_206_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18314_ input81/X input82/X VGND VGND VPWR VPWR _20138_/A sky130_fd_sc_hd__or2b_4
XFILLER_31_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34360_ _35704_/CLK _34360_/D VGND VGND VPWR VPWR _34360_/Q sky130_fd_sc_hd__dfxtp_1
X_31572_ _31572_/A VGND VGND VPWR VPWR _35998_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19294_ _20134_/A VGND VGND VPWR VPWR _19294_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_826 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33311_ _35551_/CLK _33311_/D VGND VGND VPWR VPWR _33311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18245_ _16060_/X _18243_/X _18244_/X _16072_/X VGND VGND VPWR VPWR _18245_/X sky130_fd_sc_hd__a22o_1
X_30523_ _30523_/A VGND VGND VPWR VPWR _35501_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34291_ _36144_/CLK _34291_/D VGND VGND VPWR VPWR _34291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36030_ _36030_/CLK _36030_/D VGND VGND VPWR VPWR _36030_/Q sky130_fd_sc_hd__dfxtp_1
X_30454_ _35469_/Q _29500_/X _30462_/S VGND VGND VPWR VPWR _30455_/A sky130_fd_sc_hd__mux2_1
X_33242_ _33818_/CLK _33242_/D VGND VGND VPWR VPWR _33242_/Q sky130_fd_sc_hd__dfxtp_1
X_18176_ _35474_/Q _35410_/Q _35346_/Q _35282_/Q _17960_/X _17961_/X VGND VGND VPWR
+ VPWR _18176_/X sky130_fd_sc_hd__mux4_1
XFILLER_237_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17127_ _17833_/A VGND VGND VPWR VPWR _17127_/X sky130_fd_sc_hd__buf_4
XFILLER_50_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33173_ _36052_/CLK _33173_/D VGND VGND VPWR VPWR _33173_/Q sky130_fd_sc_hd__dfxtp_1
X_30385_ _35436_/Q _29398_/X _30399_/S VGND VGND VPWR VPWR _30386_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17058_ _17054_/X _17057_/X _16779_/X VGND VGND VPWR VPWR _17090_/A sky130_fd_sc_hd__o21ba_1
X_32124_ _35964_/CLK _32124_/D VGND VGND VPWR VPWR _32124_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16009_ _17960_/A VGND VGND VPWR VPWR _16009_/X sky130_fd_sc_hd__buf_6
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32055_ _35830_/CLK _32055_/D VGND VGND VPWR VPWR _32055_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31006_ _35731_/Q input58/X _31010_/S VGND VGND VPWR VPWR _31007_/A sky130_fd_sc_hd__mux2_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35814_ _35814_/CLK _35814_/D VGND VGND VPWR VPWR _35814_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35745_ _35810_/CLK _35745_/D VGND VGND VPWR VPWR _35745_/Q sky130_fd_sc_hd__dfxtp_1
X_20971_ _35422_/Q _35358_/Q _35294_/Q _35230_/Q _20795_/X _20796_/X VGND VGND VPWR
+ VPWR _20971_/X sky130_fd_sc_hd__mux4_1
X_32957_ _36029_/CLK _32957_/D VGND VGND VPWR VPWR _32957_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_281_CLK clkbuf_6_59__f_CLK/X VGND VGND VPWR VPWR _36096_/CLK sky130_fd_sc_hd__clkbuf_16
X_22710_ _32912_/Q _32848_/Q _32784_/Q _32720_/Q _20584_/X _20587_/X VGND VGND VPWR
+ VPWR _22710_/X sky130_fd_sc_hd__mux4_1
XFILLER_241_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31908_ _31956_/S VGND VGND VPWR VPWR _31927_/S sky130_fd_sc_hd__buf_4
XFILLER_199_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35676_ _35804_/CLK _35676_/D VGND VGND VPWR VPWR _35676_/Q sky130_fd_sc_hd__dfxtp_1
X_23690_ _23064_/X _32335_/Q _23694_/S VGND VGND VPWR VPWR _23691_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32888_ _32891_/CLK _32888_/D VGND VGND VPWR VPWR _32888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22641_ _22505_/X _22639_/X _22640_/X _22510_/X VGND VGND VPWR VPWR _22641_/X sky130_fd_sc_hd__a22o_1
X_34627_ _34690_/CLK _34627_/D VGND VGND VPWR VPWR _34627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31839_ _23252_/X _36125_/Q _31843_/S VGND VGND VPWR VPWR _31840_/A sky130_fd_sc_hd__mux2_1
XFILLER_179_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25360_ _33152_/Q _23429_/X _25374_/S VGND VGND VPWR VPWR _25361_/A sky130_fd_sc_hd__mux2_1
X_22572_ _22568_/X _22571_/X _22471_/X VGND VGND VPWR VPWR _22573_/D sky130_fd_sc_hd__o21ba_1
X_34558_ _35071_/CLK _34558_/D VGND VGND VPWR VPWR _34558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24311_ _24311_/A VGND VGND VPWR VPWR _32687_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33509_ _34146_/CLK _33509_/D VGND VGND VPWR VPWR _33509_/Q sky130_fd_sc_hd__dfxtp_1
X_21523_ _22582_/A VGND VGND VPWR VPWR _21523_/X sky130_fd_sc_hd__buf_6
XFILLER_194_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25291_ _25291_/A VGND VGND VPWR VPWR _33119_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34489_ _35193_/CLK _34489_/D VGND VGND VPWR VPWR _34489_/Q sky130_fd_sc_hd__dfxtp_1
X_27030_ _27030_/A VGND VGND VPWR VPWR _33940_/D sky130_fd_sc_hd__clkbuf_1
X_36228_ _36229_/CLK _36228_/D VGND VGND VPWR VPWR _36228_/Q sky130_fd_sc_hd__dfxtp_1
X_24242_ _24242_/A VGND VGND VPWR VPWR _32656_/D sky130_fd_sc_hd__clkbuf_1
X_21454_ _33388_/Q _33324_/Q _33260_/Q _33196_/Q _21374_/X _21375_/X VGND VGND VPWR
+ VPWR _21454_/X sky130_fd_sc_hd__mux4_1
XFILLER_108_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20405_ _20401_/X _20404_/X _20138_/X VGND VGND VPWR VPWR _20427_/A sky130_fd_sc_hd__o21ba_2
XFILLER_135_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36159_ _36159_/CLK _36159_/D VGND VGND VPWR VPWR _36159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24173_ _24173_/A VGND VGND VPWR VPWR _32623_/D sky130_fd_sc_hd__clkbuf_1
X_21385_ _32874_/Q _32810_/Q _32746_/Q _32682_/Q _21240_/X _21241_/X VGND VGND VPWR
+ VPWR _21385_/X sky130_fd_sc_hd__mux4_1
XFILLER_208_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23124_ _23124_/A VGND VGND VPWR VPWR _32101_/D sky130_fd_sc_hd__clkbuf_1
X_20336_ _20332_/X _20335_/X _20171_/X VGND VGND VPWR VPWR _20337_/D sky130_fd_sc_hd__o21ba_1
X_28981_ _34801_/Q _27118_/X _28985_/S VGND VGND VPWR VPWR _28982_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27932_ _27776_/X _34305_/Q _27944_/S VGND VGND VPWR VPWR _27933_/A sky130_fd_sc_hd__mux2_1
X_23055_ input50/X VGND VGND VPWR VPWR _23055_/X sky130_fd_sc_hd__buf_2
XTAP_6026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20267_ _35211_/Q _35147_/Q _35083_/Q _32267_/Q _20016_/X _20017_/X VGND VGND VPWR
+ VPWR _20267_/X sky130_fd_sc_hd__mux4_1
XFILLER_157_1380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22006_ _34172_/Q _34108_/Q _34044_/Q _33980_/Q _21693_/X _21694_/X VGND VGND VPWR
+ VPWR _22006_/X sky130_fd_sc_hd__mux4_1
XTAP_6059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20198_ _20159_/X _20196_/X _20197_/X _20162_/X VGND VGND VPWR VPWR _20198_/X sky130_fd_sc_hd__a22o_1
XTAP_5325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27863_ _27673_/X _34272_/Q _27881_/S VGND VGND VPWR VPWR _27864_/A sky130_fd_sc_hd__mux2_1
XTAP_5336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29602_ _35065_/Q _29438_/X _29610_/S VGND VGND VPWR VPWR _29603_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26814_ _26814_/A VGND VGND VPWR VPWR _33837_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27794_ input44/X VGND VGND VPWR VPWR _27794_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29533_ _35032_/Q _29336_/X _29547_/S VGND VGND VPWR VPWR _29534_/A sky130_fd_sc_hd__mux2_1
XTAP_4668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26745_ _33805_/Q _23472_/X _26753_/S VGND VGND VPWR VPWR _26746_/A sky130_fd_sc_hd__mux2_1
X_23957_ _23052_/X _32523_/Q _23969_/S VGND VGND VPWR VPWR _23958_/A sky130_fd_sc_hd__mux2_1
XTAP_3934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_272_CLK clkbuf_6_57__f_CLK/X VGND VGND VPWR VPWR _35715_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22908_ _22908_/A VGND VGND VPWR VPWR _32028_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29464_ _35009_/Q _29463_/X _29482_/S VGND VGND VPWR VPWR _29465_/A sky130_fd_sc_hd__mux2_1
XTAP_3978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26676_ _33772_/Q _23299_/X _26690_/S VGND VGND VPWR VPWR _26677_/A sky130_fd_sc_hd__mux2_1
XTAP_3989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23888_ _22949_/X _32490_/Q _23906_/S VGND VGND VPWR VPWR _23889_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28415_ _27692_/X _34534_/Q _28421_/S VGND VGND VPWR VPWR _28416_/A sky130_fd_sc_hd__mux2_1
X_22839_ _22835_/X _22838_/X _22457_/A VGND VGND VPWR VPWR _22847_/C sky130_fd_sc_hd__o21ba_1
X_25627_ _25675_/S VGND VGND VPWR VPWR _25646_/S sky130_fd_sc_hd__buf_4
XFILLER_16_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29395_ input14/X VGND VGND VPWR VPWR _29395_/X sky130_fd_sc_hd__buf_2
XFILLER_112_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16360_ _16353_/X _16355_/X _16358_/X _16359_/X VGND VGND VPWR VPWR _16360_/X sky130_fd_sc_hd__a22o_1
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28346_ _28346_/A VGND VGND VPWR VPWR _34501_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25558_ _24821_/X _33245_/Q _25562_/S VGND VGND VPWR VPWR _25559_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24509_ _24509_/A VGND VGND VPWR VPWR _32781_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16291_ _16285_/X _16290_/X _16044_/X _16046_/X VGND VGND VPWR VPWR _16312_/B sky130_fd_sc_hd__o211a_1
X_28277_ _28277_/A VGND VGND VPWR VPWR _34468_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25489_ _25489_/A VGND VGND VPWR VPWR _33212_/D sky130_fd_sc_hd__clkbuf_1
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_240_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18030_ _34701_/Q _34637_/Q _34573_/Q _34509_/Q _17998_/X _17999_/X VGND VGND VPWR
+ VPWR _18030_/X sky130_fd_sc_hd__mux4_1
X_27228_ _27228_/A VGND VGND VPWR VPWR _34004_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_818 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27159_ _27230_/S VGND VGND VPWR VPWR _27187_/S sky130_fd_sc_hd__buf_6
XFILLER_165_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30170_ _30170_/A VGND VGND VPWR VPWR _35334_/D sky130_fd_sc_hd__clkbuf_1
X_19981_ _19806_/X _19979_/X _19980_/X _19809_/X VGND VGND VPWR VPWR _19981_/X sky130_fd_sc_hd__a22o_1
XFILLER_126_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18932_ _33382_/Q _33318_/Q _33254_/Q _33190_/Q _18721_/X _18722_/X VGND VGND VPWR
+ VPWR _18932_/X sky130_fd_sc_hd__mux4_1
XFILLER_239_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18863_ _33636_/Q _33572_/Q _33508_/Q _33444_/Q _18794_/X _18795_/X VGND VGND VPWR
+ VPWR _18863_/X sky130_fd_sc_hd__mux4_1
XFILLER_79_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17814_ _35719_/Q _32229_/Q _35591_/Q _35527_/Q _17670_/X _17671_/X VGND VGND VPWR
+ VPWR _17814_/X sky130_fd_sc_hd__mux4_1
XFILLER_239_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33860_ _33924_/CLK _33860_/D VGND VGND VPWR VPWR _33860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18794_ _20206_/A VGND VGND VPWR VPWR _18794_/X sky130_fd_sc_hd__buf_6
XFILLER_227_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_902 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32811_ _32875_/CLK _32811_/D VGND VGND VPWR VPWR _32811_/Q sky130_fd_sc_hd__dfxtp_1
X_17745_ _35461_/Q _35397_/Q _35333_/Q _35269_/Q _17607_/X _17608_/X VGND VGND VPWR
+ VPWR _17745_/X sky130_fd_sc_hd__mux4_1
X_33791_ _36095_/CLK _33791_/D VGND VGND VPWR VPWR _33791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_263_CLK clkbuf_6_62__f_CLK/X VGND VGND VPWR VPWR _36101_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_63_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35530_ _35723_/CLK _35530_/D VGND VGND VPWR VPWR _35530_/Q sky130_fd_sc_hd__dfxtp_1
X_32742_ _32873_/CLK _32742_/D VGND VGND VPWR VPWR _32742_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17676_ _33091_/Q _32067_/Q _35843_/Q _35779_/Q _17431_/X _17432_/X VGND VGND VPWR
+ VPWR _17676_/X sky130_fd_sc_hd__mux4_1
XFILLER_35_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19415_ _34675_/Q _34611_/Q _34547_/Q _34483_/Q _19239_/X _19240_/X VGND VGND VPWR
+ VPWR _19415_/X sky130_fd_sc_hd__mux4_1
X_35461_ _35845_/CLK _35461_/D VGND VGND VPWR VPWR _35461_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16627_ _16627_/A _16627_/B _16627_/C _16627_/D VGND VGND VPWR VPWR _16628_/A sky130_fd_sc_hd__or4_2
X_32673_ _35875_/CLK _32673_/D VGND VGND VPWR VPWR _32673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34412_ _36142_/CLK _34412_/D VGND VGND VPWR VPWR _34412_/Q sky130_fd_sc_hd__dfxtp_1
X_19346_ _34417_/Q _36145_/Q _34289_/Q _34225_/Q _19176_/X _19177_/X VGND VGND VPWR
+ VPWR _19346_/X sky130_fd_sc_hd__mux4_1
X_31624_ _27745_/X _36023_/Q _31636_/S VGND VGND VPWR VPWR _31625_/A sky130_fd_sc_hd__mux2_1
X_35392_ _35839_/CLK _35392_/D VGND VGND VPWR VPWR _35392_/Q sky130_fd_sc_hd__dfxtp_1
X_16558_ _34915_/Q _34851_/Q _34787_/Q _34723_/Q _16454_/X _16455_/X VGND VGND VPWR
+ VPWR _16558_/X sky130_fd_sc_hd__mux4_1
XFILLER_56_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34343_ _35559_/CLK _34343_/D VGND VGND VPWR VPWR _34343_/Q sky130_fd_sc_hd__dfxtp_1
X_31555_ _27639_/X _35990_/Q _31573_/S VGND VGND VPWR VPWR _31556_/A sky130_fd_sc_hd__mux2_1
XFILLER_175_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19277_ _34927_/Q _34863_/Q _34799_/Q _34735_/Q _19107_/X _19108_/X VGND VGND VPWR
+ VPWR _19277_/X sky130_fd_sc_hd__mux4_1
XFILLER_176_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16489_ _16452_/X _16487_/X _16488_/X _16457_/X VGND VGND VPWR VPWR _16489_/X sky130_fd_sc_hd__a22o_1
XFILLER_206_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18228_ _17153_/A _18226_/X _18227_/X _17156_/A VGND VGND VPWR VPWR _18228_/X sky130_fd_sc_hd__a22o_1
X_30506_ _30506_/A VGND VGND VPWR VPWR _35493_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_248_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34274_ _36210_/CLK _34274_/D VGND VGND VPWR VPWR _34274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31486_ _31486_/A VGND VGND VPWR VPWR _35957_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36013_ _36013_/CLK _36013_/D VGND VGND VPWR VPWR _36013_/Q sky130_fd_sc_hd__dfxtp_1
X_33225_ _33420_/CLK _33225_/D VGND VGND VPWR VPWR _33225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18159_ _33682_/Q _33618_/Q _33554_/Q _33490_/Q _17906_/X _17907_/X VGND VGND VPWR
+ VPWR _18159_/X sky130_fd_sc_hd__mux4_1
X_30437_ _35461_/Q _29475_/X _30441_/S VGND VGND VPWR VPWR _30438_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33156_ _35779_/CLK _33156_/D VGND VGND VPWR VPWR _33156_/Q sky130_fd_sc_hd__dfxtp_1
X_21170_ _22582_/A VGND VGND VPWR VPWR _21170_/X sky130_fd_sc_hd__buf_6
X_30368_ _35428_/Q _29373_/X _30378_/S VGND VGND VPWR VPWR _30369_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20121_ _34695_/Q _34631_/Q _34567_/Q _34503_/Q _19945_/X _19946_/X VGND VGND VPWR
+ VPWR _20121_/X sky130_fd_sc_hd__mux4_1
X_32107_ _35949_/CLK _32107_/D VGND VGND VPWR VPWR _32107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_217_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30299_ _30299_/A VGND VGND VPWR VPWR _35395_/D sky130_fd_sc_hd__clkbuf_1
X_33087_ _35839_/CLK _33087_/D VGND VGND VPWR VPWR _33087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20052_ _34437_/Q _36165_/Q _34309_/Q _34245_/Q _19882_/X _19883_/X VGND VGND VPWR
+ VPWR _20052_/X sky130_fd_sc_hd__mux4_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32038_ _35755_/CLK _32038_/D VGND VGND VPWR VPWR _32038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_217_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24860_ _24860_/A VGND VGND VPWR VPWR _32937_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_246_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23811_ _23039_/X _32391_/Q _23811_/S VGND VGND VPWR VPWR _23812_/A sky130_fd_sc_hd__mux2_1
XFILLER_227_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24791_ _24791_/A VGND VGND VPWR VPWR _32915_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33989_ _34183_/CLK _33989_/D VGND VGND VPWR VPWR _33989_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_254_CLK clkbuf_6_63__f_CLK/X VGND VGND VPWR VPWR _34182_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_213_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26530_ _24858_/X _33705_/Q _26530_/S VGND VGND VPWR VPWR _26531_/A sky130_fd_sc_hd__mux2_1
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35728_ _35728_/CLK _35728_/D VGND VGND VPWR VPWR _35728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23742_ _22937_/X _32358_/Q _23748_/S VGND VGND VPWR VPWR _23743_/A sky130_fd_sc_hd__mux2_1
XFILLER_214_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20954_ _22366_/A VGND VGND VPWR VPWR _20954_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26461_ _26461_/A VGND VGND VPWR VPWR _33672_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35659_ _35724_/CLK _35659_/D VGND VGND VPWR VPWR _35659_/Q sky130_fd_sc_hd__dfxtp_1
X_23673_ _23039_/X _32327_/Q _23673_/S VGND VGND VPWR VPWR _23674_/A sky130_fd_sc_hd__mux2_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20885_ _20618_/X _20883_/X _20884_/X _20627_/X VGND VGND VPWR VPWR _20885_/X sky130_fd_sc_hd__a22o_1
XFILLER_42_938 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28200_ _27773_/X _34432_/Q _28214_/S VGND VGND VPWR VPWR _28201_/A sky130_fd_sc_hd__mux2_1
X_25412_ _25412_/A VGND VGND VPWR VPWR _33175_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29180_ _29180_/A VGND VGND VPWR VPWR _34895_/D sky130_fd_sc_hd__clkbuf_1
X_22624_ _35661_/Q _35021_/Q _34381_/Q _33741_/Q _22450_/X _22451_/X VGND VGND VPWR
+ VPWR _22624_/X sky130_fd_sc_hd__mux4_1
X_26392_ _33640_/Q _23286_/X _26394_/S VGND VGND VPWR VPWR _26393_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28131_ _28131_/A VGND VGND VPWR VPWR _34399_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25343_ _33144_/Q _23402_/X _25353_/S VGND VGND VPWR VPWR _25344_/A sky130_fd_sc_hd__mux2_1
X_22555_ _22373_/X _22553_/X _22554_/X _22377_/X VGND VGND VPWR VPWR _22555_/X sky130_fd_sc_hd__a22o_1
XFILLER_107_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_976 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28062_ _28062_/A VGND VGND VPWR VPWR _34366_/D sky130_fd_sc_hd__clkbuf_1
X_21506_ _21500_/X _21505_/X _21398_/X VGND VGND VPWR VPWR _21514_/C sky130_fd_sc_hd__o21ba_1
X_25274_ _33111_/Q _23234_/X _25290_/S VGND VGND VPWR VPWR _25275_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22486_ _32905_/Q _32841_/Q _32777_/Q _32713_/Q _22299_/X _22300_/X VGND VGND VPWR
+ VPWR _22486_/X sky130_fd_sc_hd__mux4_1
XFILLER_108_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27013_ _33932_/Q _23469_/X _27023_/S VGND VGND VPWR VPWR _27014_/A sky130_fd_sc_hd__mux2_1
X_24225_ _32648_/Q _23453_/X _24243_/S VGND VGND VPWR VPWR _24226_/A sky130_fd_sc_hd__mux2_1
XFILLER_181_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21437_ _34667_/Q _34603_/Q _34539_/Q _34475_/Q _21186_/X _21187_/X VGND VGND VPWR
+ VPWR _21437_/X sky130_fd_sc_hd__mux4_1
XFILLER_68_1303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24156_ _24156_/A VGND VGND VPWR VPWR _32615_/D sky130_fd_sc_hd__clkbuf_1
X_21368_ _21364_/X _21367_/X _21059_/X VGND VGND VPWR VPWR _21369_/D sky130_fd_sc_hd__o21ba_1
XFILLER_163_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23107_ _23107_/A VGND VGND VPWR VPWR _32093_/D sky130_fd_sc_hd__clkbuf_1
X_20319_ _32141_/Q _32333_/Q _32397_/Q _35917_/Q _20286_/X _20074_/X VGND VGND VPWR
+ VPWR _20319_/X sky130_fd_sc_hd__mux4_1
X_24087_ _23042_/X _32584_/Q _24105_/S VGND VGND VPWR VPWR _24088_/A sky130_fd_sc_hd__mux2_1
X_28964_ _34793_/Q _27093_/X _28964_/S VGND VGND VPWR VPWR _28965_/A sky130_fd_sc_hd__mux2_1
X_21299_ _33640_/Q _33576_/Q _33512_/Q _33448_/Q _21094_/X _21095_/X VGND VGND VPWR
+ VPWR _21299_/X sky130_fd_sc_hd__mux4_1
XFILLER_107_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23038_ _23038_/A VGND VGND VPWR VPWR _32070_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27915_ _27751_/X _34297_/Q _27923_/S VGND VGND VPWR VPWR _27916_/A sky130_fd_sc_hd__mux2_1
XTAP_5111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28895_ _34760_/Q _27189_/X _28913_/S VGND VGND VPWR VPWR _28896_/A sky130_fd_sc_hd__mux2_1
XTAP_5122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_493_CLK clkbuf_6_3__f_CLK/X VGND VGND VPWR VPWR _35625_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_5144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27846_ _27649_/X _34264_/Q _27860_/S VGND VGND VPWR VPWR _27847_/A sky130_fd_sc_hd__mux2_1
XFILLER_209_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27777_ _27776_/X _34241_/Q _27795_/S VGND VGND VPWR VPWR _27778_/A sky130_fd_sc_hd__mux2_1
XTAP_4465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24989_ _24988_/X _32979_/Q _24995_/S VGND VGND VPWR VPWR _24990_/A sky130_fd_sc_hd__mux2_1
XTAP_4476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_245_CLK clkbuf_6_61__f_CLK/X VGND VGND VPWR VPWR _33425_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29516_ _35026_/Q _29515_/X _29525_/S VGND VGND VPWR VPWR _29517_/A sky130_fd_sc_hd__mux2_1
XTAP_3753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17530_ _33151_/Q _36031_/Q _33023_/Q _32959_/Q _17415_/X _17416_/X VGND VGND VPWR
+ VPWR _17530_/X sky130_fd_sc_hd__mux4_1
X_26728_ _33797_/Q _23444_/X _26732_/S VGND VGND VPWR VPWR _26729_/A sky130_fd_sc_hd__mux2_1
XTAP_4498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17461_ _35709_/Q _32218_/Q _35581_/Q _35517_/Q _17317_/X _17318_/X VGND VGND VPWR
+ VPWR _17461_/X sky130_fd_sc_hd__mux4_1
X_29447_ input32/X VGND VGND VPWR VPWR _29447_/X sky130_fd_sc_hd__buf_2
X_26659_ _33764_/Q _23274_/X _26669_/S VGND VGND VPWR VPWR _26660_/A sky130_fd_sc_hd__mux2_1
XFILLER_232_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19200_ _18945_/X _19198_/X _19199_/X _18948_/X VGND VGND VPWR VPWR _19200_/X sky130_fd_sc_hd__a22o_1
X_16412_ _34399_/Q _36127_/Q _34271_/Q _34207_/Q _16170_/X _16171_/X VGND VGND VPWR
+ VPWR _16412_/X sky130_fd_sc_hd__mux4_1
XFILLER_60_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29378_ _29378_/A VGND VGND VPWR VPWR _34981_/D sky130_fd_sc_hd__clkbuf_1
X_17392_ _35451_/Q _35387_/Q _35323_/Q _35259_/Q _17254_/X _17255_/X VGND VGND VPWR
+ VPWR _17392_/X sky130_fd_sc_hd__mux4_1
XFILLER_220_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19131_ _35627_/Q _34987_/Q _34347_/Q _33707_/Q _19091_/X _19092_/X VGND VGND VPWR
+ VPWR _19131_/X sky130_fd_sc_hd__mux4_1
X_16343_ _16339_/X _16342_/X _16104_/X VGND VGND VPWR VPWR _16344_/D sky130_fd_sc_hd__o21ba_1
XFILLER_13_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28329_ _28329_/A VGND VGND VPWR VPWR _34493_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16274_ _16274_/A _16274_/B _16274_/C _16274_/D VGND VGND VPWR VPWR _16275_/A sky130_fd_sc_hd__or4_1
X_19062_ _34665_/Q _34601_/Q _34537_/Q _34473_/Q _18886_/X _18887_/X VGND VGND VPWR
+ VPWR _19062_/X sky130_fd_sc_hd__mux4_1
X_31340_ _31340_/A VGND VGND VPWR VPWR _35888_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18013_ _33933_/Q _33869_/Q _33805_/Q _36109_/Q _17730_/X _17731_/X VGND VGND VPWR
+ VPWR _18013_/X sky130_fd_sc_hd__mux4_1
XFILLER_16_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_218_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31271_ _27822_/X _35856_/Q _31273_/S VGND VGND VPWR VPWR _31272_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1086 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33010_ _36017_/CLK _33010_/D VGND VGND VPWR VPWR _33010_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30222_ _35359_/Q _29357_/X _30222_/S VGND VGND VPWR VPWR _30223_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30153_ _35326_/Q _29453_/X _30171_/S VGND VGND VPWR VPWR _30154_/A sky130_fd_sc_hd__mux2_1
X_19964_ _33155_/Q _36035_/Q _33027_/Q _32963_/Q _19715_/X _19716_/X VGND VGND VPWR
+ VPWR _19964_/X sky130_fd_sc_hd__mux4_1
X_18915_ _18592_/X _18913_/X _18914_/X _18595_/X VGND VGND VPWR VPWR _18915_/X sky130_fd_sc_hd__a22o_1
XTAP_7080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34961_ _34961_/CLK _34961_/D VGND VGND VPWR VPWR _34961_/Q sky130_fd_sc_hd__dfxtp_1
X_30084_ _30084_/A VGND VGND VPWR VPWR _35293_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19895_ _19859_/X _19893_/X _19894_/X _19862_/X VGND VGND VPWR VPWR _19895_/X sky130_fd_sc_hd__a22o_1
XFILLER_141_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_484_CLK _35560_/CLK VGND VGND VPWR VPWR _33897_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_95_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33912_ _36090_/CLK _33912_/D VGND VGND VPWR VPWR _33912_/Q sky130_fd_sc_hd__dfxtp_1
X_18846_ _35619_/Q _34979_/Q _34339_/Q _33699_/Q _18738_/X _18739_/X VGND VGND VPWR
+ VPWR _18846_/X sky130_fd_sc_hd__mux4_1
X_34892_ _34957_/CLK _34892_/D VGND VGND VPWR VPWR _34892_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_954 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33843_ _36085_/CLK _33843_/D VGND VGND VPWR VPWR _33843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18777_ _35681_/Q _32188_/Q _35553_/Q _35489_/Q _18558_/X _18559_/X VGND VGND VPWR
+ VPWR _18777_/X sky130_fd_sc_hd__mux4_1
X_15989_ input67/X input68/X VGND VGND VPWR VPWR _17771_/A sky130_fd_sc_hd__nor2_4
XFILLER_209_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_236_CLK clkbuf_6_54__f_CLK/X VGND VGND VPWR VPWR _36165_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17728_ _17552_/X _17726_/X _17727_/X _17557_/X VGND VGND VPWR VPWR _17728_/X sky130_fd_sc_hd__a22o_1
XFILLER_209_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33774_ _36077_/CLK _33774_/D VGND VGND VPWR VPWR _33774_/Q sky130_fd_sc_hd__dfxtp_1
X_30986_ _35721_/Q input47/X _31002_/S VGND VGND VPWR VPWR _30987_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35513_ _35577_/CLK _35513_/D VGND VGND VPWR VPWR _35513_/Q sky130_fd_sc_hd__dfxtp_1
X_32725_ _35989_/CLK _32725_/D VGND VGND VPWR VPWR _32725_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17659_ _33411_/Q _33347_/Q _33283_/Q _33219_/Q _17480_/X _17481_/X VGND VGND VPWR
+ VPWR _17659_/X sky130_fd_sc_hd__mux4_1
XFILLER_35_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35444_ _35446_/CLK _35444_/D VGND VGND VPWR VPWR _35444_/Q sky130_fd_sc_hd__dfxtp_1
X_20670_ _33046_/Q _32022_/Q _35798_/Q _35734_/Q _20667_/X _20669_/X VGND VGND VPWR
+ VPWR _20670_/X sky130_fd_sc_hd__mux4_1
X_32656_ _36049_/CLK _32656_/D VGND VGND VPWR VPWR _32656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31607_ _27720_/X _36015_/Q _31615_/S VGND VGND VPWR VPWR _31608_/A sky130_fd_sc_hd__mux2_1
X_19329_ _32625_/Q _32561_/Q _32497_/Q _35953_/Q _19223_/X _19007_/X VGND VGND VPWR
+ VPWR _19329_/X sky130_fd_sc_hd__mux4_1
X_35375_ _35694_/CLK _35375_/D VGND VGND VPWR VPWR _35375_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32587_ _35980_/CLK _32587_/D VGND VGND VPWR VPWR _32587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34326_ _35673_/CLK _34326_/D VGND VGND VPWR VPWR _34326_/Q sky130_fd_sc_hd__dfxtp_1
X_22340_ _22020_/X _22338_/X _22339_/X _22024_/X VGND VGND VPWR VPWR _22340_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31538_ _31538_/A VGND VGND VPWR VPWR _35982_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34257_ _36177_/CLK _34257_/D VGND VGND VPWR VPWR _34257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22271_ _22400_/A VGND VGND VPWR VPWR _22271_/X sky130_fd_sc_hd__buf_4
XFILLER_192_968 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31469_ _31469_/A VGND VGND VPWR VPWR _35949_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24010_ _24010_/A VGND VGND VPWR VPWR _32547_/D sky130_fd_sc_hd__clkbuf_1
X_33208_ _36090_/CLK _33208_/D VGND VGND VPWR VPWR _33208_/Q sky130_fd_sc_hd__dfxtp_1
X_21222_ _21047_/X _21220_/X _21221_/X _21050_/X VGND VGND VPWR VPWR _21222_/X sky130_fd_sc_hd__a22o_1
XFILLER_219_1314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34188_ _34188_/CLK _34188_/D VGND VGND VPWR VPWR _34188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21153_ _21147_/X _21152_/X _21045_/X VGND VGND VPWR VPWR _21161_/C sky130_fd_sc_hd__o21ba_1
X_33139_ _36020_/CLK _33139_/D VGND VGND VPWR VPWR _33139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20104_ _33927_/Q _33863_/Q _33799_/Q _36103_/Q _20030_/X _20031_/X VGND VGND VPWR
+ VPWR _20104_/X sky130_fd_sc_hd__mux4_1
XFILLER_63_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25961_ _24818_/X _33436_/Q _25967_/S VGND VGND VPWR VPWR _25962_/A sky130_fd_sc_hd__mux2_1
XFILLER_132_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21084_ _34657_/Q _34593_/Q _34529_/Q _34465_/Q _20833_/X _20834_/X VGND VGND VPWR
+ VPWR _21084_/X sky130_fd_sc_hd__mux4_1
XFILLER_8_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_475_CLK clkbuf_6_10__f_CLK/X VGND VGND VPWR VPWR _33902_/CLK sky130_fd_sc_hd__clkbuf_16
X_27700_ _27700_/A VGND VGND VPWR VPWR _34216_/D sky130_fd_sc_hd__clkbuf_1
X_20035_ _32645_/Q _32581_/Q _32517_/Q _35973_/Q _19929_/X _19713_/X VGND VGND VPWR
+ VPWR _20035_/X sky130_fd_sc_hd__mux4_1
XFILLER_115_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24912_ _24911_/X _32954_/Q _24921_/S VGND VGND VPWR VPWR _24913_/A sky130_fd_sc_hd__mux2_1
XFILLER_246_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25892_ _25892_/A VGND VGND VPWR VPWR _33403_/D sky130_fd_sc_hd__clkbuf_1
X_28680_ _34659_/Q _27075_/X _28692_/S VGND VGND VPWR VPWR _28681_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27631_ _34194_/Q _27220_/X _27637_/S VGND VGND VPWR VPWR _27632_/A sky130_fd_sc_hd__mux2_1
XFILLER_218_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24843_ input6/X VGND VGND VPWR VPWR _24843_/X sky130_fd_sc_hd__buf_4
XTAP_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_227_CLK clkbuf_6_55__f_CLK/X VGND VGND VPWR VPWR _34064_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_39_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24774_ _23052_/X _32907_/Q _24786_/S VGND VGND VPWR VPWR _24775_/A sky130_fd_sc_hd__mux2_1
X_27562_ _34161_/Q _27118_/X _27566_/S VGND VGND VPWR VPWR _27563_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21986_ _32891_/Q _32827_/Q _32763_/Q _32699_/Q _21946_/X _21947_/X VGND VGND VPWR
+ VPWR _21986_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_6_57__f_CLK clkbuf_5_28_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_57__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_27_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29301_ _29301_/A VGND VGND VPWR VPWR _34952_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23725_ _22912_/X _32350_/Q _23727_/S VGND VGND VPWR VPWR _23726_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26513_ _26513_/A VGND VGND VPWR VPWR _33696_/D sky130_fd_sc_hd__clkbuf_1
X_20937_ _34653_/Q _34589_/Q _34525_/Q _34461_/Q _20833_/X _20834_/X VGND VGND VPWR
+ VPWR _20937_/X sky130_fd_sc_hd__mux4_1
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27493_ _27493_/A VGND VGND VPWR VPWR _34128_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29232_ _34920_/Q _27090_/X _29234_/S VGND VGND VPWR VPWR _29233_/A sky130_fd_sc_hd__mux2_1
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26444_ _26444_/A VGND VGND VPWR VPWR _33664_/D sky130_fd_sc_hd__clkbuf_1
X_23656_ _23656_/A VGND VGND VPWR VPWR _32318_/D sky130_fd_sc_hd__clkbuf_1
X_20868_ _35163_/Q _35099_/Q _35035_/Q _32155_/Q _20683_/X _20685_/X VGND VGND VPWR
+ VPWR _20868_/X sky130_fd_sc_hd__mux4_1
XFILLER_186_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22607_ _22607_/A _22607_/B _22607_/C _22607_/D VGND VGND VPWR VPWR _22608_/A sky130_fd_sc_hd__or4_4
XFILLER_168_932 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29163_ _29163_/A VGND VGND VPWR VPWR _34887_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26375_ _26486_/S VGND VGND VPWR VPWR _26394_/S sky130_fd_sc_hd__buf_6
XFILLER_35_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23587_ _22912_/X _32286_/Q _23589_/S VGND VGND VPWR VPWR _23588_/A sky130_fd_sc_hd__mux2_1
XFILLER_224_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20799_ _20660_/X _20797_/X _20798_/X _20672_/X VGND VGND VPWR VPWR _20799_/X sky130_fd_sc_hd__a22o_1
X_28114_ _27646_/X _34391_/Q _28130_/S VGND VGND VPWR VPWR _28115_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25326_ _33136_/Q _23340_/X _25332_/S VGND VGND VPWR VPWR _25327_/A sky130_fd_sc_hd__mux2_1
X_22538_ _34954_/Q _34890_/Q _34826_/Q _34762_/Q _22466_/X _22467_/X VGND VGND VPWR
+ VPWR _22538_/X sky130_fd_sc_hd__mux4_1
XFILLER_155_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29094_ _29094_/A VGND VGND VPWR VPWR _34854_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25257_ _33104_/Q _23481_/X _25259_/S VGND VGND VPWR VPWR _25258_/A sky130_fd_sc_hd__mux2_1
X_28045_ _28045_/A VGND VGND VPWR VPWR _34358_/D sky130_fd_sc_hd__clkbuf_1
X_22469_ _22469_/A VGND VGND VPWR VPWR _22469_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_154_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24208_ _32640_/Q _23429_/X _24222_/S VGND VGND VPWR VPWR _24209_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25188_ _33071_/Q _23316_/X _25196_/S VGND VGND VPWR VPWR _25189_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24139_ _24139_/A VGND VGND VPWR VPWR _32607_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1008 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29996_ _30065_/S VGND VGND VPWR VPWR _30015_/S sky130_fd_sc_hd__buf_6
XFILLER_150_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28947_ _28947_/A VGND VGND VPWR VPWR _34784_/D sky130_fd_sc_hd__clkbuf_1
X_16961_ _32879_/Q _32815_/Q _32751_/Q _32687_/Q _16640_/X _16641_/X VGND VGND VPWR
+ VPWR _16961_/X sky130_fd_sc_hd__mux4_1
X_18700_ _18661_/X _18698_/X _18699_/X _18665_/X VGND VGND VPWR VPWR _18700_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_466_CLK clkbuf_6_11__f_CLK/X VGND VGND VPWR VPWR _35181_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_238_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19680_ _19506_/X _19676_/X _19679_/X _19509_/X VGND VGND VPWR VPWR _19680_/X sky130_fd_sc_hd__a22o_1
XFILLER_231_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28878_ _34752_/Q _27165_/X _28892_/S VGND VGND VPWR VPWR _28879_/A sky130_fd_sc_hd__mux2_1
X_16892_ _33133_/Q _36013_/Q _33005_/Q _32941_/Q _16709_/X _16710_/X VGND VGND VPWR
+ VPWR _16892_/X sky130_fd_sc_hd__mux4_1
XFILLER_204_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18631_ _35613_/Q _34973_/Q _34333_/Q _33693_/Q _18353_/X _18355_/X VGND VGND VPWR
+ VPWR _18631_/X sky130_fd_sc_hd__mux4_1
X_27829_ _27828_/X _34258_/Q _27838_/S VGND VGND VPWR VPWR _27830_/A sky130_fd_sc_hd__mux2_1
XTAP_4240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_218_CLK clkbuf_6_53__f_CLK/X VGND VGND VPWR VPWR _36169_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_58_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18562_ _18348_/X _18560_/X _18561_/X _18358_/X VGND VGND VPWR VPWR _18562_/X sky130_fd_sc_hd__a22o_1
X_30840_ _35652_/Q input41/X _30846_/S VGND VGND VPWR VPWR _30841_/A sky130_fd_sc_hd__mux2_1
XTAP_4284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1096 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17513_ _17866_/A VGND VGND VPWR VPWR _17513_/X sky130_fd_sc_hd__buf_4
XTAP_3583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18493_ _35609_/Q _34969_/Q _34329_/Q _33689_/Q _18353_/X _18355_/X VGND VGND VPWR
+ VPWR _18493_/X sky130_fd_sc_hd__mux4_1
XTAP_3594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30771_ _35619_/Q input5/X _30783_/S VGND VGND VPWR VPWR _30772_/A sky130_fd_sc_hd__mux2_1
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32510_ _36031_/CLK _32510_/D VGND VGND VPWR VPWR _32510_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17444_ _17444_/A VGND VGND VPWR VPWR _31996_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33490_ _33875_/CLK _33490_/D VGND VGND VPWR VPWR _33490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32441_ _33895_/CLK _32441_/D VGND VGND VPWR VPWR _32441_/Q sky130_fd_sc_hd__dfxtp_1
X_17375_ _17199_/X _17373_/X _17374_/X _17204_/X VGND VGND VPWR VPWR _17375_/X sky130_fd_sc_hd__a22o_1
XFILLER_229_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_807 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19114_ _19114_/A _19114_/B _19114_/C _19114_/D VGND VGND VPWR VPWR _19115_/A sky130_fd_sc_hd__or4_2
X_35160_ _35160_/CLK _35160_/D VGND VGND VPWR VPWR _35160_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16326_ _32093_/Q _32285_/Q _32349_/Q _35869_/Q _16221_/X _17867_/A VGND VGND VPWR
+ VPWR _16326_/X sky130_fd_sc_hd__mux4_1
X_32372_ _32882_/CLK _32372_/D VGND VGND VPWR VPWR _32372_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34111_ _35454_/CLK _34111_/D VGND VGND VPWR VPWR _34111_/Q sky130_fd_sc_hd__dfxtp_1
X_19045_ _33897_/Q _33833_/Q _33769_/Q _36073_/Q _18971_/X _18972_/X VGND VGND VPWR
+ VPWR _19045_/X sky130_fd_sc_hd__mux4_1
X_31323_ _31323_/A VGND VGND VPWR VPWR _35880_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_199_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35091_ _36114_/CLK _35091_/D VGND VGND VPWR VPWR _35091_/Q sky130_fd_sc_hd__dfxtp_1
X_16257_ _16253_/X _16256_/X _16044_/X _16046_/X VGND VGND VPWR VPWR _16274_/B sky130_fd_sc_hd__o211a_1
XFILLER_174_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34042_ _35320_/CLK _34042_/D VGND VGND VPWR VPWR _34042_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput204 _36237_/Q VGND VGND VPWR VPWR D2[55] sky130_fd_sc_hd__buf_2
X_31254_ _31281_/S VGND VGND VPWR VPWR _31273_/S sky130_fd_sc_hd__buf_4
X_16188_ _32089_/Q _32281_/Q _32345_/Q _35865_/Q _16032_/X _17867_/A VGND VGND VPWR
+ VPWR _16188_/X sky130_fd_sc_hd__mux4_1
Xoutput215 _36189_/Q VGND VGND VPWR VPWR D2[7] sky130_fd_sc_hd__buf_2
Xoutput226 _32423_/Q VGND VGND VPWR VPWR D3[17] sky130_fd_sc_hd__buf_2
XFILLER_99_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30205_ _30205_/A VGND VGND VPWR VPWR _35350_/D sky130_fd_sc_hd__clkbuf_1
Xoutput237 _32433_/Q VGND VGND VPWR VPWR D3[27] sky130_fd_sc_hd__buf_2
XFILLER_126_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput248 _32443_/Q VGND VGND VPWR VPWR D3[37] sky130_fd_sc_hd__buf_2
XFILLER_114_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput259 _32453_/Q VGND VGND VPWR VPWR D3[47] sky130_fd_sc_hd__buf_2
X_31185_ _27695_/X _35815_/Q _31189_/S VGND VGND VPWR VPWR _31186_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19947_ _34690_/Q _34626_/Q _34562_/Q _34498_/Q _19945_/X _19946_/X VGND VGND VPWR
+ VPWR _19947_/X sky130_fd_sc_hd__mux4_1
XFILLER_4_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30136_ _35318_/Q _29429_/X _30150_/S VGND VGND VPWR VPWR _30137_/A sky130_fd_sc_hd__mux2_1
X_35993_ _35993_/CLK _35993_/D VGND VGND VPWR VPWR _35993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_457_CLK clkbuf_leaf_49_CLK/A VGND VGND VPWR VPWR _35820_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_96_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34944_ _36161_/CLK _34944_/D VGND VGND VPWR VPWR _34944_/Q sky130_fd_sc_hd__dfxtp_1
X_30067_ _30877_/A _31147_/B VGND VGND VPWR VPWR _30200_/S sky130_fd_sc_hd__nor2_8
X_19878_ _19874_/X _19877_/X _19804_/X VGND VGND VPWR VPWR _19888_/C sky130_fd_sc_hd__o21ba_1
XFILLER_95_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18829_ _18829_/A _18829_/B _18829_/C _18829_/D VGND VGND VPWR VPWR _18830_/A sky130_fd_sc_hd__or4_2
XFILLER_95_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34875_ _34941_/CLK _34875_/D VGND VGND VPWR VPWR _34875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_243_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_209_CLK clkbuf_6_54__f_CLK/X VGND VGND VPWR VPWR _34698_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33826_ _36066_/CLK _33826_/D VGND VGND VPWR VPWR _33826_/Q sky130_fd_sc_hd__dfxtp_1
X_21840_ _33399_/Q _33335_/Q _33271_/Q _33207_/Q _21727_/X _21728_/X VGND VGND VPWR
+ VPWR _21840_/X sky130_fd_sc_hd__mux4_1
XFILLER_243_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33757_ _33821_/CLK _33757_/D VGND VGND VPWR VPWR _33757_/Q sky130_fd_sc_hd__dfxtp_1
X_21771_ _21446_/X _21769_/X _21770_/X _21451_/X VGND VGND VPWR VPWR _21771_/X sky130_fd_sc_hd__a22o_1
X_30969_ _35713_/Q input38/X _30981_/S VGND VGND VPWR VPWR _30970_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_1354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23510_ _23510_/A VGND VGND VPWR VPWR _32250_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_212_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20722_ _20630_/X _20720_/X _20721_/X _20641_/X VGND VGND VPWR VPWR _20722_/X sky130_fd_sc_hd__a22o_1
X_32708_ _35973_/CLK _32708_/D VGND VGND VPWR VPWR _32708_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24490_ _24490_/A VGND VGND VPWR VPWR _32772_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33688_ _35609_/CLK _33688_/D VGND VGND VPWR VPWR _33688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_1218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23441_ input41/X VGND VGND VPWR VPWR _23441_/X sky130_fd_sc_hd__buf_6
XFILLER_17_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35427_ _35814_/CLK _35427_/D VGND VGND VPWR VPWR _35427_/Q sky130_fd_sc_hd__dfxtp_1
X_20653_ _22598_/A VGND VGND VPWR VPWR _20653_/X sky130_fd_sc_hd__buf_6
X_32639_ _35903_/CLK _32639_/D VGND VGND VPWR VPWR _32639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26160_ _26160_/A VGND VGND VPWR VPWR _33530_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35358_ _35677_/CLK _35358_/D VGND VGND VPWR VPWR _35358_/Q sky130_fd_sc_hd__dfxtp_1
X_23372_ _23372_/A VGND VGND VPWR VPWR _32201_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_176_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20584_ _22506_/A VGND VGND VPWR VPWR _20584_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_176_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25111_ _25111_/A VGND VGND VPWR VPWR _33035_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34309_ _36165_/CLK _34309_/D VGND VGND VPWR VPWR _34309_/Q sky130_fd_sc_hd__dfxtp_1
X_22323_ _22319_/X _22322_/X _22118_/X VGND VGND VPWR VPWR _22324_/D sky130_fd_sc_hd__o21ba_1
XFILLER_99_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26091_ _26091_/A VGND VGND VPWR VPWR _33497_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35289_ _35674_/CLK _35289_/D VGND VGND VPWR VPWR _35289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25042_ _25042_/A VGND VGND VPWR VPWR _33002_/D sky130_fd_sc_hd__clkbuf_1
X_22254_ _22254_/A _22254_/B _22254_/C _22254_/D VGND VGND VPWR VPWR _22255_/A sky130_fd_sc_hd__or4_4
XFILLER_3_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21205_ _33125_/Q _36005_/Q _32997_/Q _32933_/Q _20956_/X _20957_/X VGND VGND VPWR
+ VPWR _21205_/X sky130_fd_sc_hd__mux4_1
XFILLER_155_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29850_ _29850_/A VGND VGND VPWR VPWR _35182_/D sky130_fd_sc_hd__clkbuf_1
X_22185_ _34944_/Q _34880_/Q _34816_/Q _34752_/Q _22113_/X _22114_/X VGND VGND VPWR
+ VPWR _22185_/X sky130_fd_sc_hd__mux4_1
X_28801_ _28801_/A VGND VGND VPWR VPWR _34715_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21136_ _21100_/X _21134_/X _21135_/X _21103_/X VGND VGND VPWR VPWR _21136_/X sky130_fd_sc_hd__a22o_1
X_29781_ _35150_/Q _29503_/X _29787_/S VGND VGND VPWR VPWR _29782_/A sky130_fd_sc_hd__mux2_1
X_26993_ _26993_/A VGND VGND VPWR VPWR _33922_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_448_CLK clkbuf_leaf_61_CLK/A VGND VGND VPWR VPWR _35883_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_247_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28732_ _34684_/Q _27152_/X _28734_/S VGND VGND VPWR VPWR _28733_/A sky130_fd_sc_hd__mux2_1
X_25944_ _25944_/A VGND VGND VPWR VPWR _33428_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21067_ _33889_/Q _33825_/Q _33761_/Q _36065_/Q _20918_/X _20919_/X VGND VGND VPWR
+ VPWR _21067_/X sky130_fd_sc_hd__mux4_1
XFILLER_24_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20018_ _35204_/Q _35140_/Q _35076_/Q _32260_/Q _20016_/X _20017_/X VGND VGND VPWR
+ VPWR _20018_/X sky130_fd_sc_hd__mux4_1
XFILLER_171_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28663_ _34651_/Q _27050_/X _28671_/S VGND VGND VPWR VPWR _28664_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25875_ _25875_/A VGND VGND VPWR VPWR _33395_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27614_ _27614_/A VGND VGND VPWR VPWR _34185_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_230_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24826_ _24826_/A VGND VGND VPWR VPWR _32926_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28594_ _27757_/X _34619_/Q _28598_/S VGND VGND VPWR VPWR _28595_/A sky130_fd_sc_hd__mux2_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27545_ _34153_/Q _27093_/X _27545_/S VGND VGND VPWR VPWR _27546_/A sky130_fd_sc_hd__mux2_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24757_ _23027_/X _32899_/Q _24765_/S VGND VGND VPWR VPWR _24758_/A sky130_fd_sc_hd__mux2_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21969_ _21758_/X _21967_/X _21968_/X _21763_/X VGND VGND VPWR VPWR _21969_/X sky130_fd_sc_hd__a22o_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23708_ _23840_/S VGND VGND VPWR VPWR _23727_/S sky130_fd_sc_hd__buf_4
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27476_ _34120_/Q _27189_/X _27494_/S VGND VGND VPWR VPWR _27477_/A sky130_fd_sc_hd__mux2_1
XFILLER_203_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24688_ _22925_/X _32866_/Q _24702_/S VGND VGND VPWR VPWR _24689_/A sky130_fd_sc_hd__mux2_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29215_ _29326_/S VGND VGND VPWR VPWR _29234_/S sky130_fd_sc_hd__buf_4
XFILLER_70_885 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26427_ _26427_/A VGND VGND VPWR VPWR _33656_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23639_ _23639_/A VGND VGND VPWR VPWR _32310_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_230_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29146_ _34879_/Q _27162_/X _29162_/S VGND VGND VPWR VPWR _29147_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_1282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17160_ _17866_/A VGND VGND VPWR VPWR _17160_/X sky130_fd_sc_hd__buf_4
X_26358_ _26358_/A VGND VGND VPWR VPWR _33623_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16111_ _33367_/Q _33303_/Q _33239_/Q _33175_/Q _16002_/X _16003_/X VGND VGND VPWR
+ VPWR _16111_/X sky130_fd_sc_hd__mux4_1
XFILLER_70_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25309_ _33128_/Q _23286_/X _25311_/S VGND VGND VPWR VPWR _25310_/A sky130_fd_sc_hd__mux2_1
X_29077_ _29077_/A VGND VGND VPWR VPWR _34846_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26289_ _26289_/A VGND VGND VPWR VPWR _33591_/D sky130_fd_sc_hd__clkbuf_1
X_17091_ _17091_/A VGND VGND VPWR VPWR _31986_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16042_ _16030_/X _16035_/X _16040_/X _16041_/X VGND VGND VPWR VPWR _16042_/X sky130_fd_sc_hd__a22o_1
XFILLER_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28028_ _28028_/A VGND VGND VPWR VPWR _34350_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_938 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19801_ _35454_/Q _35390_/Q _35326_/Q _35262_/Q _19554_/X _19555_/X VGND VGND VPWR
+ VPWR _19801_/X sky130_fd_sc_hd__mux4_1
XFILLER_215_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17993_ _17704_/X _17991_/X _17992_/X _17707_/X VGND VGND VPWR VPWR _17993_/X sky130_fd_sc_hd__a22o_1
X_29979_ _29979_/A VGND VGND VPWR VPWR _35243_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_439_CLK clkbuf_6_36__f_CLK/X VGND VGND VPWR VPWR _36017_/CLK sky130_fd_sc_hd__clkbuf_16
X_19732_ _20236_/A VGND VGND VPWR VPWR _19732_/X sky130_fd_sc_hd__buf_4
XFILLER_111_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16944_ _34414_/Q _36142_/Q _34286_/Q _34222_/Q _16876_/X _16877_/X VGND VGND VPWR
+ VPWR _16944_/X sky130_fd_sc_hd__mux4_1
X_32990_ _33119_/CLK _32990_/D VGND VGND VPWR VPWR _32990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31941_ _31941_/A VGND VGND VPWR VPWR _36173_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_1275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19663_ _20016_/A VGND VGND VPWR VPWR _19663_/X sky130_fd_sc_hd__buf_6
X_16875_ _16800_/X _16873_/X _16874_/X _16803_/X VGND VGND VPWR VPWR _16875_/X sky130_fd_sc_hd__a22o_1
XFILLER_65_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18614_ _33629_/Q _33565_/Q _33501_/Q _33437_/Q _18441_/X _18442_/X VGND VGND VPWR
+ VPWR _18614_/X sky130_fd_sc_hd__mux4_1
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34660_ _34913_/CLK _34660_/D VGND VGND VPWR VPWR _34660_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19594_ _34680_/Q _34616_/Q _34552_/Q _34488_/Q _19592_/X _19593_/X VGND VGND VPWR
+ VPWR _19594_/X sky130_fd_sc_hd__mux4_1
X_31872_ _31872_/A VGND VGND VPWR VPWR _36140_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33611_ _34187_/CLK _33611_/D VGND VGND VPWR VPWR _33611_/Q sky130_fd_sc_hd__dfxtp_1
X_18545_ _34139_/Q _34075_/Q _34011_/Q _33947_/Q _18309_/X _18311_/X VGND VGND VPWR
+ VPWR _18545_/X sky130_fd_sc_hd__mux4_1
XFILLER_52_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30823_ _35644_/Q input32/X _30825_/S VGND VGND VPWR VPWR _30824_/A sky130_fd_sc_hd__mux2_1
X_34591_ _35544_/CLK _34591_/D VGND VGND VPWR VPWR _34591_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_40__f_CLK clkbuf_5_20_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_40__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_209_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33542_ _34179_/CLK _33542_/D VGND VGND VPWR VPWR _33542_/Q sky130_fd_sc_hd__dfxtp_1
X_18476_ _18476_/A _18476_/B _18476_/C _18476_/D VGND VGND VPWR VPWR _18477_/A sky130_fd_sc_hd__or4_1
X_30754_ _35611_/Q input56/X _30762_/S VGND VGND VPWR VPWR _30755_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_863 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17427_ _35708_/Q _32217_/Q _35580_/Q _35516_/Q _17317_/X _17318_/X VGND VGND VPWR
+ VPWR _17427_/X sky130_fd_sc_hd__mux4_1
X_33473_ _34180_/CLK _33473_/D VGND VGND VPWR VPWR _33473_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30685_ _30685_/A VGND VGND VPWR VPWR _35578_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35212_ _35212_/CLK _35212_/D VGND VGND VPWR VPWR _35212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32424_ _36068_/CLK _32424_/D VGND VGND VPWR VPWR _32424_/Q sky130_fd_sc_hd__dfxtp_1
X_36192_ _36207_/CLK _36192_/D VGND VGND VPWR VPWR _36192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17358_ _33082_/Q _32058_/Q _35834_/Q _35770_/Q _17078_/X _17079_/X VGND VGND VPWR
+ VPWR _17358_/X sky130_fd_sc_hd__mux4_1
XFILLER_174_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16309_ _34908_/Q _34844_/Q _34780_/Q _34716_/Q _16096_/X _16098_/X VGND VGND VPWR
+ VPWR _16309_/X sky130_fd_sc_hd__mux4_1
X_35143_ _35657_/CLK _35143_/D VGND VGND VPWR VPWR _35143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32355_ _32356_/CLK _32355_/D VGND VGND VPWR VPWR _32355_/Q sky130_fd_sc_hd__dfxtp_1
X_17289_ _33080_/Q _32056_/Q _35832_/Q _35768_/Q _17078_/X _17079_/X VGND VGND VPWR
+ VPWR _17289_/X sky130_fd_sc_hd__mux4_1
X_31306_ _27673_/X _35872_/Q _31324_/S VGND VGND VPWR VPWR _31307_/A sky130_fd_sc_hd__mux2_1
X_19028_ _18950_/X _19024_/X _19027_/X _18953_/X VGND VGND VPWR VPWR _19028_/X sky130_fd_sc_hd__a22o_1
X_35074_ _35655_/CLK _35074_/D VGND VGND VPWR VPWR _35074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32286_ _35870_/CLK _32286_/D VGND VGND VPWR VPWR _32286_/Q sky130_fd_sc_hd__dfxtp_1
X_34025_ _35624_/CLK _34025_/D VGND VGND VPWR VPWR _34025_/Q sky130_fd_sc_hd__dfxtp_1
X_31237_ _31237_/A VGND VGND VPWR VPWR _35839_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31168_ _27670_/X _35807_/Q _31168_/S VGND VGND VPWR VPWR _31169_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30119_ _35310_/Q _29404_/X _30129_/S VGND VGND VPWR VPWR _30120_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23990_ _22900_/X _32538_/Q _24000_/S VGND VGND VPWR VPWR _23991_/A sky130_fd_sc_hd__mux2_1
X_35976_ _35976_/CLK _35976_/D VGND VGND VPWR VPWR _35976_/Q sky130_fd_sc_hd__dfxtp_1
X_31099_ _31099_/A VGND VGND VPWR VPWR _35774_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22941_ _22940_/X _32039_/Q _22947_/S VGND VGND VPWR VPWR _22942_/A sky130_fd_sc_hd__mux2_1
X_34927_ _34927_/CLK _34927_/D VGND VGND VPWR VPWR _34927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_928 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25660_ _25660_/A VGND VGND VPWR VPWR _33293_/D sky130_fd_sc_hd__clkbuf_1
X_22872_ _20648_/X _22870_/X _22871_/X _20658_/X VGND VGND VPWR VPWR _22872_/X sky130_fd_sc_hd__a22o_1
XFILLER_186_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34858_ _35692_/CLK _34858_/D VGND VGND VPWR VPWR _34858_/Q sky130_fd_sc_hd__dfxtp_1
X_24611_ _24659_/S VGND VGND VPWR VPWR _24630_/S sky130_fd_sc_hd__buf_4
X_21823_ _33078_/Q _32054_/Q _35830_/Q _35766_/Q _21678_/X _21679_/X VGND VGND VPWR
+ VPWR _21823_/X sky130_fd_sc_hd__mux4_1
X_33809_ _34440_/CLK _33809_/D VGND VGND VPWR VPWR _33809_/Q sky130_fd_sc_hd__dfxtp_1
X_25591_ _25591_/A VGND VGND VPWR VPWR _33260_/D sky130_fd_sc_hd__clkbuf_1
X_34789_ _34790_/CLK _34789_/D VGND VGND VPWR VPWR _34789_/Q sky130_fd_sc_hd__dfxtp_1
X_27330_ _34051_/Q _27174_/X _27338_/S VGND VGND VPWR VPWR _27331_/A sky130_fd_sc_hd__mux2_1
X_24542_ _22909_/X _32797_/Q _24546_/S VGND VGND VPWR VPWR _24543_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21754_ _34676_/Q _34612_/Q _34548_/Q _34484_/Q _21539_/X _21540_/X VGND VGND VPWR
+ VPWR _21754_/X sky130_fd_sc_hd__mux4_1
XFILLER_227_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20705_ _20689_/X _20702_/X _20704_/X VGND VGND VPWR VPWR _20706_/D sky130_fd_sc_hd__o21ba_1
XFILLER_52_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27261_ _34018_/Q _27072_/X _27275_/S VGND VGND VPWR VPWR _27262_/A sky130_fd_sc_hd__mux2_1
X_24473_ _24473_/A VGND VGND VPWR VPWR _32764_/D sky130_fd_sc_hd__clkbuf_1
X_21685_ _21400_/X _21683_/X _21684_/X _21403_/X VGND VGND VPWR VPWR _21685_/X sky130_fd_sc_hd__a22o_1
XFILLER_138_902 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29000_ _34810_/Q _27146_/X _29006_/S VGND VGND VPWR VPWR _29001_/A sky130_fd_sc_hd__mux2_1
X_26212_ _26212_/A VGND VGND VPWR VPWR _33555_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23424_ _32220_/Q _23384_/X _23424_/S VGND VGND VPWR VPWR _23425_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27192_ _27192_/A VGND VGND VPWR VPWR _33992_/D sky130_fd_sc_hd__clkbuf_1
X_20636_ _20661_/A VGND VGND VPWR VPWR _22433_/A sky130_fd_sc_hd__buf_12
XFILLER_123_1433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26143_ _26143_/A VGND VGND VPWR VPWR _33522_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23355_ _32194_/Q _23283_/X _23359_/S VGND VGND VPWR VPWR _23356_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20567_ _33109_/Q _32085_/Q _35861_/Q _35797_/Q _18379_/X _18380_/X VGND VGND VPWR
+ VPWR _20567_/X sky130_fd_sc_hd__mux4_1
XFILLER_221_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22306_ _35652_/Q _35012_/Q _34372_/Q _33732_/Q _22097_/X _22098_/X VGND VGND VPWR
+ VPWR _22306_/X sky130_fd_sc_hd__mux4_1
XFILLER_166_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26074_ _24985_/X _33490_/Q _26080_/S VGND VGND VPWR VPWR _26075_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23286_ input10/X VGND VGND VPWR VPWR _23286_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_164_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20498_ _19453_/A _20496_/X _20497_/X _19456_/A VGND VGND VPWR VPWR _20498_/X sky130_fd_sc_hd__a22o_1
X_29902_ _29902_/A VGND VGND VPWR VPWR _35207_/D sky130_fd_sc_hd__clkbuf_1
X_25025_ _25025_/A VGND VGND VPWR VPWR _32994_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22237_ _22232_/X _22236_/X _22093_/X _22094_/X VGND VGND VPWR VPWR _22254_/B sky130_fd_sc_hd__o211a_1
XFILLER_65_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29833_ _29833_/A VGND VGND VPWR VPWR _35174_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22168_ _32128_/Q _32320_/Q _32384_/Q _35904_/Q _21880_/X _22021_/X VGND VGND VPWR
+ VPWR _22168_/X sky130_fd_sc_hd__mux4_1
XFILLER_120_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21119_ _21115_/X _21118_/X _21045_/X VGND VGND VPWR VPWR _21129_/C sky130_fd_sc_hd__o21ba_1
XTAP_6967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29764_ _35142_/Q _29478_/X _29766_/S VGND VGND VPWR VPWR _29765_/A sky130_fd_sc_hd__mux2_1
XTAP_6978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22099_ _35646_/Q _35006_/Q _34366_/Q _33726_/Q _22097_/X _22098_/X VGND VGND VPWR
+ VPWR _22099_/X sky130_fd_sc_hd__mux4_1
X_26976_ _26976_/A VGND VGND VPWR VPWR _33914_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28715_ _28784_/S VGND VGND VPWR VPWR _28734_/S sky130_fd_sc_hd__buf_4
XFILLER_247_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25927_ _24967_/X _33420_/Q _25937_/S VGND VGND VPWR VPWR _25928_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29695_ _35109_/Q _29376_/X _29703_/S VGND VGND VPWR VPWR _29696_/A sky130_fd_sc_hd__mux2_1
XFILLER_219_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28646_ _27834_/X _34644_/Q _28648_/S VGND VGND VPWR VPWR _28647_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16660_ _16447_/X _16656_/X _16659_/X _16450_/X VGND VGND VPWR VPWR _16660_/X sky130_fd_sc_hd__a22o_1
XFILLER_210_1450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25858_ _24865_/X _33387_/Q _25874_/S VGND VGND VPWR VPWR _25859_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_903 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24809_ input34/X VGND VGND VPWR VPWR _24809_/X sky130_fd_sc_hd__clkbuf_4
X_28577_ _27732_/X _34611_/Q _28577_/S VGND VGND VPWR VPWR _28578_/A sky130_fd_sc_hd__mux2_1
X_16591_ _34404_/Q _36132_/Q _34276_/Q _34212_/Q _16523_/X _16524_/X VGND VGND VPWR
+ VPWR _16591_/X sky130_fd_sc_hd__mux4_1
X_25789_ _25789_/A VGND VGND VPWR VPWR _33354_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_222_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18330_ _20212_/A VGND VGND VPWR VPWR _18330_/X sky130_fd_sc_hd__buf_4
XFILLER_188_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27528_ _27528_/A VGND VGND VPWR VPWR _34144_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18261_ _17158_/A _18259_/X _18260_/X _17163_/A VGND VGND VPWR VPWR _18261_/X sky130_fd_sc_hd__a22o_1
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27459_ _34112_/Q _27165_/X _27473_/S VGND VGND VPWR VPWR _27460_/A sky130_fd_sc_hd__mux2_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17212_ _32630_/Q _32566_/Q _32502_/Q _35958_/Q _16923_/X _17060_/X VGND VGND VPWR
+ VPWR _17212_/X sky130_fd_sc_hd__mux4_1
XFILLER_129_913 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18192_ _33427_/Q _33363_/Q _33299_/Q _33235_/Q _16037_/X _16039_/X VGND VGND VPWR
+ VPWR _18192_/X sky130_fd_sc_hd__mux4_1
X_30470_ _35477_/Q _29524_/X _30470_/S VGND VGND VPWR VPWR _30471_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17143_ _35700_/Q _32208_/Q _35572_/Q _35508_/Q _16964_/X _16965_/X VGND VGND VPWR
+ VPWR _17143_/X sky130_fd_sc_hd__mux4_1
X_29129_ _34871_/Q _27137_/X _29141_/S VGND VGND VPWR VPWR _29130_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32140_ _32909_/CLK _32140_/D VGND VGND VPWR VPWR _32140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17074_ _35698_/Q _32206_/Q _35570_/Q _35506_/Q _16964_/X _16965_/X VGND VGND VPWR
+ VPWR _17074_/X sky130_fd_sc_hd__mux4_1
XFILLER_7_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16025_ _17907_/A VGND VGND VPWR VPWR _16025_/X sky130_fd_sc_hd__buf_4
XFILLER_237_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32071_ _35974_/CLK _32071_/D VGND VGND VPWR VPWR _32071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_1214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31022_ _35738_/Q input45/X _31032_/S VGND VGND VPWR VPWR _31023_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_1326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35830_ _35830_/CLK _35830_/D VGND VGND VPWR VPWR _35830_/Q sky130_fd_sc_hd__dfxtp_1
X_17976_ _34188_/Q _34124_/Q _34060_/Q _33996_/Q _17799_/X _17800_/X VGND VGND VPWR
+ VPWR _17976_/X sky130_fd_sc_hd__mux4_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19715_ _20286_/A VGND VGND VPWR VPWR _19715_/X sky130_fd_sc_hd__buf_6
X_16927_ _17986_/A VGND VGND VPWR VPWR _16927_/X sky130_fd_sc_hd__buf_6
X_32973_ _36045_/CLK _32973_/D VGND VGND VPWR VPWR _32973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35761_ _36147_/CLK _35761_/D VGND VGND VPWR VPWR _35761_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34712_ _34907_/CLK _34712_/D VGND VGND VPWR VPWR _34712_/Q sky130_fd_sc_hd__dfxtp_1
X_31924_ _31924_/A VGND VGND VPWR VPWR _36165_/D sky130_fd_sc_hd__clkbuf_1
X_19646_ _20133_/A VGND VGND VPWR VPWR _19646_/X sky130_fd_sc_hd__buf_4
X_16858_ _16852_/X _16857_/X _16779_/X VGND VGND VPWR VPWR _16882_/A sky130_fd_sc_hd__o21ba_1
X_35692_ _35692_/CLK _35692_/D VGND VGND VPWR VPWR _35692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34643_ _36115_/CLK _34643_/D VGND VGND VPWR VPWR _34643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31855_ _31855_/A VGND VGND VPWR VPWR _36132_/D sky130_fd_sc_hd__clkbuf_1
X_19577_ _32632_/Q _32568_/Q _32504_/Q _35960_/Q _19576_/X _19360_/X VGND VGND VPWR
+ VPWR _19577_/X sky130_fd_sc_hd__mux4_1
XFILLER_94_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16789_ _16783_/X _16786_/X _16787_/X _16788_/X VGND VGND VPWR VPWR _16814_/B sky130_fd_sc_hd__o211a_1
XFILLER_207_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18528_ _18348_/X _18526_/X _18527_/X _18358_/X VGND VGND VPWR VPWR _18528_/X sky130_fd_sc_hd__a22o_1
X_30806_ _30875_/S VGND VGND VPWR VPWR _30825_/S sky130_fd_sc_hd__buf_6
X_34574_ _35664_/CLK _34574_/D VGND VGND VPWR VPWR _34574_/Q sky130_fd_sc_hd__dfxtp_1
X_31786_ _36100_/Q input41/X _31792_/S VGND VGND VPWR VPWR _31787_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33525_ _34099_/CLK _33525_/D VGND VGND VPWR VPWR _33525_/Q sky130_fd_sc_hd__dfxtp_1
X_18459_ _18455_/X _18458_/X _18344_/X _18346_/X VGND VGND VPWR VPWR _18476_/B sky130_fd_sc_hd__o211a_1
X_30737_ _30737_/A VGND VGND VPWR VPWR _35603_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36244_ _36245_/CLK _36244_/D VGND VGND VPWR VPWR _36244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33456_ _34035_/CLK _33456_/D VGND VGND VPWR VPWR _33456_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21470_ _33068_/Q _32044_/Q _35820_/Q _35756_/Q _21325_/X _21326_/X VGND VGND VPWR
+ VPWR _21470_/X sky130_fd_sc_hd__mux4_1
XFILLER_119_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30668_ _30668_/A VGND VGND VPWR VPWR _35570_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20421_ _35216_/Q _35152_/Q _35088_/Q _32272_/Q _18392_/X _18394_/X VGND VGND VPWR
+ VPWR _20421_/X sky130_fd_sc_hd__mux4_1
X_32407_ _34148_/CLK _32407_/D VGND VGND VPWR VPWR _32407_/Q sky130_fd_sc_hd__dfxtp_1
X_36175_ _36175_/CLK _36175_/D VGND VGND VPWR VPWR _36175_/Q sky130_fd_sc_hd__dfxtp_1
X_33387_ _36076_/CLK _33387_/D VGND VGND VPWR VPWR _33387_/Q sky130_fd_sc_hd__dfxtp_1
X_30599_ _35538_/Q _29515_/X _30605_/S VGND VGND VPWR VPWR _30600_/A sky130_fd_sc_hd__mux2_1
XFILLER_179_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35126_ _35126_/CLK _35126_/D VGND VGND VPWR VPWR _35126_/Q sky130_fd_sc_hd__dfxtp_1
X_23140_ _22959_/X _32109_/Q _23152_/S VGND VGND VPWR VPWR _23141_/A sky130_fd_sc_hd__mux2_1
X_20352_ _20348_/X _20351_/X _20146_/X _20147_/X VGND VGND VPWR VPWR _20367_/B sky130_fd_sc_hd__o211a_1
X_32338_ _35922_/CLK _32338_/D VGND VGND VPWR VPWR _32338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23071_ _23070_/X _32081_/Q _23071_/S VGND VGND VPWR VPWR _23072_/A sky130_fd_sc_hd__mux2_1
X_35057_ _35377_/CLK _35057_/D VGND VGND VPWR VPWR _35057_/Q sky130_fd_sc_hd__dfxtp_1
X_32269_ _35213_/CLK _32269_/D VGND VGND VPWR VPWR _32269_/Q sky130_fd_sc_hd__dfxtp_1
X_20283_ _32652_/Q _32588_/Q _32524_/Q _35980_/Q _20282_/X _20066_/X VGND VGND VPWR
+ VPWR _20283_/X sky130_fd_sc_hd__mux4_1
XTAP_6208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34008_ _34331_/CLK _34008_/D VGND VGND VPWR VPWR _34008_/Q sky130_fd_sc_hd__dfxtp_1
X_22022_ _32124_/Q _32316_/Q _32380_/Q _35900_/Q _21880_/X _22021_/X VGND VGND VPWR
+ VPWR _22022_/X sky130_fd_sc_hd__mux4_1
XTAP_6219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26830_ _33845_/Q _23393_/X _26846_/S VGND VGND VPWR VPWR _26831_/A sky130_fd_sc_hd__mux2_1
XTAP_5529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26761_ _33813_/Q _23498_/X _26761_/S VGND VGND VPWR VPWR _26762_/A sky130_fd_sc_hd__mux2_1
XTAP_4828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23973_ _23076_/X _32531_/Q _23977_/S VGND VGND VPWR VPWR _23974_/A sky130_fd_sc_hd__mux2_1
X_35959_ _36023_/CLK _35959_/D VGND VGND VPWR VPWR _35959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28500_ _28500_/A VGND VGND VPWR VPWR _34574_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25712_ _24849_/X _33318_/Q _25718_/S VGND VGND VPWR VPWR _25713_/A sky130_fd_sc_hd__mux2_1
X_29480_ _29480_/A VGND VGND VPWR VPWR _35014_/D sky130_fd_sc_hd__clkbuf_1
X_22924_ _22924_/A VGND VGND VPWR VPWR _32033_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26692_ _26761_/S VGND VGND VPWR VPWR _26711_/S sky130_fd_sc_hd__buf_4
XFILLER_217_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28431_ _28431_/A VGND VGND VPWR VPWR _34541_/D sky130_fd_sc_hd__clkbuf_1
X_25643_ _25643_/A VGND VGND VPWR VPWR _33285_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22855_ _22851_/X _22854_/X _22438_/A VGND VGND VPWR VPWR _22877_/A sky130_fd_sc_hd__o21ba_1
XFILLER_25_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28362_ _27813_/X _34509_/Q _28370_/S VGND VGND VPWR VPWR _28363_/A sky130_fd_sc_hd__mux2_1
X_21806_ _22512_/A VGND VGND VPWR VPWR _21806_/X sky130_fd_sc_hd__buf_6
X_22786_ _22782_/X _22785_/X _22471_/A VGND VGND VPWR VPWR _22787_/D sky130_fd_sc_hd__o21ba_1
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25574_ _25574_/A VGND VGND VPWR VPWR _33252_/D sky130_fd_sc_hd__clkbuf_1
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27313_ _34043_/Q _27149_/X _27317_/S VGND VGND VPWR VPWR _27314_/A sky130_fd_sc_hd__mux2_1
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24525_ _24525_/A VGND VGND VPWR VPWR _32789_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21737_ _32116_/Q _32308_/Q _32372_/Q _35892_/Q _21527_/X _21668_/X VGND VGND VPWR
+ VPWR _21737_/X sky130_fd_sc_hd__mux4_1
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28293_ _27711_/X _34476_/Q _28307_/S VGND VGND VPWR VPWR _28294_/A sky130_fd_sc_hd__mux2_1
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27244_ _34010_/Q _27047_/X _27254_/S VGND VGND VPWR VPWR _27245_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21668_ _22374_/A VGND VGND VPWR VPWR _21668_/X sky130_fd_sc_hd__clkbuf_4
X_24456_ _22980_/X _32756_/Q _24474_/S VGND VGND VPWR VPWR _24457_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20619_ _20661_/A VGND VGND VPWR VPWR _22582_/A sky130_fd_sc_hd__buf_12
X_23407_ _23407_/A VGND VGND VPWR VPWR _32214_/D sky130_fd_sc_hd__clkbuf_1
X_27175_ _33987_/Q _27174_/X _27187_/S VGND VGND VPWR VPWR _27176_/A sky130_fd_sc_hd__mux2_1
X_24387_ _23079_/X _32724_/Q _24389_/S VGND VGND VPWR VPWR _24388_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_1274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21599_ _35696_/Q _32204_/Q _35568_/Q _35504_/Q _21564_/X _21565_/X VGND VGND VPWR
+ VPWR _21599_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26126_ _24861_/X _33514_/Q _26144_/S VGND VGND VPWR VPWR _26127_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23338_ _32186_/Q _23261_/X _23359_/S VGND VGND VPWR VPWR _23339_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_798 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26057_ _26057_/A VGND VGND VPWR VPWR _33481_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23269_ _32162_/Q _23268_/X _23290_/S VGND VGND VPWR VPWR _23270_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_6_4__f_CLK clkbuf_5_2_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_4__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_25008_ _25008_/A VGND VGND VPWR VPWR _32986_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17830_ _33672_/Q _33608_/Q _33544_/Q _33480_/Q _17553_/X _17554_/X VGND VGND VPWR
+ VPWR _17830_/X sky130_fd_sc_hd__mux4_1
X_29816_ _29816_/A VGND VGND VPWR VPWR _35166_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17761_ _33414_/Q _33350_/Q _33286_/Q _33222_/Q _17480_/X _17481_/X VGND VGND VPWR
+ VPWR _17761_/X sky130_fd_sc_hd__mux4_1
X_29747_ _29795_/S VGND VGND VPWR VPWR _29766_/S sky130_fd_sc_hd__buf_4
XFILLER_19_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26959_ _26959_/A VGND VGND VPWR VPWR _33906_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19500_ _20206_/A VGND VGND VPWR VPWR _19500_/X sky130_fd_sc_hd__buf_6
X_16712_ _17910_/A VGND VGND VPWR VPWR _16712_/X sky130_fd_sc_hd__clkbuf_4
X_29678_ _35101_/Q _29351_/X _29682_/S VGND VGND VPWR VPWR _29679_/A sky130_fd_sc_hd__mux2_1
X_17692_ _33924_/Q _33860_/Q _33796_/Q _36100_/Q _17377_/X _17378_/X VGND VGND VPWR
+ VPWR _17692_/X sky130_fd_sc_hd__mux4_1
XFILLER_130_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19431_ _19153_/X _19429_/X _19430_/X _19156_/X VGND VGND VPWR VPWR _19431_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28629_ _28629_/A VGND VGND VPWR VPWR _34635_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_207_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16643_ _16361_/X _16639_/X _16642_/X _16365_/X VGND VGND VPWR VPWR _16643_/X sky130_fd_sc_hd__a22o_1
XFILLER_74_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31640_ _31640_/A VGND VGND VPWR VPWR _36030_/D sky130_fd_sc_hd__clkbuf_1
X_19362_ _20286_/A VGND VGND VPWR VPWR _19362_/X sky130_fd_sc_hd__buf_4
X_16574_ _17986_/A VGND VGND VPWR VPWR _16574_/X sky130_fd_sc_hd__buf_4
XFILLER_90_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18313_ _18301_/X _18304_/X _18307_/X _18312_/X VGND VGND VPWR VPWR _18313_/X sky130_fd_sc_hd__a22o_1
XFILLER_43_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31571_ _27667_/X _35998_/Q _31573_/S VGND VGND VPWR VPWR _31572_/A sky130_fd_sc_hd__mux2_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19293_ _20133_/A VGND VGND VPWR VPWR _19293_/X sky130_fd_sc_hd__buf_4
XFILLER_176_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33310_ _33821_/CLK _33310_/D VGND VGND VPWR VPWR _33310_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18244_ _34964_/Q _34900_/Q _34836_/Q _34772_/Q _16083_/X _16085_/X VGND VGND VPWR
+ VPWR _18244_/X sky130_fd_sc_hd__mux4_1
X_30522_ _35501_/Q _29401_/X _30534_/S VGND VGND VPWR VPWR _30523_/A sky130_fd_sc_hd__mux2_1
XFILLER_187_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_838 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34290_ _36143_/CLK _34290_/D VGND VGND VPWR VPWR _34290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33241_ _33753_/CLK _33241_/D VGND VGND VPWR VPWR _33241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18175_ _15981_/X _18173_/X _18174_/X _15991_/X VGND VGND VPWR VPWR _18175_/X sky130_fd_sc_hd__a22o_1
X_30453_ _30453_/A VGND VGND VPWR VPWR _35468_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17126_ _16846_/X _17124_/X _17125_/X _16851_/X VGND VGND VPWR VPWR _17126_/X sky130_fd_sc_hd__a22o_1
XFILLER_15_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33172_ _36052_/CLK _33172_/D VGND VGND VPWR VPWR _33172_/Q sky130_fd_sc_hd__dfxtp_1
X_30384_ _30384_/A VGND VGND VPWR VPWR _35435_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32123_ _35962_/CLK _32123_/D VGND VGND VPWR VPWR _32123_/Q sky130_fd_sc_hd__dfxtp_1
X_17057_ _16853_/X _17055_/X _17056_/X _16856_/X VGND VGND VPWR VPWR _17057_/X sky130_fd_sc_hd__a22o_1
XFILLER_48_1120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16008_ _16061_/A VGND VGND VPWR VPWR _17960_/A sky130_fd_sc_hd__buf_12
X_32054_ _35765_/CLK _32054_/D VGND VGND VPWR VPWR _32054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31005_ _31005_/A VGND VGND VPWR VPWR _35730_/D sky130_fd_sc_hd__clkbuf_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35813_ _35814_/CLK _35813_/D VGND VGND VPWR VPWR _35813_/Q sky130_fd_sc_hd__dfxtp_1
X_17959_ _17704_/X _17957_/X _17958_/X _17707_/X VGND VGND VPWR VPWR _17959_/X sky130_fd_sc_hd__a22o_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20970_ _20892_/X _20968_/X _20969_/X _20895_/X VGND VGND VPWR VPWR _20970_/X sky130_fd_sc_hd__a22o_1
X_35744_ _35810_/CLK _35744_/D VGND VGND VPWR VPWR _35744_/Q sky130_fd_sc_hd__dfxtp_1
X_32956_ _35451_/CLK _32956_/D VGND VGND VPWR VPWR _32956_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31907_ _31907_/A VGND VGND VPWR VPWR _36157_/D sky130_fd_sc_hd__clkbuf_1
X_19629_ _34425_/Q _36153_/Q _34297_/Q _34233_/Q _19529_/X _19530_/X VGND VGND VPWR
+ VPWR _19629_/X sky130_fd_sc_hd__mux4_1
X_35675_ _35804_/CLK _35675_/D VGND VGND VPWR VPWR _35675_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32887_ _32887_/CLK _32887_/D VGND VGND VPWR VPWR _32887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22640_ _34190_/Q _34126_/Q _34062_/Q _33998_/Q _22399_/X _22400_/X VGND VGND VPWR
+ VPWR _22640_/X sky130_fd_sc_hd__mux4_1
X_31838_ _31838_/A VGND VGND VPWR VPWR _36124_/D sky130_fd_sc_hd__clkbuf_1
X_34626_ _34626_/CLK _34626_/D VGND VGND VPWR VPWR _34626_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22571_ _22464_/X _22569_/X _22570_/X _22469_/X VGND VGND VPWR VPWR _22571_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_833 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34557_ _36152_/CLK _34557_/D VGND VGND VPWR VPWR _34557_/Q sky130_fd_sc_hd__dfxtp_1
X_31769_ _36092_/Q input32/X _31771_/S VGND VGND VPWR VPWR _31770_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21522_ _21518_/X _21521_/X _21379_/X VGND VGND VPWR VPWR _21548_/A sky130_fd_sc_hd__o21ba_1
X_24310_ _22965_/X _32687_/Q _24318_/S VGND VGND VPWR VPWR _24311_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25290_ _33119_/Q _23258_/X _25290_/S VGND VGND VPWR VPWR _25291_/A sky130_fd_sc_hd__mux2_1
X_33508_ _34151_/CLK _33508_/D VGND VGND VPWR VPWR _33508_/Q sky130_fd_sc_hd__dfxtp_1
X_34488_ _35193_/CLK _34488_/D VGND VGND VPWR VPWR _34488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24241_ _32656_/Q _23481_/X _24243_/S VGND VGND VPWR VPWR _24242_/A sky130_fd_sc_hd__mux2_1
X_36227_ _36229_/CLK _36227_/D VGND VGND VPWR VPWR _36227_/Q sky130_fd_sc_hd__dfxtp_1
X_33439_ _36191_/CLK _33439_/D VGND VGND VPWR VPWR _33439_/Q sky130_fd_sc_hd__dfxtp_1
X_21453_ _22512_/A VGND VGND VPWR VPWR _21453_/X sky130_fd_sc_hd__buf_4
XFILLER_147_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20404_ _20212_/X _20402_/X _20403_/X _20215_/X VGND VGND VPWR VPWR _20404_/X sky130_fd_sc_hd__a22o_1
XFILLER_193_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36158_ _36159_/CLK _36158_/D VGND VGND VPWR VPWR _36158_/Q sky130_fd_sc_hd__dfxtp_1
X_24172_ _32623_/Q _23316_/X _24180_/S VGND VGND VPWR VPWR _24173_/A sky130_fd_sc_hd__mux2_1
X_21384_ _32106_/Q _32298_/Q _32362_/Q _35882_/Q _21174_/X _21315_/X VGND VGND VPWR
+ VPWR _21384_/X sky130_fd_sc_hd__mux4_1
X_23123_ _22934_/X _32101_/Q _23131_/S VGND VGND VPWR VPWR _23124_/A sky130_fd_sc_hd__mux2_1
X_20335_ _20164_/X _20333_/X _20334_/X _20169_/X VGND VGND VPWR VPWR _20335_/X sky130_fd_sc_hd__a22o_1
X_35109_ _35168_/CLK _35109_/D VGND VGND VPWR VPWR _35109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36089_ _36090_/CLK _36089_/D VGND VGND VPWR VPWR _36089_/Q sky130_fd_sc_hd__dfxtp_1
X_28980_ _28980_/A VGND VGND VPWR VPWR _34800_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27931_ _27931_/A VGND VGND VPWR VPWR _34304_/D sky130_fd_sc_hd__clkbuf_1
X_23054_ _23054_/A VGND VGND VPWR VPWR _32075_/D sky130_fd_sc_hd__clkbuf_1
X_20266_ _34699_/Q _34635_/Q _34571_/Q _34507_/Q _19945_/X _19946_/X VGND VGND VPWR
+ VPWR _20266_/X sky130_fd_sc_hd__mux4_1
XFILLER_116_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22005_ _33660_/Q _33596_/Q _33532_/Q _33468_/Q _21800_/X _21801_/X VGND VGND VPWR
+ VPWR _22005_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_963 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27862_ _27973_/S VGND VGND VPWR VPWR _27881_/S sky130_fd_sc_hd__buf_4
XFILLER_49_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_248_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20197_ _35209_/Q _35145_/Q _35081_/Q _32265_/Q _20016_/X _20017_/X VGND VGND VPWR
+ VPWR _20197_/X sky130_fd_sc_hd__mux4_1
XTAP_5326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29601_ _29601_/A VGND VGND VPWR VPWR _35064_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26813_ _33837_/Q _23302_/X _26825_/S VGND VGND VPWR VPWR _26814_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27793_ _27793_/A VGND VGND VPWR VPWR _34246_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29532_ _29532_/A VGND VGND VPWR VPWR _35031_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26744_ _26744_/A VGND VGND VPWR VPWR _33804_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23956_ _23956_/A VGND VGND VPWR VPWR _32522_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29463_ input38/X VGND VGND VPWR VPWR _29463_/X sky130_fd_sc_hd__clkbuf_4
X_22907_ _22906_/X _32028_/Q _22916_/S VGND VGND VPWR VPWR _22908_/A sky130_fd_sc_hd__mux2_1
XFILLER_244_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26675_ _26675_/A VGND VGND VPWR VPWR _33771_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_229_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23887_ _23977_/S VGND VGND VPWR VPWR _23906_/S sky130_fd_sc_hd__buf_4
XFILLER_217_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28414_ _28414_/A VGND VGND VPWR VPWR _34533_/D sky130_fd_sc_hd__clkbuf_1
X_25626_ _25626_/A VGND VGND VPWR VPWR _33277_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22838_ _20601_/X _22836_/X _22837_/X _20607_/X VGND VGND VPWR VPWR _22838_/X sky130_fd_sc_hd__a22o_1
X_29394_ _29394_/A VGND VGND VPWR VPWR _34986_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_227_1040 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28345_ _27788_/X _34501_/Q _28349_/S VGND VGND VPWR VPWR _28346_/A sky130_fd_sc_hd__mux2_1
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25557_ _25557_/A VGND VGND VPWR VPWR _33244_/D sky130_fd_sc_hd__clkbuf_1
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22769_ _32146_/Q _32338_/Q _32402_/Q _35922_/Q _22586_/X _21611_/A VGND VGND VPWR
+ VPWR _22769_/X sky130_fd_sc_hd__mux4_1
XFILLER_24_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24508_ _23058_/X _32781_/Q _24516_/S VGND VGND VPWR VPWR _24509_/A sky130_fd_sc_hd__mux2_1
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16290_ _16030_/X _16286_/X _16289_/X _16041_/X VGND VGND VPWR VPWR _16290_/X sky130_fd_sc_hd__a22o_1
X_28276_ _27686_/X _34468_/Q _28286_/S VGND VGND VPWR VPWR _28277_/A sky130_fd_sc_hd__mux2_1
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25488_ _24917_/X _33212_/Q _25490_/S VGND VGND VPWR VPWR _25489_/A sky130_fd_sc_hd__mux2_1
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27227_ _34004_/Q _27226_/X _27230_/S VGND VGND VPWR VPWR _27228_/A sky130_fd_sc_hd__mux2_1
XFILLER_200_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24439_ _22956_/X _32748_/Q _24453_/S VGND VGND VPWR VPWR _24440_/A sky130_fd_sc_hd__mux2_1
XFILLER_205_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27158_ input35/X VGND VGND VPWR VPWR _27158_/X sky130_fd_sc_hd__buf_4
XFILLER_125_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26109_ _24837_/X _33506_/Q _26123_/S VGND VGND VPWR VPWR _26110_/A sky130_fd_sc_hd__mux2_1
X_19980_ _35203_/Q _35139_/Q _35075_/Q _32259_/Q _19663_/X _19664_/X VGND VGND VPWR
+ VPWR _19980_/X sky130_fd_sc_hd__mux4_1
XFILLER_181_863 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27089_ _27089_/A VGND VGND VPWR VPWR _33959_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18931_ _18793_/X _18929_/X _18930_/X _18798_/X VGND VGND VPWR VPWR _18931_/X sky130_fd_sc_hd__a22o_1
XFILLER_180_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18862_ _18862_/A VGND VGND VPWR VPWR _32419_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17813_ _17809_/X _17812_/X _17493_/X _17494_/X VGND VGND VPWR VPWR _17828_/B sky130_fd_sc_hd__o211a_1
XFILLER_122_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18793_ _20205_/A VGND VGND VPWR VPWR _18793_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_212_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32810_ _32914_/CLK _32810_/D VGND VGND VPWR VPWR _32810_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_248_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17744_ _17704_/X _17742_/X _17743_/X _17707_/X VGND VGND VPWR VPWR _17744_/X sky130_fd_sc_hd__a22o_1
XFILLER_236_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33790_ _35711_/CLK _33790_/D VGND VGND VPWR VPWR _33790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32741_ _32869_/CLK _32741_/D VGND VGND VPWR VPWR _32741_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17675_ _35459_/Q _35395_/Q _35331_/Q _35267_/Q _17607_/X _17608_/X VGND VGND VPWR
+ VPWR _17675_/X sky130_fd_sc_hd__mux4_1
XFILLER_235_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_247_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19414_ _19410_/X _19413_/X _19098_/X VGND VGND VPWR VPWR _19422_/C sky130_fd_sc_hd__o21ba_1
X_35460_ _35843_/CLK _35460_/D VGND VGND VPWR VPWR _35460_/Q sky130_fd_sc_hd__dfxtp_1
X_16626_ _16622_/X _16625_/X _16459_/X VGND VGND VPWR VPWR _16627_/D sky130_fd_sc_hd__o21ba_1
X_32672_ _33119_/CLK _32672_/D VGND VGND VPWR VPWR _32672_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34411_ _36141_/CLK _34411_/D VGND VGND VPWR VPWR _34411_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_5_10_0_CLK clkbuf_5_9_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_10_0_CLK/X sky130_fd_sc_hd__clkbuf_8
X_19345_ _19100_/X _19343_/X _19344_/X _19103_/X VGND VGND VPWR VPWR _19345_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31623_ _31623_/A VGND VGND VPWR VPWR _36022_/D sky130_fd_sc_hd__clkbuf_1
X_35391_ _35456_/CLK _35391_/D VGND VGND VPWR VPWR _35391_/Q sky130_fd_sc_hd__dfxtp_1
X_16557_ _34403_/Q _36131_/Q _34275_/Q _34211_/Q _16523_/X _16524_/X VGND VGND VPWR
+ VPWR _16557_/X sky130_fd_sc_hd__mux4_1
XFILLER_210_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34342_ _35620_/CLK _34342_/D VGND VGND VPWR VPWR _34342_/Q sky130_fd_sc_hd__dfxtp_1
X_31554_ _31686_/S VGND VGND VPWR VPWR _31573_/S sky130_fd_sc_hd__clkbuf_8
X_19276_ _34415_/Q _36143_/Q _34287_/Q _34223_/Q _19176_/X _19177_/X VGND VGND VPWR
+ VPWR _19276_/X sky130_fd_sc_hd__mux4_1
XFILLER_203_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16488_ _34913_/Q _34849_/Q _34785_/Q _34721_/Q _16454_/X _16455_/X VGND VGND VPWR
+ VPWR _16488_/X sky130_fd_sc_hd__mux4_1
XFILLER_143_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18227_ _33172_/Q _36052_/Q _33044_/Q _32980_/Q _16032_/X _17161_/A VGND VGND VPWR
+ VPWR _18227_/X sky130_fd_sc_hd__mux4_1
X_30505_ _35493_/Q _29376_/X _30513_/S VGND VGND VPWR VPWR _30506_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34273_ _36128_/CLK _34273_/D VGND VGND VPWR VPWR _34273_/Q sky130_fd_sc_hd__dfxtp_1
X_31485_ _27739_/X _35957_/Q _31501_/S VGND VGND VPWR VPWR _31486_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_5_25_0_CLK clkbuf_2_3_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_25_0_CLK/X sky130_fd_sc_hd__clkbuf_8
X_36012_ _36141_/CLK _36012_/D VGND VGND VPWR VPWR _36012_/Q sky130_fd_sc_hd__dfxtp_1
X_33224_ _33420_/CLK _33224_/D VGND VGND VPWR VPWR _33224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30436_ _30436_/A VGND VGND VPWR VPWR _35460_/D sky130_fd_sc_hd__clkbuf_1
X_18158_ _18158_/A VGND VGND VPWR VPWR _32017_/D sky130_fd_sc_hd__clkbuf_1
X_17109_ _35635_/Q _34995_/Q _34355_/Q _33715_/Q _16791_/X _16792_/X VGND VGND VPWR
+ VPWR _17109_/X sky130_fd_sc_hd__mux4_1
X_33155_ _35779_/CLK _33155_/D VGND VGND VPWR VPWR _33155_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18089_ _18085_/X _18088_/X _17857_/X VGND VGND VPWR VPWR _18097_/C sky130_fd_sc_hd__o21ba_1
XFILLER_132_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30367_ _30367_/A VGND VGND VPWR VPWR _35427_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_176_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20120_ _20116_/X _20119_/X _19804_/X VGND VGND VPWR VPWR _20128_/C sky130_fd_sc_hd__o21ba_1
XFILLER_144_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32106_ _35949_/CLK _32106_/D VGND VGND VPWR VPWR _32106_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33086_ _35454_/CLK _33086_/D VGND VGND VPWR VPWR _33086_/Q sky130_fd_sc_hd__dfxtp_1
X_30298_ _35395_/Q _29469_/X _30306_/S VGND VGND VPWR VPWR _30299_/A sky130_fd_sc_hd__mux2_1
X_20051_ _19806_/X _20049_/X _20050_/X _19809_/X VGND VGND VPWR VPWR _20051_/X sky130_fd_sc_hd__a22o_1
X_32037_ _35814_/CLK _32037_/D VGND VGND VPWR VPWR _32037_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23810_ _23810_/A VGND VGND VPWR VPWR _32390_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24790_ _23076_/X _32915_/Q _24794_/S VGND VGND VPWR VPWR _24791_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33988_ _34180_/CLK _33988_/D VGND VGND VPWR VPWR _33988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35727_ _35727_/CLK _35727_/D VGND VGND VPWR VPWR _35727_/Q sky130_fd_sc_hd__dfxtp_1
X_20953_ _22505_/A VGND VGND VPWR VPWR _20953_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_38_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23741_ _23741_/A VGND VGND VPWR VPWR _32357_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_226_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32939_ _36010_/CLK _32939_/D VGND VGND VPWR VPWR _32939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26460_ _33672_/Q _23453_/X _26478_/S VGND VGND VPWR VPWR _26461_/A sky130_fd_sc_hd__mux2_1
XFILLER_187_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35658_ _35658_/CLK _35658_/D VGND VGND VPWR VPWR _35658_/Q sky130_fd_sc_hd__dfxtp_1
X_20884_ _33116_/Q _35996_/Q _32988_/Q _32924_/Q _20624_/X _20625_/X VGND VGND VPWR
+ VPWR _20884_/X sky130_fd_sc_hd__mux4_1
X_23672_ _23672_/A VGND VGND VPWR VPWR _32326_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25411_ _24803_/X _33175_/Q _25427_/S VGND VGND VPWR VPWR _25412_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22623_ _35725_/Q _32236_/Q _35597_/Q _35533_/Q _20593_/X _20595_/X VGND VGND VPWR
+ VPWR _22623_/X sky130_fd_sc_hd__mux4_1
X_34609_ _34611_/CLK _34609_/D VGND VGND VPWR VPWR _34609_/Q sky130_fd_sc_hd__dfxtp_1
X_26391_ _26391_/A VGND VGND VPWR VPWR _33639_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35589_ _35718_/CLK _35589_/D VGND VGND VPWR VPWR _35589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28130_ _27670_/X _34399_/Q _28130_/S VGND VGND VPWR VPWR _28131_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22554_ _32907_/Q _32843_/Q _32779_/Q _32715_/Q _22299_/X _22300_/X VGND VGND VPWR
+ VPWR _22554_/X sky130_fd_sc_hd__mux4_1
X_25342_ _25342_/A VGND VGND VPWR VPWR _33143_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21505_ _21250_/X _21503_/X _21504_/X _21253_/X VGND VGND VPWR VPWR _21505_/X sky130_fd_sc_hd__a22o_1
X_28061_ _34366_/Q _27158_/X _28079_/S VGND VGND VPWR VPWR _28062_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25273_ _25273_/A VGND VGND VPWR VPWR _33110_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22485_ _32137_/Q _32329_/Q _32393_/Q _35913_/Q _22233_/X _22374_/X VGND VGND VPWR
+ VPWR _22485_/X sky130_fd_sc_hd__mux4_1
XFILLER_195_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27012_ _27012_/A VGND VGND VPWR VPWR _33931_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24224_ _24251_/S VGND VGND VPWR VPWR _24243_/S sky130_fd_sc_hd__buf_4
X_21436_ _21432_/X _21435_/X _21398_/X VGND VGND VPWR VPWR _21444_/C sky130_fd_sc_hd__o21ba_1
XFILLER_107_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_17__f_CLK clkbuf_5_8_0_CLK/X VGND VGND VPWR VPWR clkbuf_leaf_99_CLK/A sky130_fd_sc_hd__clkbuf_16
X_24155_ _32615_/Q _23283_/X _24159_/S VGND VGND VPWR VPWR _24156_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_190_CLK clkbuf_6_48__f_CLK/X VGND VGND VPWR VPWR _32655_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_135_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21367_ _21052_/X _21365_/X _21366_/X _21057_/X VGND VGND VPWR VPWR _21367_/X sky130_fd_sc_hd__a22o_1
XFILLER_107_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23106_ _22909_/X _32093_/Q _23110_/S VGND VGND VPWR VPWR _23107_/A sky130_fd_sc_hd__mux2_1
X_20318_ _20065_/X _20316_/X _20317_/X _20071_/X VGND VGND VPWR VPWR _20318_/X sky130_fd_sc_hd__a22o_1
XFILLER_190_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24086_ _24113_/S VGND VGND VPWR VPWR _24105_/S sky130_fd_sc_hd__buf_4
XFILLER_122_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28963_ _28963_/A VGND VGND VPWR VPWR _34792_/D sky130_fd_sc_hd__clkbuf_1
X_21298_ _21298_/A VGND VGND VPWR VPWR _36199_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23037_ _23036_/X _32070_/Q _23040_/S VGND VGND VPWR VPWR _23038_/A sky130_fd_sc_hd__mux2_1
X_27914_ _27914_/A VGND VGND VPWR VPWR _34296_/D sky130_fd_sc_hd__clkbuf_1
X_20249_ _20245_/X _20248_/X _20138_/X VGND VGND VPWR VPWR _20273_/A sky130_fd_sc_hd__o21ba_2
XFILLER_67_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28894_ _28921_/S VGND VGND VPWR VPWR _28913_/S sky130_fd_sc_hd__buf_4
XTAP_5101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27845_ _27845_/A VGND VGND VPWR VPWR _34263_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_847 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27776_ input38/X VGND VGND VPWR VPWR _27776_/X sky130_fd_sc_hd__buf_2
XTAP_4455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24988_ input58/X VGND VGND VPWR VPWR _24988_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29515_ input57/X VGND VGND VPWR VPWR _29515_/X sky130_fd_sc_hd__buf_2
XTAP_4477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26727_ _26727_/A VGND VGND VPWR VPWR _33796_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23939_ _23939_/A VGND VGND VPWR VPWR _32514_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29446_ _29446_/A VGND VGND VPWR VPWR _35003_/D sky130_fd_sc_hd__clkbuf_1
X_17460_ _17456_/X _17459_/X _17140_/X _17141_/X VGND VGND VPWR VPWR _17475_/B sky130_fd_sc_hd__o211a_1
XFILLER_205_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26658_ _26658_/A VGND VGND VPWR VPWR _33763_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16411_ _16078_/X _16409_/X _16410_/X _16088_/X VGND VGND VPWR VPWR _16411_/X sky130_fd_sc_hd__a22o_1
X_25609_ _24896_/X _33269_/Q _25625_/S VGND VGND VPWR VPWR _25610_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29377_ _34981_/Q _29376_/X _29389_/S VGND VGND VPWR VPWR _29378_/A sky130_fd_sc_hd__mux2_1
X_17391_ _17351_/X _17389_/X _17390_/X _17354_/X VGND VGND VPWR VPWR _17391_/X sky130_fd_sc_hd__a22o_1
XFILLER_242_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26589_ _24945_/X _33733_/Q _26593_/S VGND VGND VPWR VPWR _26590_/A sky130_fd_sc_hd__mux2_1
XFILLER_246_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19130_ _35691_/Q _32199_/Q _35563_/Q _35499_/Q _18911_/X _18912_/X VGND VGND VPWR
+ VPWR _19130_/X sky130_fd_sc_hd__mux4_1
X_16342_ _16091_/X _16340_/X _16341_/X _16101_/X VGND VGND VPWR VPWR _16342_/X sky130_fd_sc_hd__a22o_1
X_28328_ _27763_/X _34493_/Q _28328_/S VGND VGND VPWR VPWR _28329_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19061_ _19057_/X _19060_/X _18745_/X VGND VGND VPWR VPWR _19069_/C sky130_fd_sc_hd__o21ba_1
X_16273_ _16269_/X _16272_/X _16104_/X VGND VGND VPWR VPWR _16274_/D sky130_fd_sc_hd__o21ba_1
X_28259_ _27661_/X _34460_/Q _28265_/S VGND VGND VPWR VPWR _28260_/A sky130_fd_sc_hd__mux2_1
X_18012_ _33421_/Q _33357_/Q _33293_/Q _33229_/Q _17833_/X _17834_/X VGND VGND VPWR
+ VPWR _18012_/X sky130_fd_sc_hd__mux4_1
XFILLER_16_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31270_ _31270_/A VGND VGND VPWR VPWR _35855_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30221_ _30221_/A VGND VGND VPWR VPWR _35358_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_181_CLK clkbuf_6_27__f_CLK/X VGND VGND VPWR VPWR _35599_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_181_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30152_ _30200_/S VGND VGND VPWR VPWR _30171_/S sky130_fd_sc_hd__buf_6
X_19963_ _32643_/Q _32579_/Q _32515_/Q _35971_/Q _19929_/X _19713_/X VGND VGND VPWR
+ VPWR _19963_/X sky130_fd_sc_hd__mux4_1
XFILLER_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18914_ _35621_/Q _34981_/Q _34341_/Q _33701_/Q _18738_/X _18739_/X VGND VGND VPWR
+ VPWR _18914_/X sky130_fd_sc_hd__mux4_1
XTAP_7070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34960_ _34961_/CLK _34960_/D VGND VGND VPWR VPWR _34960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30083_ _35293_/Q _29351_/X _30087_/S VGND VGND VPWR VPWR _30084_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19894_ _33921_/Q _33857_/Q _33793_/Q _36097_/Q _19677_/X _19678_/X VGND VGND VPWR
+ VPWR _19894_/X sky130_fd_sc_hd__mux4_1
XTAP_7092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_214_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33911_ _33911_/CLK _33911_/D VGND VGND VPWR VPWR _33911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18845_ _35683_/Q _32190_/Q _35555_/Q _35491_/Q _18558_/X _18559_/X VGND VGND VPWR
+ VPWR _18845_/X sky130_fd_sc_hd__mux4_1
X_34891_ _34957_/CLK _34891_/D VGND VGND VPWR VPWR _34891_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_966 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18776_ _18772_/X _18775_/X _18734_/X _18735_/X VGND VGND VPWR VPWR _18791_/B sky130_fd_sc_hd__o211a_1
X_33842_ _34099_/CLK _33842_/D VGND VGND VPWR VPWR _33842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_212_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15988_ _33622_/Q _33558_/Q _33494_/Q _33430_/Q _15984_/X _15987_/X VGND VGND VPWR
+ VPWR _15988_/X sky130_fd_sc_hd__mux4_1
XFILLER_94_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17727_ _34181_/Q _34117_/Q _34053_/Q _33989_/Q _17446_/X _17447_/X VGND VGND VPWR
+ VPWR _17727_/X sky130_fd_sc_hd__mux4_1
X_33773_ _34093_/CLK _33773_/D VGND VGND VPWR VPWR _33773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30985_ _30985_/A VGND VGND VPWR VPWR _35720_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_208_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35512_ _35768_/CLK _35512_/D VGND VGND VPWR VPWR _35512_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_235_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17658_ _17552_/X _17656_/X _17657_/X _17557_/X VGND VGND VPWR VPWR _17658_/X sky130_fd_sc_hd__a22o_1
X_32724_ _32869_/CLK _32724_/D VGND VGND VPWR VPWR _32724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16609_ _16361_/X _16607_/X _16608_/X _16365_/X VGND VGND VPWR VPWR _16609_/X sky130_fd_sc_hd__a22o_1
XFILLER_211_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32655_ _32655_/CLK _32655_/D VGND VGND VPWR VPWR _32655_/Q sky130_fd_sc_hd__dfxtp_1
X_35443_ _35764_/CLK _35443_/D VGND VGND VPWR VPWR _35443_/Q sky130_fd_sc_hd__dfxtp_1
X_17589_ _17589_/A VGND VGND VPWR VPWR _32000_/D sky130_fd_sc_hd__buf_4
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19328_ _19322_/X _19327_/X _19079_/X VGND VGND VPWR VPWR _19350_/A sky130_fd_sc_hd__o21ba_1
X_31606_ _31606_/A VGND VGND VPWR VPWR _36014_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32586_ _35978_/CLK _32586_/D VGND VGND VPWR VPWR _32586_/Q sky130_fd_sc_hd__dfxtp_1
X_35374_ _35438_/CLK _35374_/D VGND VGND VPWR VPWR _35374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34325_ _36181_/CLK _34325_/D VGND VGND VPWR VPWR _34325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31537_ _27816_/X _35982_/Q _31543_/S VGND VGND VPWR VPWR _31538_/A sky130_fd_sc_hd__mux2_1
X_19259_ _19006_/X _19257_/X _19258_/X _19012_/X VGND VGND VPWR VPWR _19259_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34256_ _36176_/CLK _34256_/D VGND VGND VPWR VPWR _34256_/Q sky130_fd_sc_hd__dfxtp_1
X_22270_ _22399_/A VGND VGND VPWR VPWR _22270_/X sky130_fd_sc_hd__buf_4
X_31468_ _27714_/X _35949_/Q _31480_/S VGND VGND VPWR VPWR _31469_/A sky130_fd_sc_hd__mux2_1
XFILLER_191_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33207_ _36087_/CLK _33207_/D VGND VGND VPWR VPWR _33207_/Q sky130_fd_sc_hd__dfxtp_1
X_21221_ _35173_/Q _35109_/Q _35045_/Q _32165_/Q _20904_/X _20905_/X VGND VGND VPWR
+ VPWR _21221_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30419_ _30419_/A VGND VGND VPWR VPWR _35452_/D sky130_fd_sc_hd__clkbuf_1
X_34187_ _34187_/CLK _34187_/D VGND VGND VPWR VPWR _34187_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_172_CLK clkbuf_6_28__f_CLK/X VGND VGND VPWR VPWR _35865_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_117_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31399_ _31399_/A VGND VGND VPWR VPWR _35916_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21152_ _20897_/X _21150_/X _21151_/X _20900_/X VGND VGND VPWR VPWR _21152_/X sky130_fd_sc_hd__a22o_1
X_33138_ _36020_/CLK _33138_/D VGND VGND VPWR VPWR _33138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20103_ _33415_/Q _33351_/Q _33287_/Q _33223_/Q _19780_/X _19781_/X VGND VGND VPWR
+ VPWR _20103_/X sky130_fd_sc_hd__mux4_1
XFILLER_137_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25960_ _25960_/A VGND VGND VPWR VPWR _33435_/D sky130_fd_sc_hd__clkbuf_1
X_33069_ _35822_/CLK _33069_/D VGND VGND VPWR VPWR _33069_/Q sky130_fd_sc_hd__dfxtp_1
X_21083_ _21079_/X _21082_/X _21045_/X VGND VGND VPWR VPWR _21091_/C sky130_fd_sc_hd__o21ba_1
XFILLER_101_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20034_ _20028_/X _20033_/X _19785_/X VGND VGND VPWR VPWR _20056_/A sky130_fd_sc_hd__o21ba_2
XFILLER_119_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24911_ input30/X VGND VGND VPWR VPWR _24911_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_113_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25891_ _24914_/X _33403_/Q _25895_/S VGND VGND VPWR VPWR _25892_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27630_ _27630_/A VGND VGND VPWR VPWR _34193_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24842_ _24842_/A VGND VGND VPWR VPWR _32931_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27561_ _27561_/A VGND VGND VPWR VPWR _34160_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24773_ _24773_/A VGND VGND VPWR VPWR _32906_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21985_ _32123_/Q _32315_/Q _32379_/Q _35899_/Q _21880_/X _21668_/X VGND VGND VPWR
+ VPWR _21985_/X sky130_fd_sc_hd__mux4_1
X_29300_ _34952_/Q _27189_/X _29318_/S VGND VGND VPWR VPWR _29301_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26512_ _24830_/X _33696_/Q _26530_/S VGND VGND VPWR VPWR _26513_/A sky130_fd_sc_hd__mux2_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23724_ _23724_/A VGND VGND VPWR VPWR _32349_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27492_ _34128_/Q _27214_/X _27494_/S VGND VGND VPWR VPWR _27493_/A sky130_fd_sc_hd__mux2_1
X_20936_ _20932_/X _20935_/X _20675_/X VGND VGND VPWR VPWR _20944_/C sky130_fd_sc_hd__o21ba_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29231_ _29231_/A VGND VGND VPWR VPWR _34919_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26443_ _33664_/Q _23429_/X _26457_/S VGND VGND VPWR VPWR _26444_/A sky130_fd_sc_hd__mux2_1
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20867_ _34651_/Q _34587_/Q _34523_/Q _34459_/Q _20833_/X _20834_/X VGND VGND VPWR
+ VPWR _20867_/X sky130_fd_sc_hd__mux4_1
X_23655_ _23011_/X _32318_/Q _23673_/S VGND VGND VPWR VPWR _23656_/A sky130_fd_sc_hd__mux2_1
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_900 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22606_ _22602_/X _22605_/X _22471_/X VGND VGND VPWR VPWR _22607_/D sky130_fd_sc_hd__o21ba_1
X_29162_ _34887_/Q _27186_/X _29162_/S VGND VGND VPWR VPWR _29163_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_944 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26374_ _26374_/A VGND VGND VPWR VPWR _33631_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20798_ _33049_/Q _32025_/Q _35801_/Q _35737_/Q _20667_/X _20669_/X VGND VGND VPWR
+ VPWR _20798_/X sky130_fd_sc_hd__mux4_1
XFILLER_179_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23586_ _23586_/A VGND VGND VPWR VPWR _32285_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28113_ _28113_/A VGND VGND VPWR VPWR _34390_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25325_ _25325_/A VGND VGND VPWR VPWR _33135_/D sky130_fd_sc_hd__clkbuf_1
X_22537_ _34442_/Q _36170_/Q _34314_/Q _34250_/Q _22535_/X _22536_/X VGND VGND VPWR
+ VPWR _22537_/X sky130_fd_sc_hd__mux4_1
XFILLER_183_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29093_ _34854_/Q _27084_/X _29099_/S VGND VGND VPWR VPWR _29094_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28044_ _34358_/Q _27134_/X _28058_/S VGND VGND VPWR VPWR _28045_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25256_ _25256_/A VGND VGND VPWR VPWR _33103_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_1071 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22468_ _34952_/Q _34888_/Q _34824_/Q _34760_/Q _22466_/X _22467_/X VGND VGND VPWR
+ VPWR _22468_/X sky130_fd_sc_hd__mux4_1
XFILLER_154_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24207_ _24207_/A VGND VGND VPWR VPWR _32639_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_163_CLK clkbuf_6_30__f_CLK/X VGND VGND VPWR VPWR _34705_/CLK sky130_fd_sc_hd__clkbuf_16
X_21419_ _33387_/Q _33323_/Q _33259_/Q _33195_/Q _21374_/X _21375_/X VGND VGND VPWR
+ VPWR _21419_/X sky130_fd_sc_hd__mux4_1
X_22399_ _22399_/A VGND VGND VPWR VPWR _22399_/X sky130_fd_sc_hd__buf_4
X_25187_ _25187_/A VGND VGND VPWR VPWR _33070_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24138_ _32607_/Q _23258_/X _24138_/S VGND VGND VPWR VPWR _24139_/A sky130_fd_sc_hd__mux2_1
X_29995_ _29995_/A VGND VGND VPWR VPWR _35251_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_1148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16960_ _32111_/Q _32303_/Q _32367_/Q _35887_/Q _16927_/X _16715_/X VGND VGND VPWR
+ VPWR _16960_/X sky130_fd_sc_hd__mux4_1
X_24069_ _24069_/A VGND VGND VPWR VPWR _32575_/D sky130_fd_sc_hd__clkbuf_1
X_28946_ _34784_/Q _27065_/X _28964_/S VGND VGND VPWR VPWR _28947_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28877_ _28877_/A VGND VGND VPWR VPWR _34751_/D sky130_fd_sc_hd__clkbuf_1
X_16891_ _32621_/Q _32557_/Q _32493_/Q _35949_/Q _16570_/X _16707_/X VGND VGND VPWR
+ VPWR _16891_/X sky130_fd_sc_hd__mux4_1
XFILLER_131_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18630_ _35677_/Q _32183_/Q _35549_/Q _35485_/Q _18558_/X _18559_/X VGND VGND VPWR
+ VPWR _18630_/X sky130_fd_sc_hd__mux4_1
X_27828_ input57/X VGND VGND VPWR VPWR _27828_/X sky130_fd_sc_hd__clkbuf_4
XTAP_4230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18561_ _35611_/Q _34971_/Q _34331_/Q _33691_/Q _18353_/X _18355_/X VGND VGND VPWR
+ VPWR _18561_/X sky130_fd_sc_hd__mux4_1
XTAP_4274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_246_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27759_ _27759_/A VGND VGND VPWR VPWR _34235_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17512_ _34430_/Q _36158_/Q _34302_/Q _34238_/Q _17229_/X _17230_/X VGND VGND VPWR
+ VPWR _17512_/X sky130_fd_sc_hd__mux4_1
XTAP_3562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18492_ _35673_/Q _32179_/Q _35545_/Q _35481_/Q _18349_/X _18350_/X VGND VGND VPWR
+ VPWR _18492_/X sky130_fd_sc_hd__mux4_1
XTAP_3584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30770_ _30770_/A VGND VGND VPWR VPWR _35618_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29429_ input26/X VGND VGND VPWR VPWR _29429_/X sky130_fd_sc_hd__buf_2
XFILLER_32_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17443_ _17443_/A _17443_/B _17443_/C _17443_/D VGND VGND VPWR VPWR _17444_/A sky130_fd_sc_hd__or4_4
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32440_ _33895_/CLK _32440_/D VGND VGND VPWR VPWR _32440_/Q sky130_fd_sc_hd__dfxtp_1
X_17374_ _34171_/Q _34107_/Q _34043_/Q _33979_/Q _17093_/X _17094_/X VGND VGND VPWR
+ VPWR _17374_/X sky130_fd_sc_hd__mux4_1
XFILLER_158_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19113_ _19104_/X _19111_/X _19112_/X VGND VGND VPWR VPWR _19114_/D sky130_fd_sc_hd__o21ba_1
XFILLER_158_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16325_ _16018_/X _16323_/X _16324_/X _16027_/X VGND VGND VPWR VPWR _16325_/X sky130_fd_sc_hd__a22o_1
XFILLER_229_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32371_ _35955_/CLK _32371_/D VGND VGND VPWR VPWR _32371_/Q sky130_fd_sc_hd__dfxtp_1
X_34110_ _34174_/CLK _34110_/D VGND VGND VPWR VPWR _34110_/Q sky130_fd_sc_hd__dfxtp_1
X_19044_ _33385_/Q _33321_/Q _33257_/Q _33193_/Q _18721_/X _18722_/X VGND VGND VPWR
+ VPWR _19044_/X sky130_fd_sc_hd__mux4_1
XFILLER_12_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31322_ _27698_/X _35880_/Q _31324_/S VGND VGND VPWR VPWR _31323_/A sky130_fd_sc_hd__mux2_1
X_35090_ _35730_/CLK _35090_/D VGND VGND VPWR VPWR _35090_/Q sky130_fd_sc_hd__dfxtp_1
X_16256_ _16030_/X _16254_/X _16255_/X _16041_/X VGND VGND VPWR VPWR _16256_/X sky130_fd_sc_hd__a22o_1
XFILLER_127_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34041_ _35641_/CLK _34041_/D VGND VGND VPWR VPWR _34041_/Q sky130_fd_sc_hd__dfxtp_1
X_31253_ _31253_/A VGND VGND VPWR VPWR _35847_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_154_CLK clkbuf_6_31__f_CLK/X VGND VGND VPWR VPWR _33875_/CLK sky130_fd_sc_hd__clkbuf_16
X_16187_ _16018_/X _16185_/X _16186_/X _16027_/X VGND VGND VPWR VPWR _16187_/X sky130_fd_sc_hd__a22o_1
Xoutput205 _36238_/Q VGND VGND VPWR VPWR D2[56] sky130_fd_sc_hd__buf_2
XFILLER_103_1294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput216 _36190_/Q VGND VGND VPWR VPWR D2[8] sky130_fd_sc_hd__buf_2
X_30204_ _35350_/Q _29328_/X _30222_/S VGND VGND VPWR VPWR _30205_/A sky130_fd_sc_hd__mux2_1
Xoutput227 _32424_/Q VGND VGND VPWR VPWR D3[18] sky130_fd_sc_hd__buf_2
Xoutput238 _32434_/Q VGND VGND VPWR VPWR D3[28] sky130_fd_sc_hd__buf_2
Xoutput249 _32444_/Q VGND VGND VPWR VPWR D3[38] sky130_fd_sc_hd__buf_2
X_31184_ _31184_/A VGND VGND VPWR VPWR _35814_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_63__f_CLK clkbuf_5_31_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_63__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_30135_ _30135_/A VGND VGND VPWR VPWR _35317_/D sky130_fd_sc_hd__clkbuf_1
X_19946_ _20299_/A VGND VGND VPWR VPWR _19946_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_138_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35992_ _35992_/CLK _35992_/D VGND VGND VPWR VPWR _35992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34943_ _36161_/CLK _34943_/D VGND VGND VPWR VPWR _34943_/Q sky130_fd_sc_hd__dfxtp_1
X_30066_ _30066_/A VGND VGND VPWR VPWR _35285_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19877_ _19656_/X _19875_/X _19876_/X _19659_/X VGND VGND VPWR VPWR _19877_/X sky130_fd_sc_hd__a22o_1
XFILLER_60_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18828_ _18822_/X _18827_/X _18759_/X VGND VGND VPWR VPWR _18829_/D sky130_fd_sc_hd__o21ba_1
X_34874_ _35448_/CLK _34874_/D VGND VGND VPWR VPWR _34874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33825_ _36065_/CLK _33825_/D VGND VGND VPWR VPWR _33825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18759_ _20171_/A VGND VGND VPWR VPWR _18759_/X sky130_fd_sc_hd__buf_2
XFILLER_243_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21770_ _34165_/Q _34101_/Q _34037_/Q _33973_/Q _21693_/X _21694_/X VGND VGND VPWR
+ VPWR _21770_/X sky130_fd_sc_hd__mux4_1
X_33756_ _33818_/CLK _33756_/D VGND VGND VPWR VPWR _33756_/Q sky130_fd_sc_hd__dfxtp_1
X_30968_ _30968_/A VGND VGND VPWR VPWR _35712_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20721_ _32855_/Q _32791_/Q _32727_/Q _32663_/Q _20637_/X _20639_/X VGND VGND VPWR
+ VPWR _20721_/X sky130_fd_sc_hd__mux4_1
XFILLER_184_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32707_ _32894_/CLK _32707_/D VGND VGND VPWR VPWR _32707_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33687_ _35801_/CLK _33687_/D VGND VGND VPWR VPWR _33687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30899_ _31010_/S VGND VGND VPWR VPWR _30918_/S sky130_fd_sc_hd__buf_4
XFILLER_223_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23440_ _23440_/A VGND VGND VPWR VPWR _32225_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20652_ _22582_/A VGND VGND VPWR VPWR _22598_/A sky130_fd_sc_hd__buf_12
X_35426_ _35553_/CLK _35426_/D VGND VGND VPWR VPWR _35426_/Q sky130_fd_sc_hd__dfxtp_1
X_32638_ _35839_/CLK _32638_/D VGND VGND VPWR VPWR _32638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23371_ _32201_/Q _23302_/X _23385_/S VGND VGND VPWR VPWR _23372_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20583_ _20661_/A VGND VGND VPWR VPWR _22506_/A sky130_fd_sc_hd__buf_12
X_35357_ _35677_/CLK _35357_/D VGND VGND VPWR VPWR _35357_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_393_CLK clkbuf_6_40__f_CLK/X VGND VGND VPWR VPWR _35703_/CLK sky130_fd_sc_hd__clkbuf_16
X_32569_ _36027_/CLK _32569_/D VGND VGND VPWR VPWR _32569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_722 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25110_ _24964_/X _33035_/Q _25122_/S VGND VGND VPWR VPWR _25111_/A sky130_fd_sc_hd__mux2_1
X_22322_ _22111_/X _22320_/X _22321_/X _22116_/X VGND VGND VPWR VPWR _22322_/X sky130_fd_sc_hd__a22o_1
X_34308_ _36164_/CLK _34308_/D VGND VGND VPWR VPWR _34308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26090_ _24809_/X _33497_/Q _26102_/S VGND VGND VPWR VPWR _26091_/A sky130_fd_sc_hd__mux2_1
X_35288_ _35799_/CLK _35288_/D VGND VGND VPWR VPWR _35288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22253_ _22249_/X _22252_/X _22118_/X VGND VGND VPWR VPWR _22254_/D sky130_fd_sc_hd__o21ba_1
X_25041_ _24861_/X _33002_/Q _25059_/S VGND VGND VPWR VPWR _25042_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_145_CLK clkbuf_6_29__f_CLK/X VGND VGND VPWR VPWR _36117_/CLK sky130_fd_sc_hd__clkbuf_16
X_34239_ _36103_/CLK _34239_/D VGND VGND VPWR VPWR _34239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_1402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21204_ _32613_/Q _32549_/Q _32485_/Q _35941_/Q _21170_/X _20954_/X VGND VGND VPWR
+ VPWR _21204_/X sky130_fd_sc_hd__mux4_1
XFILLER_219_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22184_ _34432_/Q _36160_/Q _34304_/Q _34240_/Q _22182_/X _22183_/X VGND VGND VPWR
+ VPWR _22184_/X sky130_fd_sc_hd__mux4_1
XFILLER_144_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28800_ _34715_/Q _27050_/X _28808_/S VGND VGND VPWR VPWR _28801_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21135_ _33891_/Q _33827_/Q _33763_/Q _36067_/Q _20918_/X _20919_/X VGND VGND VPWR
+ VPWR _21135_/X sky130_fd_sc_hd__mux4_1
X_29780_ _29780_/A VGND VGND VPWR VPWR _35149_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26992_ _33922_/Q _23435_/X _27002_/S VGND VGND VPWR VPWR _26993_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28731_ _28731_/A VGND VGND VPWR VPWR _34683_/D sky130_fd_sc_hd__clkbuf_1
X_25943_ _24991_/X _33428_/Q _25945_/S VGND VGND VPWR VPWR _25944_/A sky130_fd_sc_hd__mux2_1
X_21066_ _33377_/Q _33313_/Q _33249_/Q _33185_/Q _21021_/X _21022_/X VGND VGND VPWR
+ VPWR _21066_/X sky130_fd_sc_hd__mux4_1
XFILLER_87_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20017_ _20017_/A VGND VGND VPWR VPWR _20017_/X sky130_fd_sc_hd__buf_4
X_28662_ _28662_/A VGND VGND VPWR VPWR _34650_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25874_ _24889_/X _33395_/Q _25874_/S VGND VGND VPWR VPWR _25875_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1029 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27613_ _34185_/Q _27193_/X _27629_/S VGND VGND VPWR VPWR _27614_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24825_ _24824_/X _32926_/Q _24828_/S VGND VGND VPWR VPWR _24826_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28593_ _28593_/A VGND VGND VPWR VPWR _34618_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27544_ _27544_/A VGND VGND VPWR VPWR _34152_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24756_ _24756_/A VGND VGND VPWR VPWR _32898_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21968_ _34938_/Q _34874_/Q _34810_/Q _34746_/Q _21760_/X _21761_/X VGND VGND VPWR
+ VPWR _21968_/X sky130_fd_sc_hd__mux4_1
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23707_ _31418_/A _27840_/A VGND VGND VPWR VPWR _23840_/S sky130_fd_sc_hd__nand2_8
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27475_ _27502_/S VGND VGND VPWR VPWR _27494_/S sky130_fd_sc_hd__buf_4
XFILLER_187_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20919_ _22451_/A VGND VGND VPWR VPWR _20919_/X sky130_fd_sc_hd__clkbuf_8
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24687_ _24687_/A VGND VGND VPWR VPWR _32865_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21899_ _21758_/X _21897_/X _21898_/X _21763_/X VGND VGND VPWR VPWR _21899_/X sky130_fd_sc_hd__a22o_1
X_29214_ _29214_/A VGND VGND VPWR VPWR _34911_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26426_ _33656_/Q _23402_/X _26436_/S VGND VGND VPWR VPWR _26427_/A sky130_fd_sc_hd__mux2_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23638_ _22987_/X _32310_/Q _23652_/S VGND VGND VPWR VPWR _23639_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29145_ _29145_/A VGND VGND VPWR VPWR _34878_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26357_ _33623_/Q _23234_/X _26373_/S VGND VGND VPWR VPWR _26358_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23569_ _31823_/A _31418_/A VGND VGND VPWR VPWR _23702_/S sky130_fd_sc_hd__nand2_8
XFILLER_11_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_384_CLK clkbuf_6_42__f_CLK/X VGND VGND VPWR VPWR _33914_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_168_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16110_ _15981_/X _16108_/X _16109_/X _15991_/X VGND VGND VPWR VPWR _16110_/X sky130_fd_sc_hd__a22o_1
XFILLER_167_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25308_ _25308_/A VGND VGND VPWR VPWR _33127_/D sky130_fd_sc_hd__clkbuf_1
X_29076_ _34846_/Q _27059_/X _29078_/S VGND VGND VPWR VPWR _29077_/A sky130_fd_sc_hd__mux2_1
X_17090_ _17090_/A _17090_/B _17090_/C _17090_/D VGND VGND VPWR VPWR _17091_/A sky130_fd_sc_hd__or4_4
X_26288_ _24902_/X _33591_/Q _26300_/S VGND VGND VPWR VPWR _26289_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_1226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16041_ _17915_/A VGND VGND VPWR VPWR _16041_/X sky130_fd_sc_hd__buf_4
X_28027_ _34350_/Q _27109_/X _28037_/S VGND VGND VPWR VPWR _28028_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_136_CLK clkbuf_6_23__f_CLK/X VGND VGND VPWR VPWR _35799_/CLK sky130_fd_sc_hd__clkbuf_16
X_25239_ _25239_/A VGND VGND VPWR VPWR _33095_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_237_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19800_ _19651_/X _19796_/X _19799_/X _19654_/X VGND VGND VPWR VPWR _19800_/X sky130_fd_sc_hd__a22o_1
XFILLER_123_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17992_ _35660_/Q _35020_/Q _34380_/Q _33740_/Q _17850_/X _17851_/X VGND VGND VPWR
+ VPWR _17992_/X sky130_fd_sc_hd__mux4_1
XFILLER_2_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29978_ _35243_/Q _29395_/X _29994_/S VGND VGND VPWR VPWR _29979_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19731_ _20235_/A VGND VGND VPWR VPWR _19731_/X sky130_fd_sc_hd__buf_6
X_16943_ _16800_/X _16941_/X _16942_/X _16803_/X VGND VGND VPWR VPWR _16943_/X sky130_fd_sc_hd__a22o_1
XFILLER_81_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28929_ _34776_/Q _27041_/X _28943_/S VGND VGND VPWR VPWR _28930_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31940_ _23472_/X _36173_/Q _31948_/S VGND VGND VPWR VPWR _31941_/A sky130_fd_sc_hd__mux2_1
X_16874_ _35180_/Q _35116_/Q _35052_/Q _32172_/Q _16657_/X _16658_/X VGND VGND VPWR
+ VPWR _16874_/X sky130_fd_sc_hd__mux4_1
X_19662_ _34682_/Q _34618_/Q _34554_/Q _34490_/Q _19592_/X _19593_/X VGND VGND VPWR
+ VPWR _19662_/X sky130_fd_sc_hd__mux4_1
XFILLER_226_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18613_ _18613_/A VGND VGND VPWR VPWR _32412_/D sky130_fd_sc_hd__clkbuf_4
XTAP_4060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31871_ _23299_/X _36140_/Q _31885_/S VGND VGND VPWR VPWR _31872_/A sky130_fd_sc_hd__mux2_1
X_19593_ _20299_/A VGND VGND VPWR VPWR _19593_/X sky130_fd_sc_hd__buf_6
XTAP_4071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_1330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33610_ _33869_/CLK _33610_/D VGND VGND VPWR VPWR _33610_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30822_ _30822_/A VGND VGND VPWR VPWR _35643_/D sky130_fd_sc_hd__clkbuf_1
X_18544_ _33627_/Q _33563_/Q _33499_/Q _33435_/Q _18441_/X _18442_/X VGND VGND VPWR
+ VPWR _18544_/X sky130_fd_sc_hd__mux4_1
XFILLER_18_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34590_ _36229_/CLK _34590_/D VGND VGND VPWR VPWR _34590_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_691 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33541_ _34179_/CLK _33541_/D VGND VGND VPWR VPWR _33541_/Q sky130_fd_sc_hd__dfxtp_1
X_18475_ _18469_/X _18474_/X _18404_/X VGND VGND VPWR VPWR _18476_/D sky130_fd_sc_hd__o21ba_1
X_30753_ _30753_/A VGND VGND VPWR VPWR _35610_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1074 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17426_ _17419_/X _17425_/X _17140_/X _17141_/X VGND VGND VPWR VPWR _17443_/B sky130_fd_sc_hd__o211a_1
XFILLER_221_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33472_ _33984_/CLK _33472_/D VGND VGND VPWR VPWR _33472_/Q sky130_fd_sc_hd__dfxtp_1
X_30684_ _35578_/Q _29441_/X _30690_/S VGND VGND VPWR VPWR _30685_/A sky130_fd_sc_hd__mux2_1
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35211_ _35212_/CLK _35211_/D VGND VGND VPWR VPWR _35211_/Q sky130_fd_sc_hd__dfxtp_1
X_32423_ _36072_/CLK _32423_/D VGND VGND VPWR VPWR _32423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17357_ _35450_/Q _35386_/Q _35322_/Q _35258_/Q _17254_/X _17255_/X VGND VGND VPWR
+ VPWR _17357_/X sky130_fd_sc_hd__mux4_1
X_36191_ _36191_/CLK _36191_/D VGND VGND VPWR VPWR _36191_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_375_CLK clkbuf_6_43__f_CLK/X VGND VGND VPWR VPWR _34877_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_105_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16308_ _34396_/Q _36124_/Q _34268_/Q _34204_/Q _16170_/X _16171_/X VGND VGND VPWR
+ VPWR _16308_/X sky130_fd_sc_hd__mux4_1
XFILLER_201_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35142_ _35718_/CLK _35142_/D VGND VGND VPWR VPWR _35142_/Q sky130_fd_sc_hd__dfxtp_1
X_32354_ _32356_/CLK _32354_/D VGND VGND VPWR VPWR _32354_/Q sky130_fd_sc_hd__dfxtp_1
X_17288_ _35448_/Q _35384_/Q _35320_/Q _35256_/Q _17254_/X _17255_/X VGND VGND VPWR
+ VPWR _17288_/X sky130_fd_sc_hd__mux4_1
XFILLER_118_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19027_ _33064_/Q _32040_/Q _35816_/Q _35752_/Q _19025_/X _19026_/X VGND VGND VPWR
+ VPWR _19027_/X sky130_fd_sc_hd__mux4_1
X_31305_ _31416_/S VGND VGND VPWR VPWR _31324_/S sky130_fd_sc_hd__clkbuf_4
X_16239_ _34906_/Q _34842_/Q _34778_/Q _34714_/Q _16096_/X _16098_/X VGND VGND VPWR
+ VPWR _16239_/X sky130_fd_sc_hd__mux4_1
XFILLER_238_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35073_ _35655_/CLK _35073_/D VGND VGND VPWR VPWR _35073_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_127_CLK clkbuf_6_21__f_CLK/X VGND VGND VPWR VPWR _34907_/CLK sky130_fd_sc_hd__clkbuf_16
X_32285_ _32797_/CLK _32285_/D VGND VGND VPWR VPWR _32285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34024_ _34146_/CLK _34024_/D VGND VGND VPWR VPWR _34024_/Q sky130_fd_sc_hd__dfxtp_1
X_31236_ _27770_/X _35839_/Q _31252_/S VGND VGND VPWR VPWR _31237_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31167_ _31167_/A VGND VGND VPWR VPWR _35806_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_1176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30118_ _30118_/A VGND VGND VPWR VPWR _35309_/D sky130_fd_sc_hd__clkbuf_1
X_19929_ _20282_/A VGND VGND VPWR VPWR _19929_/X sky130_fd_sc_hd__buf_6
XFILLER_214_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35975_ _35975_/CLK _35975_/D VGND VGND VPWR VPWR _35975_/Q sky130_fd_sc_hd__dfxtp_1
X_31098_ _35774_/Q input35/X _31116_/S VGND VGND VPWR VPWR _31099_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_214_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30049_ _35277_/Q _29500_/X _30057_/S VGND VGND VPWR VPWR _30050_/A sky130_fd_sc_hd__mux2_1
X_34926_ _34926_/CLK _34926_/D VGND VGND VPWR VPWR _34926_/Q sky130_fd_sc_hd__dfxtp_1
X_22940_ input9/X VGND VGND VPWR VPWR _22940_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_116_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22871_ _35221_/Q _35157_/Q _35093_/Q _32277_/Q _20692_/X _20694_/X VGND VGND VPWR
+ VPWR _22871_/X sky130_fd_sc_hd__mux4_1
X_34857_ _34921_/CLK _34857_/D VGND VGND VPWR VPWR _34857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24610_ _24610_/A VGND VGND VPWR VPWR _32829_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33808_ _36113_/CLK _33808_/D VGND VGND VPWR VPWR _33808_/Q sky130_fd_sc_hd__dfxtp_1
X_21822_ _35446_/Q _35382_/Q _35318_/Q _35254_/Q _21501_/X _21502_/X VGND VGND VPWR
+ VPWR _21822_/X sky130_fd_sc_hd__mux4_1
X_25590_ _24868_/X _33260_/Q _25604_/S VGND VGND VPWR VPWR _25591_/A sky130_fd_sc_hd__mux2_1
X_34788_ _34790_/CLK _34788_/D VGND VGND VPWR VPWR _34788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24541_ _24541_/A VGND VGND VPWR VPWR _32796_/D sky130_fd_sc_hd__clkbuf_1
X_33739_ _35724_/CLK _33739_/D VGND VGND VPWR VPWR _33739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21753_ _21753_/A VGND VGND VPWR VPWR _21753_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_54_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20704_ _22471_/A VGND VGND VPWR VPWR _20704_/X sky130_fd_sc_hd__clkbuf_4
X_27260_ _27260_/A VGND VGND VPWR VPWR _34017_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24472_ _23005_/X _32764_/Q _24474_/S VGND VGND VPWR VPWR _24473_/A sky130_fd_sc_hd__mux2_1
X_21684_ _35186_/Q _35122_/Q _35058_/Q _32209_/Q _21610_/X _21611_/X VGND VGND VPWR
+ VPWR _21684_/X sky130_fd_sc_hd__mux4_1
X_26211_ _24988_/X _33555_/Q _26215_/S VGND VGND VPWR VPWR _26212_/A sky130_fd_sc_hd__mux2_1
X_35409_ _35859_/CLK _35409_/D VGND VGND VPWR VPWR _35409_/Q sky130_fd_sc_hd__dfxtp_1
X_23423_ _23423_/A VGND VGND VPWR VPWR _32219_/D sky130_fd_sc_hd__clkbuf_1
X_27191_ _33992_/Q _27189_/X _27218_/S VGND VGND VPWR VPWR _27192_/A sky130_fd_sc_hd__mux2_1
X_20635_ _32086_/Q _32278_/Q _32342_/Q _35862_/Q _20632_/X _22467_/A VGND VGND VPWR
+ VPWR _20635_/X sky130_fd_sc_hd__mux4_1
XFILLER_138_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_366_CLK clkbuf_6_41__f_CLK/X VGND VGND VPWR VPWR _35192_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_32_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26142_ _24886_/X _33522_/Q _26144_/S VGND VGND VPWR VPWR _26143_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20566_ _35477_/Q _35413_/Q _35349_/Q _35285_/Q _18309_/X _18311_/X VGND VGND VPWR
+ VPWR _20566_/X sky130_fd_sc_hd__mux4_1
X_23354_ _23354_/A VGND VGND VPWR VPWR _32193_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22305_ _35716_/Q _32226_/Q _35588_/Q _35524_/Q _22270_/X _22271_/X VGND VGND VPWR
+ VPWR _22305_/X sky130_fd_sc_hd__mux4_1
X_26073_ _26073_/A VGND VGND VPWR VPWR _33489_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_118_CLK clkbuf_6_20__f_CLK/X VGND VGND VPWR VPWR _36229_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_164_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20497_ _33171_/Q _36051_/Q _33043_/Q _32979_/Q _18332_/X _19461_/A VGND VGND VPWR
+ VPWR _20497_/X sky130_fd_sc_hd__mux4_1
X_23285_ _23285_/A VGND VGND VPWR VPWR _32167_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29901_ _35207_/Q _29481_/X _29901_/S VGND VGND VPWR VPWR _29902_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25024_ _24837_/X _32994_/Q _25038_/S VGND VGND VPWR VPWR _25025_/A sky130_fd_sc_hd__mux2_1
X_22236_ _22020_/X _22234_/X _22235_/X _22024_/X VGND VGND VPWR VPWR _22236_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22167_ _22012_/X _22165_/X _22166_/X _22018_/X VGND VGND VPWR VPWR _22167_/X sky130_fd_sc_hd__a22o_1
X_29832_ _35174_/Q _29379_/X _29838_/S VGND VGND VPWR VPWR _29833_/A sky130_fd_sc_hd__mux2_1
XTAP_6924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21118_ _20897_/X _21116_/X _21117_/X _20900_/X VGND VGND VPWR VPWR _21118_/X sky130_fd_sc_hd__a22o_1
XTAP_6957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29763_ _29763_/A VGND VGND VPWR VPWR _35141_/D sky130_fd_sc_hd__clkbuf_1
X_22098_ _22451_/A VGND VGND VPWR VPWR _22098_/X sky130_fd_sc_hd__buf_4
XFILLER_8_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26975_ _33914_/Q _23408_/X _26981_/S VGND VGND VPWR VPWR _26976_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25926_ _25926_/A VGND VGND VPWR VPWR _33419_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_247_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28714_ _28714_/A VGND VGND VPWR VPWR _34675_/D sky130_fd_sc_hd__clkbuf_1
X_21049_ _35168_/Q _35104_/Q _35040_/Q _32160_/Q _20904_/X _20905_/X VGND VGND VPWR
+ VPWR _21049_/X sky130_fd_sc_hd__mux4_1
X_29694_ _29694_/A VGND VGND VPWR VPWR _35108_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28645_ _28645_/A VGND VGND VPWR VPWR _34643_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25857_ _25857_/A VGND VGND VPWR VPWR _33386_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24808_ _24808_/A VGND VGND VPWR VPWR _32920_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28576_ _28576_/A VGND VGND VPWR VPWR _34610_/D sky130_fd_sc_hd__clkbuf_1
X_16590_ _16447_/X _16588_/X _16589_/X _16450_/X VGND VGND VPWR VPWR _16590_/X sky130_fd_sc_hd__a22o_1
X_25788_ _24961_/X _33354_/Q _25802_/S VGND VGND VPWR VPWR _25789_/A sky130_fd_sc_hd__mux2_1
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27527_ _34144_/Q _27065_/X _27545_/S VGND VGND VPWR VPWR _27528_/A sky130_fd_sc_hd__mux2_1
XFILLER_243_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24739_ _24739_/A VGND VGND VPWR VPWR _32890_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18260_ _32917_/Q _32853_/Q _32789_/Q _32725_/Q _15984_/X _15987_/X VGND VGND VPWR
+ VPWR _18260_/X sky130_fd_sc_hd__mux4_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27458_ _27458_/A VGND VGND VPWR VPWR _34111_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17211_ _17205_/X _17210_/X _17132_/X VGND VGND VPWR VPWR _17235_/A sky130_fd_sc_hd__o21ba_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26409_ _33648_/Q _23340_/X _26415_/S VGND VGND VPWR VPWR _26410_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18191_ _17905_/X _18189_/X _18190_/X _17910_/X VGND VGND VPWR VPWR _18191_/X sky130_fd_sc_hd__a22o_1
X_27389_ _34079_/Q _27062_/X _27389_/S VGND VGND VPWR VPWR _27390_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_357_CLK clkbuf_6_46__f_CLK/X VGND VGND VPWR VPWR _35644_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_204_1244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29128_ _29128_/A VGND VGND VPWR VPWR _34870_/D sky130_fd_sc_hd__clkbuf_1
X_17142_ _17136_/X _17139_/X _17140_/X _17141_/X VGND VGND VPWR VPWR _17167_/B sky130_fd_sc_hd__o211a_1
XFILLER_204_1277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29059_ _29191_/S VGND VGND VPWR VPWR _29078_/S sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_109_CLK clkbuf_6_22__f_CLK/X VGND VGND VPWR VPWR _34135_/CLK sky130_fd_sc_hd__clkbuf_16
X_17073_ _17066_/X _17072_/X _16787_/X _16788_/X VGND VGND VPWR VPWR _17090_/B sky130_fd_sc_hd__o211a_1
XFILLER_171_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16024_ _17906_/A VGND VGND VPWR VPWR _16024_/X sky130_fd_sc_hd__clkbuf_8
X_32070_ _35974_/CLK _32070_/D VGND VGND VPWR VPWR _32070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31021_ _31021_/A VGND VGND VPWR VPWR _35737_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_836 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17975_ _33676_/Q _33612_/Q _33548_/Q _33484_/Q _17906_/X _17907_/X VGND VGND VPWR
+ VPWR _17975_/X sky130_fd_sc_hd__mux4_1
XFILLER_215_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19714_ _32636_/Q _32572_/Q _32508_/Q _35964_/Q _19576_/X _19713_/X VGND VGND VPWR
+ VPWR _19714_/X sky130_fd_sc_hd__mux4_1
X_35760_ _36147_/CLK _35760_/D VGND VGND VPWR VPWR _35760_/Q sky130_fd_sc_hd__dfxtp_1
X_16926_ _16706_/X _16924_/X _16925_/X _16712_/X VGND VGND VPWR VPWR _16926_/X sky130_fd_sc_hd__a22o_1
X_32972_ _36044_/CLK _32972_/D VGND VGND VPWR VPWR _32972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34711_ _34904_/CLK _34711_/D VGND VGND VPWR VPWR _34711_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31923_ _23444_/X _36165_/Q _31927_/S VGND VGND VPWR VPWR _31924_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19645_ _32122_/Q _32314_/Q _32378_/Q _35898_/Q _19580_/X _19368_/X VGND VGND VPWR
+ VPWR _19645_/X sky130_fd_sc_hd__mux4_1
XFILLER_226_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16857_ _16853_/X _16854_/X _16855_/X _16856_/X VGND VGND VPWR VPWR _16857_/X sky130_fd_sc_hd__a22o_1
X_35691_ _35691_/CLK _35691_/D VGND VGND VPWR VPWR _35691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34642_ _34708_/CLK _34642_/D VGND VGND VPWR VPWR _34642_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19576_ _20282_/A VGND VGND VPWR VPWR _19576_/X sky130_fd_sc_hd__buf_6
X_31854_ _23274_/X _36132_/Q _31864_/S VGND VGND VPWR VPWR _31855_/A sky130_fd_sc_hd__mux2_1
X_16788_ _17847_/A VGND VGND VPWR VPWR _16788_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_209_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_1169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18527_ _35610_/Q _34970_/Q _34330_/Q _33690_/Q _18353_/X _18355_/X VGND VGND VPWR
+ VPWR _18527_/X sky130_fd_sc_hd__mux4_1
X_30805_ _30805_/A VGND VGND VPWR VPWR _35635_/D sky130_fd_sc_hd__clkbuf_1
X_34573_ _35213_/CLK _34573_/D VGND VGND VPWR VPWR _34573_/Q sky130_fd_sc_hd__dfxtp_1
X_31785_ _31785_/A VGND VGND VPWR VPWR _36099_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33524_ _34099_/CLK _33524_/D VGND VGND VPWR VPWR _33524_/Q sky130_fd_sc_hd__dfxtp_1
X_18458_ _18330_/X _18456_/X _18457_/X _18341_/X VGND VGND VPWR VPWR _18458_/X sky130_fd_sc_hd__a22o_1
XFILLER_209_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30736_ _35603_/Q _29518_/X _30740_/S VGND VGND VPWR VPWR _30737_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_1030 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36243_ _36245_/CLK _36243_/D VGND VGND VPWR VPWR _36243_/Q sky130_fd_sc_hd__dfxtp_1
X_17409_ _33916_/Q _33852_/Q _33788_/Q _36092_/Q _17377_/X _17378_/X VGND VGND VPWR
+ VPWR _17409_/X sky130_fd_sc_hd__mux4_1
X_18389_ _18378_/X _18381_/X _18386_/X _18388_/X VGND VGND VPWR VPWR _18389_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_348_CLK clkbuf_6_47__f_CLK/X VGND VGND VPWR VPWR _35454_/CLK sky130_fd_sc_hd__clkbuf_16
X_33455_ _34991_/CLK _33455_/D VGND VGND VPWR VPWR _33455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30667_ _35570_/Q _29416_/X _30669_/S VGND VGND VPWR VPWR _30668_/A sky130_fd_sc_hd__mux2_1
X_20420_ _34704_/Q _34640_/Q _34576_/Q _34512_/Q _20298_/X _20299_/X VGND VGND VPWR
+ VPWR _20420_/X sky130_fd_sc_hd__mux4_1
XFILLER_140_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32406_ _34148_/CLK _32406_/D VGND VGND VPWR VPWR _32406_/Q sky130_fd_sc_hd__dfxtp_1
X_36174_ _36175_/CLK _36174_/D VGND VGND VPWR VPWR _36174_/Q sky130_fd_sc_hd__dfxtp_1
X_30598_ _30598_/A VGND VGND VPWR VPWR _35537_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33386_ _36076_/CLK _33386_/D VGND VGND VPWR VPWR _33386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20351_ _20073_/X _20349_/X _20350_/X _20077_/X VGND VGND VPWR VPWR _20351_/X sky130_fd_sc_hd__a22o_1
X_35125_ _35829_/CLK _35125_/D VGND VGND VPWR VPWR _35125_/Q sky130_fd_sc_hd__dfxtp_1
X_32337_ _32911_/CLK _32337_/D VGND VGND VPWR VPWR _32337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23070_ input55/X VGND VGND VPWR VPWR _23070_/X sky130_fd_sc_hd__buf_2
X_32268_ _35147_/CLK _32268_/D VGND VGND VPWR VPWR _32268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20282_ _20282_/A VGND VGND VPWR VPWR _20282_/X sky130_fd_sc_hd__buf_6
X_35056_ _35056_/CLK _35056_/D VGND VGND VPWR VPWR _35056_/Q sky130_fd_sc_hd__dfxtp_1
X_22021_ _22374_/A VGND VGND VPWR VPWR _22021_/X sky130_fd_sc_hd__clkbuf_4
XTAP_6209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34007_ _34007_/CLK _34007_/D VGND VGND VPWR VPWR _34007_/Q sky130_fd_sc_hd__dfxtp_1
X_31219_ _27745_/X _35831_/Q _31231_/S VGND VGND VPWR VPWR _31220_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32199_ _34987_/CLK _32199_/D VGND VGND VPWR VPWR _32199_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26760_ _26760_/A VGND VGND VPWR VPWR _33812_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23972_ _23972_/A VGND VGND VPWR VPWR _32530_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35958_ _36021_/CLK _35958_/D VGND VGND VPWR VPWR _35958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25711_ _25711_/A VGND VGND VPWR VPWR _33317_/D sky130_fd_sc_hd__clkbuf_1
X_34909_ _34911_/CLK _34909_/D VGND VGND VPWR VPWR _34909_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_1135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22923_ _22922_/X _32033_/Q _22947_/S VGND VGND VPWR VPWR _22924_/A sky130_fd_sc_hd__mux2_1
X_26691_ _26691_/A VGND VGND VPWR VPWR _33779_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35889_ _35952_/CLK _35889_/D VGND VGND VPWR VPWR _35889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28430_ _27714_/X _34541_/Q _28442_/S VGND VGND VPWR VPWR _28431_/A sky130_fd_sc_hd__mux2_1
X_25642_ _24945_/X _33285_/Q _25646_/S VGND VGND VPWR VPWR _25643_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22854_ _20630_/X _22852_/X _22853_/X _20641_/X VGND VGND VPWR VPWR _22854_/X sky130_fd_sc_hd__a22o_1
XFILLER_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28361_ _28361_/A VGND VGND VPWR VPWR _34508_/D sky130_fd_sc_hd__clkbuf_1
X_21805_ _21799_/X _21802_/X _21803_/X _21804_/X VGND VGND VPWR VPWR _21805_/X sky130_fd_sc_hd__a22o_1
XFILLER_45_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25573_ _24843_/X _33252_/Q _25583_/S VGND VGND VPWR VPWR _25574_/A sky130_fd_sc_hd__mux2_1
X_22785_ _20660_/X _22783_/X _22784_/X _20672_/X VGND VGND VPWR VPWR _22785_/X sky130_fd_sc_hd__a22o_1
XFILLER_169_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27312_ _27312_/A VGND VGND VPWR VPWR _34042_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_213_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24524_ _23082_/X _32789_/Q _24524_/S VGND VGND VPWR VPWR _24525_/A sky130_fd_sc_hd__mux2_1
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28292_ _28292_/A VGND VGND VPWR VPWR _34475_/D sky130_fd_sc_hd__clkbuf_1
X_21736_ _21659_/X _21734_/X _21735_/X _21665_/X VGND VGND VPWR VPWR _21736_/X sky130_fd_sc_hd__a22o_1
XFILLER_212_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27243_ _27243_/A VGND VGND VPWR VPWR _34009_/D sky130_fd_sc_hd__clkbuf_1
X_24455_ _24524_/S VGND VGND VPWR VPWR _24474_/S sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_339_CLK clkbuf_6_45__f_CLK/X VGND VGND VPWR VPWR _32889_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_185_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21667_ _22512_/A VGND VGND VPWR VPWR _21667_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_8_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_1114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23406_ _32214_/Q _23405_/X _23418_/S VGND VGND VPWR VPWR _23407_/A sky130_fd_sc_hd__mux2_1
X_20618_ _22505_/A VGND VGND VPWR VPWR _20618_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_177_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27174_ input40/X VGND VGND VPWR VPWR _27174_/X sky130_fd_sc_hd__buf_4
XFILLER_32_1136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24386_ _24386_/A VGND VGND VPWR VPWR _32723_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21598_ _22459_/A VGND VGND VPWR VPWR _21598_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_6_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26125_ _26215_/S VGND VGND VPWR VPWR _26144_/S sky130_fd_sc_hd__buf_4
X_23337_ _23499_/S VGND VGND VPWR VPWR _23359_/S sky130_fd_sc_hd__buf_4
X_20549_ _33685_/Q _33621_/Q _33557_/Q _33493_/Q _18324_/X _18325_/X VGND VGND VPWR
+ VPWR _20549_/X sky130_fd_sc_hd__mux4_1
XFILLER_126_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26056_ _24958_/X _33481_/Q _26072_/S VGND VGND VPWR VPWR _26057_/A sky130_fd_sc_hd__mux2_1
X_23268_ input4/X VGND VGND VPWR VPWR _23268_/X sky130_fd_sc_hd__buf_4
X_25007_ _24812_/X _32986_/Q _25017_/S VGND VGND VPWR VPWR _25008_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22219_ _22215_/X _22218_/X _22118_/X VGND VGND VPWR VPWR _22220_/D sky130_fd_sc_hd__o21ba_1
XFILLER_193_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23199_ _23046_/X _32137_/Q _23215_/S VGND VGND VPWR VPWR _23200_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29815_ _35166_/Q _29354_/X _29817_/S VGND VGND VPWR VPWR _29816_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17760_ _17552_/X _17758_/X _17759_/X _17557_/X VGND VGND VPWR VPWR _17760_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29746_ _29746_/A VGND VGND VPWR VPWR _35133_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26958_ _33906_/Q _23381_/X _26960_/S VGND VGND VPWR VPWR _26959_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16711_ _33128_/Q _36008_/Q _33000_/Q _32936_/Q _16709_/X _16710_/X VGND VGND VPWR
+ VPWR _16711_/X sky130_fd_sc_hd__mux4_1
X_17691_ _33412_/Q _33348_/Q _33284_/Q _33220_/Q _17480_/X _17481_/X VGND VGND VPWR
+ VPWR _17691_/X sky130_fd_sc_hd__mux4_1
X_25909_ _25909_/A VGND VGND VPWR VPWR _33411_/D sky130_fd_sc_hd__clkbuf_1
X_26889_ _26889_/A VGND VGND VPWR VPWR _33873_/D sky130_fd_sc_hd__clkbuf_1
X_29677_ _29677_/A VGND VGND VPWR VPWR _35100_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19430_ _33908_/Q _33844_/Q _33780_/Q _36084_/Q _19324_/X _19325_/X VGND VGND VPWR
+ VPWR _19430_/X sky130_fd_sc_hd__mux4_1
XFILLER_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16642_ _32870_/Q _32806_/Q _32742_/Q _32678_/Q _16640_/X _16641_/X VGND VGND VPWR
+ VPWR _16642_/X sky130_fd_sc_hd__mux4_1
X_28628_ _27807_/X _34635_/Q _28640_/S VGND VGND VPWR VPWR _28629_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_831 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19361_ _32626_/Q _32562_/Q _32498_/Q _35954_/Q _19223_/X _19360_/X VGND VGND VPWR
+ VPWR _19361_/X sky130_fd_sc_hd__mux4_1
X_16573_ _16353_/X _16571_/X _16572_/X _16359_/X VGND VGND VPWR VPWR _16573_/X sky130_fd_sc_hd__a22o_1
X_28559_ _27704_/X _34602_/Q _28577_/S VGND VGND VPWR VPWR _28560_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18312_ _33878_/Q _33814_/Q _33750_/Q _36054_/Q _18309_/X _18311_/X VGND VGND VPWR
+ VPWR _18312_/X sky130_fd_sc_hd__mux4_1
X_31570_ _31570_/A VGND VGND VPWR VPWR _35997_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19292_ _32112_/Q _32304_/Q _32368_/Q _35888_/Q _19227_/X _19015_/X VGND VGND VPWR
+ VPWR _19292_/X sky130_fd_sc_hd__mux4_1
XFILLER_204_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18243_ _34452_/Q _36180_/Q _34324_/Q _34260_/Q _16067_/X _16069_/X VGND VGND VPWR
+ VPWR _18243_/X sky130_fd_sc_hd__mux4_1
XFILLER_187_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30521_ _30521_/A VGND VGND VPWR VPWR _35500_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_203_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18174_ _35666_/Q _35026_/Q _34386_/Q _33746_/Q _16112_/X _16113_/X VGND VGND VPWR
+ VPWR _18174_/X sky130_fd_sc_hd__mux4_1
X_30452_ _35468_/Q _29497_/X _30462_/S VGND VGND VPWR VPWR _30453_/A sky130_fd_sc_hd__mux2_1
X_33240_ _36057_/CLK _33240_/D VGND VGND VPWR VPWR _33240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17125_ _34164_/Q _34100_/Q _34036_/Q _33972_/Q _17093_/X _17094_/X VGND VGND VPWR
+ VPWR _17125_/X sky130_fd_sc_hd__mux4_1
X_33171_ _35857_/CLK _33171_/D VGND VGND VPWR VPWR _33171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30383_ _35435_/Q _29395_/X _30399_/S VGND VGND VPWR VPWR _30384_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32122_ _35962_/CLK _32122_/D VGND VGND VPWR VPWR _32122_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_1438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17056_ _33906_/Q _33842_/Q _33778_/Q _36082_/Q _17024_/X _17025_/X VGND VGND VPWR
+ VPWR _17056_/X sky130_fd_sc_hd__mux4_1
X_16007_ _17915_/A VGND VGND VPWR VPWR _16007_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_48_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32053_ _35126_/CLK _32053_/D VGND VGND VPWR VPWR _32053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_502_CLK clkbuf_6_2__f_CLK/X VGND VGND VPWR VPWR _33828_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_112_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31004_ _35730_/Q input57/X _31010_/S VGND VGND VPWR VPWR _31005_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1078 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35812_ _35812_/CLK _35812_/D VGND VGND VPWR VPWR _35812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17958_ _35659_/Q _35019_/Q _34379_/Q _33739_/Q _17850_/X _17851_/X VGND VGND VPWR
+ VPWR _17958_/X sky130_fd_sc_hd__mux4_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35743_ _35743_/CLK _35743_/D VGND VGND VPWR VPWR _35743_/Q sky130_fd_sc_hd__dfxtp_1
X_16909_ _16800_/X _16907_/X _16908_/X _16803_/X VGND VGND VPWR VPWR _16909_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_1387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32955_ _35191_/CLK _32955_/D VGND VGND VPWR VPWR _32955_/Q sky130_fd_sc_hd__dfxtp_1
X_17889_ _35721_/Q _32232_/Q _35593_/Q _35529_/Q _17670_/X _17671_/X VGND VGND VPWR
+ VPWR _17889_/X sky130_fd_sc_hd__mux4_1
XFILLER_122_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31906_ _23417_/X _36157_/Q _31906_/S VGND VGND VPWR VPWR _31907_/A sky130_fd_sc_hd__mux2_1
X_19628_ _19453_/X _19626_/X _19627_/X _19456_/X VGND VGND VPWR VPWR _19628_/X sky130_fd_sc_hd__a22o_1
XFILLER_214_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35674_ _35674_/CLK _35674_/D VGND VGND VPWR VPWR _35674_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32886_ _32901_/CLK _32886_/D VGND VGND VPWR VPWR _32886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34625_ _34690_/CLK _34625_/D VGND VGND VPWR VPWR _34625_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31837_ _23249_/X _36124_/Q _31843_/S VGND VGND VPWR VPWR _31838_/A sky130_fd_sc_hd__mux2_1
XFILLER_179_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19559_ _19553_/X _19558_/X _19451_/X VGND VGND VPWR VPWR _19567_/C sky130_fd_sc_hd__o21ba_1
XFILLER_179_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22570_ _34955_/Q _34891_/Q _34827_/Q _34763_/Q _22466_/X _22467_/X VGND VGND VPWR
+ VPWR _22570_/X sky130_fd_sc_hd__mux4_1
XFILLER_224_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34556_ _35193_/CLK _34556_/D VGND VGND VPWR VPWR _34556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31768_ _31768_/A VGND VGND VPWR VPWR _36091_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_845 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21521_ _21453_/X _21519_/X _21520_/X _21456_/X VGND VGND VPWR VPWR _21521_/X sky130_fd_sc_hd__a22o_1
X_33507_ _34151_/CLK _33507_/D VGND VGND VPWR VPWR _33507_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30719_ _30719_/A VGND VGND VPWR VPWR _35594_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_179_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34487_ _36024_/CLK _34487_/D VGND VGND VPWR VPWR _34487_/Q sky130_fd_sc_hd__dfxtp_1
X_31699_ _31699_/A VGND VGND VPWR VPWR _36058_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36226_ _36229_/CLK _36226_/D VGND VGND VPWR VPWR _36226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24240_ _24240_/A VGND VGND VPWR VPWR _32655_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33438_ _36191_/CLK _33438_/D VGND VGND VPWR VPWR _33438_/Q sky130_fd_sc_hd__dfxtp_1
X_21452_ _21446_/X _21449_/X _21450_/X _21451_/X VGND VGND VPWR VPWR _21452_/X sky130_fd_sc_hd__a22o_1
XFILLER_31_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20403_ _33936_/Q _33872_/Q _33808_/Q _36112_/Q _18362_/X _18364_/X VGND VGND VPWR
+ VPWR _20403_/X sky130_fd_sc_hd__mux4_1
XFILLER_135_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36157_ _36157_/CLK _36157_/D VGND VGND VPWR VPWR _36157_/Q sky130_fd_sc_hd__dfxtp_1
X_21383_ _21306_/X _21381_/X _21382_/X _21312_/X VGND VGND VPWR VPWR _21383_/X sky130_fd_sc_hd__a22o_1
X_24171_ _24171_/A VGND VGND VPWR VPWR _32622_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33369_ _36057_/CLK _33369_/D VGND VGND VPWR VPWR _33369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35108_ _35553_/CLK _35108_/D VGND VGND VPWR VPWR _35108_/Q sky130_fd_sc_hd__dfxtp_1
X_23122_ _23122_/A VGND VGND VPWR VPWR _32100_/D sky130_fd_sc_hd__clkbuf_1
X_20334_ _34957_/Q _34893_/Q _34829_/Q _34765_/Q _20166_/X _20167_/X VGND VGND VPWR
+ VPWR _20334_/X sky130_fd_sc_hd__mux4_1
XFILLER_134_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36088_ _36090_/CLK _36088_/D VGND VGND VPWR VPWR _36088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27930_ _27773_/X _34304_/Q _27944_/S VGND VGND VPWR VPWR _27931_/A sky130_fd_sc_hd__mux2_1
X_35039_ _35610_/CLK _35039_/D VGND VGND VPWR VPWR _35039_/Q sky130_fd_sc_hd__dfxtp_1
X_20265_ _20259_/X _20264_/X _20157_/X VGND VGND VPWR VPWR _20273_/C sky130_fd_sc_hd__o21ba_1
X_23053_ _23052_/X _32075_/Q _23071_/S VGND VGND VPWR VPWR _23054_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22004_ _22004_/A VGND VGND VPWR VPWR _36219_/D sky130_fd_sc_hd__clkbuf_2
X_27861_ _27861_/A VGND VGND VPWR VPWR _34271_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20196_ _34697_/Q _34633_/Q _34569_/Q _34505_/Q _19945_/X _19946_/X VGND VGND VPWR
+ VPWR _20196_/X sky130_fd_sc_hd__mux4_1
XTAP_5305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29600_ _35064_/Q _29435_/X _29610_/S VGND VGND VPWR VPWR _29601_/A sky130_fd_sc_hd__mux2_1
XTAP_4604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26812_ _26812_/A VGND VGND VPWR VPWR _33836_/D sky130_fd_sc_hd__clkbuf_1
X_27792_ _27791_/X _34246_/Q _27795_/S VGND VGND VPWR VPWR _27793_/A sky130_fd_sc_hd__mux2_1
XTAP_5349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29531_ _35031_/Q _29333_/X _29547_/S VGND VGND VPWR VPWR _29532_/A sky130_fd_sc_hd__mux2_1
X_26743_ _33804_/Q _23469_/X _26753_/S VGND VGND VPWR VPWR _26744_/A sky130_fd_sc_hd__mux2_1
XTAP_4648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23955_ _23049_/X _32522_/Q _23969_/S VGND VGND VPWR VPWR _23956_/A sky130_fd_sc_hd__mux2_1
XTAP_3914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_854 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29462_ _29462_/A VGND VGND VPWR VPWR _35008_/D sky130_fd_sc_hd__clkbuf_1
X_22906_ input61/X VGND VGND VPWR VPWR _22906_/X sky130_fd_sc_hd__buf_2
XTAP_3947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26674_ _33771_/Q _23296_/X _26690_/S VGND VGND VPWR VPWR _26675_/A sky130_fd_sc_hd__mux2_1
XFILLER_57_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23886_ _23886_/A VGND VGND VPWR VPWR _32489_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_244_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25625_ _24920_/X _33277_/Q _25625_/S VGND VGND VPWR VPWR _25626_/A sky130_fd_sc_hd__mux2_1
X_28413_ _27689_/X _34533_/Q _28421_/S VGND VGND VPWR VPWR _28414_/A sky130_fd_sc_hd__mux2_1
XFILLER_189_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22837_ _33108_/Q _32084_/Q _35860_/Q _35796_/Q _20679_/X _20680_/X VGND VGND VPWR
+ VPWR _22837_/X sky130_fd_sc_hd__mux4_1
X_29393_ _34986_/Q _29391_/X _29420_/S VGND VGND VPWR VPWR _29394_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28344_ _28344_/A VGND VGND VPWR VPWR _34500_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25556_ _24818_/X _33244_/Q _25562_/S VGND VGND VPWR VPWR _25557_/A sky130_fd_sc_hd__mux2_1
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22768_ _21753_/A _22766_/X _22767_/X _21756_/A VGND VGND VPWR VPWR _22768_/X sky130_fd_sc_hd__a22o_1
XFILLER_25_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24507_ _24507_/A VGND VGND VPWR VPWR _32780_/D sky130_fd_sc_hd__clkbuf_1
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21719_ _34931_/Q _34867_/Q _34803_/Q _34739_/Q _21407_/X _21408_/X VGND VGND VPWR
+ VPWR _21719_/X sky130_fd_sc_hd__mux4_1
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28275_ _28275_/A VGND VGND VPWR VPWR _34467_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_839 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25487_ _25487_/A VGND VGND VPWR VPWR _33211_/D sky130_fd_sc_hd__clkbuf_1
X_22699_ _33680_/Q _33616_/Q _33552_/Q _33488_/Q _22506_/X _22507_/X VGND VGND VPWR
+ VPWR _22699_/X sky130_fd_sc_hd__mux4_1
XFILLER_200_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27226_ input59/X VGND VGND VPWR VPWR _27226_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_169_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24438_ _24438_/A VGND VGND VPWR VPWR _32747_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27157_ _27157_/A VGND VGND VPWR VPWR _33981_/D sky130_fd_sc_hd__clkbuf_1
X_24369_ _23052_/X _32715_/Q _24381_/S VGND VGND VPWR VPWR _24370_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26108_ _26108_/A VGND VGND VPWR VPWR _33505_/D sky130_fd_sc_hd__clkbuf_1
X_27088_ _33959_/Q _27087_/X _27094_/S VGND VGND VPWR VPWR _27089_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26039_ _24933_/X _33473_/Q _26051_/S VGND VGND VPWR VPWR _26040_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18930_ _34150_/Q _34086_/Q _34022_/Q _33958_/Q _18687_/X _18688_/X VGND VGND VPWR
+ VPWR _18930_/X sky130_fd_sc_hd__mux4_1
XFILLER_234_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_40_CLK clkbuf_6_7__f_CLK/X VGND VGND VPWR VPWR _35941_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_134_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18861_ _18861_/A _18861_/B _18861_/C _18861_/D VGND VGND VPWR VPWR _18862_/A sky130_fd_sc_hd__or4_2
XTAP_6540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17812_ _17773_/X _17810_/X _17811_/X _17777_/X VGND VGND VPWR VPWR _17812_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18792_ _18792_/A VGND VGND VPWR VPWR _32417_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17743_ _35653_/Q _35013_/Q _34373_/Q _33733_/Q _17497_/X _17498_/X VGND VGND VPWR
+ VPWR _17743_/X sky130_fd_sc_hd__mux4_1
XFILLER_134_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29729_ _35125_/Q _29426_/X _29745_/S VGND VGND VPWR VPWR _29730_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32740_ _32804_/CLK _32740_/D VGND VGND VPWR VPWR _32740_/Q sky130_fd_sc_hd__dfxtp_1
X_17674_ _17351_/X _17672_/X _17673_/X _17354_/X VGND VGND VPWR VPWR _17674_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19413_ _19303_/X _19411_/X _19412_/X _19306_/X VGND VGND VPWR VPWR _19413_/X sky130_fd_sc_hd__a22o_1
XFILLER_78_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16625_ _16452_/X _16623_/X _16624_/X _16457_/X VGND VGND VPWR VPWR _16625_/X sky130_fd_sc_hd__a22o_1
X_32671_ _35870_/CLK _32671_/D VGND VGND VPWR VPWR _32671_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34410_ _34413_/CLK _34410_/D VGND VGND VPWR VPWR _34410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19344_ _35185_/Q _35121_/Q _35057_/Q _32198_/Q _19310_/X _19311_/X VGND VGND VPWR
+ VPWR _19344_/X sky130_fd_sc_hd__mux4_1
X_31622_ _27742_/X _36022_/Q _31636_/S VGND VGND VPWR VPWR _31623_/A sky130_fd_sc_hd__mux2_1
X_16556_ _16447_/X _16554_/X _16555_/X _16450_/X VGND VGND VPWR VPWR _16556_/X sky130_fd_sc_hd__a22o_1
X_35390_ _35454_/CLK _35390_/D VGND VGND VPWR VPWR _35390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34341_ _35620_/CLK _34341_/D VGND VGND VPWR VPWR _34341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31553_ _31553_/A _31553_/B VGND VGND VPWR VPWR _31686_/S sky130_fd_sc_hd__nand2_8
X_16487_ _34401_/Q _36129_/Q _34273_/Q _34209_/Q _16170_/X _16171_/X VGND VGND VPWR
+ VPWR _16487_/X sky130_fd_sc_hd__mux4_2
X_19275_ _19100_/X _19273_/X _19274_/X _19103_/X VGND VGND VPWR VPWR _19275_/X sky130_fd_sc_hd__a22o_1
XFILLER_206_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18226_ _32660_/Q _32596_/Q _32532_/Q _35988_/Q _17982_/X _16877_/A VGND VGND VPWR
+ VPWR _18226_/X sky130_fd_sc_hd__mux4_1
X_30504_ _30504_/A VGND VGND VPWR VPWR _35492_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_176_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34272_ _36128_/CLK _34272_/D VGND VGND VPWR VPWR _34272_/Q sky130_fd_sc_hd__dfxtp_1
X_31484_ _31484_/A VGND VGND VPWR VPWR _35956_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36011_ _36011_/CLK _36011_/D VGND VGND VPWR VPWR _36011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33223_ _36101_/CLK _33223_/D VGND VGND VPWR VPWR _33223_/Q sky130_fd_sc_hd__dfxtp_1
X_30435_ _35460_/Q _29472_/X _30441_/S VGND VGND VPWR VPWR _30436_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18157_ _18157_/A _18157_/B _18157_/C _18157_/D VGND VGND VPWR VPWR _18158_/A sky130_fd_sc_hd__or4_4
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17108_ _35699_/Q _32207_/Q _35571_/Q _35507_/Q _16964_/X _16965_/X VGND VGND VPWR
+ VPWR _17108_/X sky130_fd_sc_hd__mux4_1
X_18088_ _16001_/X _18086_/X _18087_/X _16007_/X VGND VGND VPWR VPWR _18088_/X sky130_fd_sc_hd__a22o_1
X_33154_ _36034_/CLK _33154_/D VGND VGND VPWR VPWR _33154_/Q sky130_fd_sc_hd__dfxtp_1
X_30366_ _35427_/Q _29370_/X _30378_/S VGND VGND VPWR VPWR _30367_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_875 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17039_ _35441_/Q _35377_/Q _35313_/Q _35249_/Q _16901_/X _16902_/X VGND VGND VPWR
+ VPWR _17039_/X sky130_fd_sc_hd__mux4_1
X_32105_ _35947_/CLK _32105_/D VGND VGND VPWR VPWR _32105_/Q sky130_fd_sc_hd__dfxtp_1
X_33085_ _35453_/CLK _33085_/D VGND VGND VPWR VPWR _33085_/Q sky130_fd_sc_hd__dfxtp_1
X_30297_ _30297_/A VGND VGND VPWR VPWR _35394_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_31_CLK clkbuf_6_5__f_CLK/X VGND VGND VPWR VPWR _36128_/CLK sky130_fd_sc_hd__clkbuf_16
X_20050_ _35205_/Q _35141_/Q _35077_/Q _32261_/Q _20016_/X _20017_/X VGND VGND VPWR
+ VPWR _20050_/X sky130_fd_sc_hd__mux4_1
X_32036_ _35814_/CLK _32036_/D VGND VGND VPWR VPWR _32036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33987_ _34183_/CLK _33987_/D VGND VGND VPWR VPWR _33987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35726_ _35727_/CLK _35726_/D VGND VGND VPWR VPWR _35726_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23740_ _22934_/X _32357_/Q _23748_/S VGND VGND VPWR VPWR _23741_/A sky130_fd_sc_hd__mux2_1
XFILLER_227_876 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20952_ _20948_/X _20951_/X _20615_/X VGND VGND VPWR VPWR _20984_/A sky130_fd_sc_hd__o21ba_1
X_32938_ _36141_/CLK _32938_/D VGND VGND VPWR VPWR _32938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_242_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35657_ _35657_/CLK _35657_/D VGND VGND VPWR VPWR _35657_/Q sky130_fd_sc_hd__dfxtp_1
X_23671_ _23036_/X _32326_/Q _23673_/S VGND VGND VPWR VPWR _23672_/A sky130_fd_sc_hd__mux2_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_98_CLK clkbuf_leaf_99_CLK/A VGND VGND VPWR VPWR _33818_/CLK sky130_fd_sc_hd__clkbuf_16
X_20883_ _32604_/Q _32540_/Q _32476_/Q _35932_/Q _20817_/X _22317_/A VGND VGND VPWR
+ VPWR _20883_/X sky130_fd_sc_hd__mux4_1
X_32869_ _32869_/CLK _32869_/D VGND VGND VPWR VPWR _32869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25410_ _25410_/A VGND VGND VPWR VPWR _33174_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22622_ _22618_/X _22621_/X _22446_/X _22447_/X VGND VGND VPWR VPWR _22637_/B sky130_fd_sc_hd__o211a_2
X_34608_ _36143_/CLK _34608_/D VGND VGND VPWR VPWR _34608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26390_ _33639_/Q _23283_/X _26394_/S VGND VGND VPWR VPWR _26391_/A sky130_fd_sc_hd__mux2_1
X_35588_ _35716_/CLK _35588_/D VGND VGND VPWR VPWR _35588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25341_ _33143_/Q _23399_/X _25353_/S VGND VGND VPWR VPWR _25342_/A sky130_fd_sc_hd__mux2_1
X_22553_ _32139_/Q _32331_/Q _32395_/Q _35915_/Q _22233_/X _22374_/X VGND VGND VPWR
+ VPWR _22553_/X sky130_fd_sc_hd__mux4_1
X_34539_ _35754_/CLK _34539_/D VGND VGND VPWR VPWR _34539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28060_ _28108_/S VGND VGND VPWR VPWR _28079_/S sky130_fd_sc_hd__buf_4
X_21504_ _33069_/Q _32045_/Q _35821_/Q _35757_/Q _21325_/X _21326_/X VGND VGND VPWR
+ VPWR _21504_/X sky130_fd_sc_hd__mux4_1
X_25272_ _33110_/Q _23225_/X _25290_/S VGND VGND VPWR VPWR _25273_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22484_ _22365_/X _22482_/X _22483_/X _22371_/X VGND VGND VPWR VPWR _22484_/X sky130_fd_sc_hd__a22o_1
X_27011_ _33931_/Q _23466_/X _27023_/S VGND VGND VPWR VPWR _27012_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24223_ _24223_/A VGND VGND VPWR VPWR _32647_/D sky130_fd_sc_hd__clkbuf_1
X_36209_ _36209_/CLK _36209_/D VGND VGND VPWR VPWR _36209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21435_ _21250_/X _21433_/X _21434_/X _21253_/X VGND VGND VPWR VPWR _21435_/X sky130_fd_sc_hd__a22o_1
XFILLER_213_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24154_ _24154_/A VGND VGND VPWR VPWR _32614_/D sky130_fd_sc_hd__clkbuf_1
X_21366_ _34921_/Q _34857_/Q _34793_/Q _34729_/Q _21054_/X _21055_/X VGND VGND VPWR
+ VPWR _21366_/X sky130_fd_sc_hd__mux4_1
XFILLER_68_1338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23105_ _23105_/A VGND VGND VPWR VPWR _32092_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20317_ _33165_/Q _36045_/Q _33037_/Q _32973_/Q _20068_/X _20069_/X VGND VGND VPWR
+ VPWR _20317_/X sky130_fd_sc_hd__mux4_1
X_24085_ _24085_/A VGND VGND VPWR VPWR _32583_/D sky130_fd_sc_hd__clkbuf_1
X_28962_ _34792_/Q _27090_/X _28964_/S VGND VGND VPWR VPWR _28963_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21297_ _21297_/A _21297_/B _21297_/C _21297_/D VGND VGND VPWR VPWR _21298_/A sky130_fd_sc_hd__or4_4
Xclkbuf_leaf_22_CLK clkbuf_6_4__f_CLK/X VGND VGND VPWR VPWR _34405_/CLK sky130_fd_sc_hd__clkbuf_16
X_23036_ input43/X VGND VGND VPWR VPWR _23036_/X sky130_fd_sc_hd__buf_2
X_27913_ _27748_/X _34296_/Q _27923_/S VGND VGND VPWR VPWR _27914_/A sky130_fd_sc_hd__mux2_1
X_20248_ _20212_/X _20246_/X _20247_/X _20215_/X VGND VGND VPWR VPWR _20248_/X sky130_fd_sc_hd__a22o_1
XFILLER_157_1190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28893_ _28893_/A VGND VGND VPWR VPWR _34759_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27844_ _27646_/X _34263_/Q _27860_/S VGND VGND VPWR VPWR _27845_/A sky130_fd_sc_hd__mux2_1
X_20179_ _33929_/Q _33865_/Q _33801_/Q _36105_/Q _20030_/X _20031_/X VGND VGND VPWR
+ VPWR _20179_/X sky130_fd_sc_hd__mux4_1
XTAP_5135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_859 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27775_ _27775_/A VGND VGND VPWR VPWR _34240_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24987_ _24987_/A VGND VGND VPWR VPWR _32978_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29514_ _29514_/A VGND VGND VPWR VPWR _35025_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26726_ _33796_/Q _23441_/X _26732_/S VGND VGND VPWR VPWR _26727_/A sky130_fd_sc_hd__mux2_1
X_23938_ _23024_/X _32514_/Q _23948_/S VGND VGND VPWR VPWR _23939_/A sky130_fd_sc_hd__mux2_1
XTAP_3744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26657_ _33763_/Q _23271_/X _26669_/S VGND VGND VPWR VPWR _26658_/A sky130_fd_sc_hd__mux2_1
X_29445_ _35003_/Q _29444_/X _29451_/S VGND VGND VPWR VPWR _29446_/A sky130_fd_sc_hd__mux2_1
XFILLER_232_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23869_ _22922_/X _32481_/Q _23885_/S VGND VGND VPWR VPWR _23870_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_89_CLK clkbuf_leaf_96_CLK/A VGND VGND VPWR VPWR _35613_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_205_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16410_ _35167_/Q _35103_/Q _35039_/Q _32159_/Q _16304_/X _16305_/X VGND VGND VPWR
+ VPWR _16410_/X sky130_fd_sc_hd__mux4_1
XFILLER_199_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25608_ _25608_/A VGND VGND VPWR VPWR _33268_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17390_ _35643_/Q _35003_/Q _34363_/Q _33723_/Q _17144_/X _17145_/X VGND VGND VPWR
+ VPWR _17390_/X sky130_fd_sc_hd__mux4_1
XFILLER_77_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26588_ _26588_/A VGND VGND VPWR VPWR _33732_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29376_ input7/X VGND VGND VPWR VPWR _29376_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_246_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16341_ _34909_/Q _34845_/Q _34781_/Q _34717_/Q _16096_/X _16098_/X VGND VGND VPWR
+ VPWR _16341_/X sky130_fd_sc_hd__mux4_1
X_25539_ _25539_/A VGND VGND VPWR VPWR _33236_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_213_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28327_ _28327_/A VGND VGND VPWR VPWR _34492_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19060_ _18950_/X _19058_/X _19059_/X _18953_/X VGND VGND VPWR VPWR _19060_/X sky130_fd_sc_hd__a22o_1
X_16272_ _16091_/X _16270_/X _16271_/X _16101_/X VGND VGND VPWR VPWR _16272_/X sky130_fd_sc_hd__a22o_1
X_28258_ _28258_/A VGND VGND VPWR VPWR _34459_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27209_ _33998_/Q _27208_/X _27218_/S VGND VGND VPWR VPWR _27210_/A sky130_fd_sc_hd__mux2_1
X_18011_ _17905_/X _18009_/X _18010_/X _17910_/X VGND VGND VPWR VPWR _18011_/X sky130_fd_sc_hd__a22o_1
XFILLER_185_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28189_ _27757_/X _34427_/Q _28193_/S VGND VGND VPWR VPWR _28190_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30220_ _35358_/Q _29354_/X _30222_/S VGND VGND VPWR VPWR _30221_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30151_ _30151_/A VGND VGND VPWR VPWR _35325_/D sky130_fd_sc_hd__clkbuf_1
X_19962_ _19958_/X _19961_/X _19785_/X VGND VGND VPWR VPWR _19986_/A sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_13_CLK clkbuf_6_3__f_CLK/X VGND VGND VPWR VPWR _35176_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_45_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18913_ _35685_/Q _32192_/Q _35557_/Q _35493_/Q _18911_/X _18912_/X VGND VGND VPWR
+ VPWR _18913_/X sky130_fd_sc_hd__mux4_2
XTAP_7060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30082_ _30082_/A VGND VGND VPWR VPWR _35292_/D sky130_fd_sc_hd__clkbuf_1
XTAP_7071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19893_ _33409_/Q _33345_/Q _33281_/Q _33217_/Q _19780_/X _19781_/X VGND VGND VPWR
+ VPWR _19893_/X sky130_fd_sc_hd__mux4_1
XFILLER_171_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33910_ _33910_/CLK _33910_/D VGND VGND VPWR VPWR _33910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18844_ _18840_/X _18843_/X _18734_/X _18735_/X VGND VGND VPWR VPWR _18861_/B sky130_fd_sc_hd__o211a_1
X_34890_ _34954_/CLK _34890_/D VGND VGND VPWR VPWR _34890_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33841_ _36085_/CLK _33841_/D VGND VGND VPWR VPWR _33841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18775_ _18661_/X _18773_/X _18774_/X _18665_/X VGND VGND VPWR VPWR _18775_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15987_ _17907_/A VGND VGND VPWR VPWR _15987_/X sky130_fd_sc_hd__buf_4
XFILLER_95_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17726_ _33669_/Q _33605_/Q _33541_/Q _33477_/Q _17553_/X _17554_/X VGND VGND VPWR
+ VPWR _17726_/X sky130_fd_sc_hd__mux4_1
XFILLER_110_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33772_ _34091_/CLK _33772_/D VGND VGND VPWR VPWR _33772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_236_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30984_ _35720_/Q input46/X _31002_/S VGND VGND VPWR VPWR _30985_/A sky130_fd_sc_hd__mux2_1
XTAP_4990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35511_ _35703_/CLK _35511_/D VGND VGND VPWR VPWR _35511_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32723_ _35922_/CLK _32723_/D VGND VGND VPWR VPWR _32723_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17657_ _34179_/Q _34115_/Q _34051_/Q _33987_/Q _17446_/X _17447_/X VGND VGND VPWR
+ VPWR _17657_/X sky130_fd_sc_hd__mux4_1
XFILLER_208_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_223_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16608_ _32869_/Q _32805_/Q _32741_/Q _32677_/Q _16287_/X _16288_/X VGND VGND VPWR
+ VPWR _16608_/X sky130_fd_sc_hd__mux4_1
X_35442_ _35828_/CLK _35442_/D VGND VGND VPWR VPWR _35442_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_6_23__f_CLK clkbuf_5_11_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_23__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_32654_ _36045_/CLK _32654_/D VGND VGND VPWR VPWR _32654_/Q sky130_fd_sc_hd__dfxtp_1
X_17588_ _17588_/A _17588_/B _17588_/C _17588_/D VGND VGND VPWR VPWR _17589_/A sky130_fd_sc_hd__or4_1
XFILLER_211_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19327_ _19153_/X _19323_/X _19326_/X _19156_/X VGND VGND VPWR VPWR _19327_/X sky130_fd_sc_hd__a22o_1
X_31605_ _27717_/X _36014_/Q _31615_/S VGND VGND VPWR VPWR _31606_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35373_ _35566_/CLK _35373_/D VGND VGND VPWR VPWR _35373_/Q sky130_fd_sc_hd__dfxtp_1
X_16539_ _33123_/Q _36003_/Q _32995_/Q _32931_/Q _16356_/X _16357_/X VGND VGND VPWR
+ VPWR _16539_/X sky130_fd_sc_hd__mux4_1
X_32585_ _35978_/CLK _32585_/D VGND VGND VPWR VPWR _32585_/Q sky130_fd_sc_hd__dfxtp_1
X_34324_ _36181_/CLK _34324_/D VGND VGND VPWR VPWR _34324_/Q sky130_fd_sc_hd__dfxtp_1
X_31536_ _31536_/A VGND VGND VPWR VPWR _35981_/D sky130_fd_sc_hd__clkbuf_1
X_19258_ _33135_/Q _36015_/Q _33007_/Q _32943_/Q _19009_/X _19010_/X VGND VGND VPWR
+ VPWR _19258_/X sky130_fd_sc_hd__mux4_1
XFILLER_176_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18209_ _18205_/X _18208_/X _17857_/A VGND VGND VPWR VPWR _18217_/C sky130_fd_sc_hd__o21ba_1
X_34255_ _36175_/CLK _34255_/D VGND VGND VPWR VPWR _34255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19189_ _19153_/X _19187_/X _19188_/X _19156_/X VGND VGND VPWR VPWR _19189_/X sky130_fd_sc_hd__a22o_1
X_31467_ _31467_/A VGND VGND VPWR VPWR _35948_/D sky130_fd_sc_hd__clkbuf_1
X_33206_ _36087_/CLK _33206_/D VGND VGND VPWR VPWR _33206_/Q sky130_fd_sc_hd__dfxtp_1
X_21220_ _34661_/Q _34597_/Q _34533_/Q _34469_/Q _21186_/X _21187_/X VGND VGND VPWR
+ VPWR _21220_/X sky130_fd_sc_hd__mux4_1
XFILLER_89_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30418_ _35452_/Q _29447_/X _30420_/S VGND VGND VPWR VPWR _30419_/A sky130_fd_sc_hd__mux2_1
X_34186_ _34186_/CLK _34186_/D VGND VGND VPWR VPWR _34186_/Q sky130_fd_sc_hd__dfxtp_1
X_31398_ _27810_/X _35916_/Q _31408_/S VGND VGND VPWR VPWR _31399_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21151_ _33059_/Q _32035_/Q _35811_/Q _35747_/Q _20972_/X _20973_/X VGND VGND VPWR
+ VPWR _21151_/X sky130_fd_sc_hd__mux4_1
X_33137_ _36017_/CLK _33137_/D VGND VGND VPWR VPWR _33137_/Q sky130_fd_sc_hd__dfxtp_1
X_30349_ _35419_/Q _29345_/X _30357_/S VGND VGND VPWR VPWR _30350_/A sky130_fd_sc_hd__mux2_1
X_20102_ _19852_/X _20098_/X _20101_/X _19857_/X VGND VGND VPWR VPWR _20102_/X sky130_fd_sc_hd__a22o_1
XFILLER_160_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21082_ _20897_/X _21080_/X _21081_/X _20900_/X VGND VGND VPWR VPWR _21082_/X sky130_fd_sc_hd__a22o_1
X_33068_ _35820_/CLK _33068_/D VGND VGND VPWR VPWR _33068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20033_ _19859_/X _20029_/X _20032_/X _19862_/X VGND VGND VPWR VPWR _20033_/X sky130_fd_sc_hd__a22o_1
XFILLER_28_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24910_ _24910_/A VGND VGND VPWR VPWR _32953_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32019_ _36207_/CLK _32019_/D VGND VGND VPWR VPWR _32019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25890_ _25890_/A VGND VGND VPWR VPWR _33402_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24841_ _24840_/X _32931_/Q _24859_/S VGND VGND VPWR VPWR _24842_/A sky130_fd_sc_hd__mux2_1
XFILLER_246_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27560_ _34160_/Q _27115_/X _27566_/S VGND VGND VPWR VPWR _27561_/A sky130_fd_sc_hd__mux2_1
XTAP_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24772_ _23049_/X _32906_/Q _24786_/S VGND VGND VPWR VPWR _24773_/A sky130_fd_sc_hd__mux2_1
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21984_ _21659_/X _21982_/X _21983_/X _21665_/X VGND VGND VPWR VPWR _21984_/X sky130_fd_sc_hd__a22o_1
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_840 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26511_ _26622_/S VGND VGND VPWR VPWR _26530_/S sky130_fd_sc_hd__buf_4
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23723_ _22909_/X _32349_/Q _23727_/S VGND VGND VPWR VPWR _23724_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35709_ _35709_/CLK _35709_/D VGND VGND VPWR VPWR _35709_/Q sky130_fd_sc_hd__dfxtp_1
X_27491_ _27491_/A VGND VGND VPWR VPWR _34127_/D sky130_fd_sc_hd__clkbuf_1
X_20935_ _20897_/X _20933_/X _20934_/X _20900_/X VGND VGND VPWR VPWR _20935_/X sky130_fd_sc_hd__a22o_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_1025 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26442_ _26442_/A VGND VGND VPWR VPWR _33663_/D sky130_fd_sc_hd__clkbuf_1
X_29230_ _34919_/Q _27087_/X _29234_/S VGND VGND VPWR VPWR _29231_/A sky130_fd_sc_hd__mux2_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23654_ _23702_/S VGND VGND VPWR VPWR _23673_/S sky130_fd_sc_hd__buf_4
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20866_ _20862_/X _20865_/X _20675_/X VGND VGND VPWR VPWR _20874_/C sky130_fd_sc_hd__o21ba_1
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_912 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22605_ _22464_/X _22603_/X _22604_/X _22469_/X VGND VGND VPWR VPWR _22605_/X sky130_fd_sc_hd__a22o_1
X_29161_ _29161_/A VGND VGND VPWR VPWR _34886_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26373_ _33631_/Q _23258_/X _26373_/S VGND VGND VPWR VPWR _26374_/A sky130_fd_sc_hd__mux2_1
X_23585_ _22909_/X _32285_/Q _23589_/S VGND VGND VPWR VPWR _23586_/A sky130_fd_sc_hd__mux2_1
X_20797_ _35417_/Q _35353_/Q _35289_/Q _35225_/Q _20795_/X _20796_/X VGND VGND VPWR
+ VPWR _20797_/X sky130_fd_sc_hd__mux4_1
XFILLER_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28112_ _27639_/X _34390_/Q _28130_/S VGND VGND VPWR VPWR _28113_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25324_ _33135_/Q _23316_/X _25332_/S VGND VGND VPWR VPWR _25325_/A sky130_fd_sc_hd__mux2_1
X_22536_ _22536_/A VGND VGND VPWR VPWR _22536_/X sky130_fd_sc_hd__buf_4
X_29092_ _29092_/A VGND VGND VPWR VPWR _34853_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28043_ _28043_/A VGND VGND VPWR VPWR _34357_/D sky130_fd_sc_hd__clkbuf_1
X_25255_ _33103_/Q _23478_/X _25259_/S VGND VGND VPWR VPWR _25256_/A sky130_fd_sc_hd__mux2_1
X_22467_ _22467_/A VGND VGND VPWR VPWR _22467_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_194_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1083 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24206_ _32639_/Q _23426_/X _24222_/S VGND VGND VPWR VPWR _24207_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_1102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21418_ _21093_/X _21416_/X _21417_/X _21098_/X VGND VGND VPWR VPWR _21418_/X sky130_fd_sc_hd__a22o_1
XFILLER_182_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25186_ _33070_/Q _23305_/X _25196_/S VGND VGND VPWR VPWR _25187_/A sky130_fd_sc_hd__mux2_1
X_22398_ _33671_/Q _33607_/Q _33543_/Q _33479_/Q _22153_/X _22154_/X VGND VGND VPWR
+ VPWR _22398_/X sky130_fd_sc_hd__mux4_1
X_24137_ _24137_/A VGND VGND VPWR VPWR _32606_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21349_ _33129_/Q _36009_/Q _33001_/Q _32937_/Q _21309_/X _21310_/X VGND VGND VPWR
+ VPWR _21349_/X sky130_fd_sc_hd__mux4_1
X_29994_ _35251_/Q _29419_/X _29994_/S VGND VGND VPWR VPWR _29995_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_235_1140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24068_ _23015_/X _32575_/Q _24084_/S VGND VGND VPWR VPWR _24069_/A sky130_fd_sc_hd__mux2_1
X_28945_ _29056_/S VGND VGND VPWR VPWR _28964_/S sky130_fd_sc_hd__buf_4
XFILLER_85_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23019_ _23018_/X _32064_/Q _23040_/S VGND VGND VPWR VPWR _23020_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28876_ _34751_/Q _27162_/X _28892_/S VGND VGND VPWR VPWR _28877_/A sky130_fd_sc_hd__mux2_1
X_16890_ _16886_/X _16889_/X _16779_/X VGND VGND VPWR VPWR _16914_/A sky130_fd_sc_hd__o21ba_1
XFILLER_1_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_938 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27827_ _27827_/A VGND VGND VPWR VPWR _34257_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18560_ _35675_/Q _32181_/Q _35547_/Q _35483_/Q _18558_/X _18559_/X VGND VGND VPWR
+ VPWR _18560_/X sky130_fd_sc_hd__mux4_1
XTAP_4264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_5_24_0_CLK clkbuf_2_3_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_24_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XTAP_4275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27758_ _27757_/X _34235_/Q _27764_/S VGND VGND VPWR VPWR _27759_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17511_ _17864_/A VGND VGND VPWR VPWR _17511_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_166_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26709_ _33788_/Q _23414_/X _26711_/S VGND VGND VPWR VPWR _26710_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_862 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18491_ _18487_/X _18490_/X _18344_/X _18346_/X VGND VGND VPWR VPWR _18508_/B sky130_fd_sc_hd__o211a_1
XTAP_3574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27689_ input7/X VGND VGND VPWR VPWR _27689_/X sky130_fd_sc_hd__buf_4
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29428_ _29428_/A VGND VGND VPWR VPWR _34997_/D sky130_fd_sc_hd__clkbuf_1
X_17442_ _17438_/X _17441_/X _17165_/X VGND VGND VPWR VPWR _17443_/D sky130_fd_sc_hd__o21ba_1
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_2_CLK clkbuf_leaf_2_CLK/A VGND VGND VPWR VPWR _36065_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_221_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29359_ _29359_/A VGND VGND VPWR VPWR _34975_/D sky130_fd_sc_hd__clkbuf_1
X_17373_ _33659_/Q _33595_/Q _33531_/Q _33467_/Q _17200_/X _17201_/X VGND VGND VPWR
+ VPWR _17373_/X sky130_fd_sc_hd__mux4_1
XFILLER_14_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19112_ _20171_/A VGND VGND VPWR VPWR _19112_/X sky130_fd_sc_hd__buf_2
X_16324_ _33117_/Q _35997_/Q _32989_/Q _32925_/Q _16024_/X _16025_/X VGND VGND VPWR
+ VPWR _16324_/X sky130_fd_sc_hd__mux4_1
XFILLER_203_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32370_ _35955_/CLK _32370_/D VGND VGND VPWR VPWR _32370_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16255_ _32859_/Q _32795_/Q _32731_/Q _32667_/Q _16037_/X _16039_/X VGND VGND VPWR
+ VPWR _16255_/X sky130_fd_sc_hd__mux4_1
XFILLER_173_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19043_ _18793_/X _19039_/X _19042_/X _18798_/X VGND VGND VPWR VPWR _19043_/X sky130_fd_sc_hd__a22o_1
X_31321_ _31321_/A VGND VGND VPWR VPWR _35879_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31252_ _27794_/X _35847_/Q _31252_/S VGND VGND VPWR VPWR _31253_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34040_ _35320_/CLK _34040_/D VGND VGND VPWR VPWR _34040_/Q sky130_fd_sc_hd__dfxtp_1
X_16186_ _33113_/Q _35993_/Q _32985_/Q _32921_/Q _16024_/X _16025_/X VGND VGND VPWR
+ VPWR _16186_/X sky130_fd_sc_hd__mux4_1
XFILLER_127_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput206 _36239_/Q VGND VGND VPWR VPWR D2[57] sky130_fd_sc_hd__buf_2
XFILLER_177_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput217 _36191_/Q VGND VGND VPWR VPWR D2[9] sky130_fd_sc_hd__buf_2
XFILLER_177_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30203_ _30335_/S VGND VGND VPWR VPWR _30222_/S sky130_fd_sc_hd__buf_6
XFILLER_127_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput228 _32425_/Q VGND VGND VPWR VPWR D3[19] sky130_fd_sc_hd__buf_2
XFILLER_47_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31183_ _27692_/X _35814_/Q _31189_/S VGND VGND VPWR VPWR _31184_/A sky130_fd_sc_hd__mux2_1
Xoutput239 _32435_/Q VGND VGND VPWR VPWR D3[29] sky130_fd_sc_hd__buf_2
XFILLER_99_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30134_ _35317_/Q _29426_/X _30150_/S VGND VGND VPWR VPWR _30135_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19945_ _20298_/A VGND VGND VPWR VPWR _19945_/X sky130_fd_sc_hd__buf_6
XFILLER_142_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35991_ _35992_/CLK _35991_/D VGND VGND VPWR VPWR _35991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_218_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34942_ _34942_/CLK _34942_/D VGND VGND VPWR VPWR _34942_/Q sky130_fd_sc_hd__dfxtp_1
X_30065_ _35285_/Q _29524_/X _30065_/S VGND VGND VPWR VPWR _30066_/A sky130_fd_sc_hd__mux2_1
X_19876_ _33088_/Q _32064_/Q _35840_/Q _35776_/Q _19731_/X _19732_/X VGND VGND VPWR
+ VPWR _19876_/X sky130_fd_sc_hd__mux4_1
XFILLER_67_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18827_ _18752_/X _18825_/X _18826_/X _18757_/X VGND VGND VPWR VPWR _18827_/X sky130_fd_sc_hd__a22o_1
X_34873_ _36153_/CLK _34873_/D VGND VGND VPWR VPWR _34873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33824_ _36065_/CLK _33824_/D VGND VGND VPWR VPWR _33824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18758_ _18752_/X _18753_/X _18756_/X _18757_/X VGND VGND VPWR VPWR _18758_/X sky130_fd_sc_hd__a22o_1
XFILLER_209_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17709_ _17864_/A VGND VGND VPWR VPWR _17709_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_188_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33755_ _35547_/CLK _33755_/D VGND VGND VPWR VPWR _33755_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30967_ _35712_/Q input37/X _30981_/S VGND VGND VPWR VPWR _30968_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18689_ _34143_/Q _34079_/Q _34015_/Q _33951_/Q _18687_/X _18688_/X VGND VGND VPWR
+ VPWR _18689_/X sky130_fd_sc_hd__mux4_1
XFILLER_93_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20720_ _32087_/Q _32279_/Q _32343_/Q _35863_/Q _20632_/X _22467_/A VGND VGND VPWR
+ VPWR _20720_/X sky130_fd_sc_hd__mux4_1
X_32706_ _32894_/CLK _32706_/D VGND VGND VPWR VPWR _32706_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33686_ _35674_/CLK _33686_/D VGND VGND VPWR VPWR _33686_/Q sky130_fd_sc_hd__dfxtp_1
X_30898_ _30898_/A VGND VGND VPWR VPWR _35679_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35425_ _35810_/CLK _35425_/D VGND VGND VPWR VPWR _35425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20651_ _35670_/Q _32175_/Q _35542_/Q _35478_/Q _20649_/X _20650_/X VGND VGND VPWR
+ VPWR _20651_/X sky130_fd_sc_hd__mux4_1
X_32637_ _35451_/CLK _32637_/D VGND VGND VPWR VPWR _32637_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35356_ _35804_/CLK _35356_/D VGND VGND VPWR VPWR _35356_/Q sky130_fd_sc_hd__dfxtp_1
X_23370_ _23370_/A VGND VGND VPWR VPWR _32200_/D sky130_fd_sc_hd__clkbuf_1
X_20582_ input71/X VGND VGND VPWR VPWR _20661_/A sky130_fd_sc_hd__buf_8
X_32568_ _35961_/CLK _32568_/D VGND VGND VPWR VPWR _32568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22321_ _34948_/Q _34884_/Q _34820_/Q _34756_/Q _22113_/X _22114_/X VGND VGND VPWR
+ VPWR _22321_/X sky130_fd_sc_hd__mux4_1
X_34307_ _36164_/CLK _34307_/D VGND VGND VPWR VPWR _34307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31519_ _31519_/A VGND VGND VPWR VPWR _35973_/D sky130_fd_sc_hd__clkbuf_1
X_35287_ _35799_/CLK _35287_/D VGND VGND VPWR VPWR _35287_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32499_ _36017_/CLK _32499_/D VGND VGND VPWR VPWR _32499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25040_ _25130_/S VGND VGND VPWR VPWR _25059_/S sky130_fd_sc_hd__buf_4
X_22252_ _22111_/X _22250_/X _22251_/X _22116_/X VGND VGND VPWR VPWR _22252_/X sky130_fd_sc_hd__a22o_1
X_34238_ _35071_/CLK _34238_/D VGND VGND VPWR VPWR _34238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21203_ _21199_/X _21202_/X _21026_/X VGND VGND VPWR VPWR _21227_/A sky130_fd_sc_hd__o21ba_1
XFILLER_156_1414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22183_ _22536_/A VGND VGND VPWR VPWR _22183_/X sky130_fd_sc_hd__buf_4
X_34169_ _35641_/CLK _34169_/D VGND VGND VPWR VPWR _34169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21134_ _33379_/Q _33315_/Q _33251_/Q _33187_/Q _21021_/X _21022_/X VGND VGND VPWR
+ VPWR _21134_/X sky130_fd_sc_hd__mux4_1
X_26991_ _26991_/A VGND VGND VPWR VPWR _33921_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28730_ _34683_/Q _27149_/X _28734_/S VGND VGND VPWR VPWR _28731_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25942_ _25942_/A VGND VGND VPWR VPWR _33427_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21065_ _20740_/X _21063_/X _21064_/X _20745_/X VGND VGND VPWR VPWR _21065_/X sky130_fd_sc_hd__a22o_1
XFILLER_219_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20016_ _20016_/A VGND VGND VPWR VPWR _20016_/X sky130_fd_sc_hd__buf_6
XFILLER_100_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28661_ _34650_/Q _27047_/X _28671_/S VGND VGND VPWR VPWR _28662_/A sky130_fd_sc_hd__mux2_1
XFILLER_189_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25873_ _25873_/A VGND VGND VPWR VPWR _33394_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27612_ _27612_/A VGND VGND VPWR VPWR _34184_/D sky130_fd_sc_hd__clkbuf_1
X_24824_ input63/X VGND VGND VPWR VPWR _24824_/X sky130_fd_sc_hd__buf_2
XFILLER_74_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28592_ _27754_/X _34618_/Q _28598_/S VGND VGND VPWR VPWR _28593_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24755_ _23024_/X _32898_/Q _24765_/S VGND VGND VPWR VPWR _24756_/A sky130_fd_sc_hd__mux2_1
X_27543_ _34152_/Q _27090_/X _27545_/S VGND VGND VPWR VPWR _27544_/A sky130_fd_sc_hd__mux2_1
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21967_ _34426_/Q _36154_/Q _34298_/Q _34234_/Q _21829_/X _21830_/X VGND VGND VPWR
+ VPWR _21967_/X sky130_fd_sc_hd__mux4_1
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23706_ _27232_/A _28786_/B VGND VGND VPWR VPWR _27840_/A sky130_fd_sc_hd__nor2_8
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27474_ _27474_/A VGND VGND VPWR VPWR _34119_/D sky130_fd_sc_hd__clkbuf_1
X_20918_ _22450_/A VGND VGND VPWR VPWR _20918_/X sky130_fd_sc_hd__buf_6
XFILLER_42_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24686_ _22922_/X _32865_/Q _24702_/S VGND VGND VPWR VPWR _24687_/A sky130_fd_sc_hd__mux2_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21898_ _34936_/Q _34872_/Q _34808_/Q _34744_/Q _21760_/X _21761_/X VGND VGND VPWR
+ VPWR _21898_/X sky130_fd_sc_hd__mux4_1
XFILLER_187_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29213_ _34911_/Q _27062_/X _29213_/S VGND VGND VPWR VPWR _29214_/A sky130_fd_sc_hd__mux2_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26425_ _26425_/A VGND VGND VPWR VPWR _33655_/D sky130_fd_sc_hd__clkbuf_1
X_23637_ _23637_/A VGND VGND VPWR VPWR _32309_/D sky130_fd_sc_hd__clkbuf_1
X_20849_ _20747_/X _20847_/X _20848_/X _20750_/X VGND VGND VPWR VPWR _20849_/X sky130_fd_sc_hd__a22o_1
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29144_ _34878_/Q _27158_/X _29162_/S VGND VGND VPWR VPWR _29145_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26356_ _26356_/A VGND VGND VPWR VPWR _33622_/D sky130_fd_sc_hd__clkbuf_1
X_23568_ _23568_/A VGND VGND VPWR VPWR _31823_/A sky130_fd_sc_hd__buf_6
XFILLER_195_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25307_ _33127_/Q _23283_/X _25311_/S VGND VGND VPWR VPWR _25308_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22519_ _33162_/Q _36042_/Q _33034_/Q _32970_/Q _22368_/X _22369_/X VGND VGND VPWR
+ VPWR _22519_/X sky130_fd_sc_hd__mux4_1
X_29075_ _29075_/A VGND VGND VPWR VPWR _34845_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_1197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26287_ _26287_/A VGND VGND VPWR VPWR _33590_/D sky130_fd_sc_hd__clkbuf_1
X_23499_ _32245_/Q _23498_/X _23499_/S VGND VGND VPWR VPWR _23500_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16040_ _32854_/Q _32790_/Q _32726_/Q _32662_/Q _16037_/X _16039_/X VGND VGND VPWR
+ VPWR _16040_/X sky130_fd_sc_hd__mux4_1
XFILLER_196_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25238_ _33095_/Q _23450_/X _25238_/S VGND VGND VPWR VPWR _25239_/A sky130_fd_sc_hd__mux2_1
X_28026_ _28026_/A VGND VGND VPWR VPWR _34349_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25169_ _33062_/Q _23280_/X _25175_/S VGND VGND VPWR VPWR _25170_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17991_ _35724_/Q _32235_/Q _35596_/Q _35532_/Q _17670_/X _17671_/X VGND VGND VPWR
+ VPWR _17991_/X sky130_fd_sc_hd__mux4_1
X_29977_ _29977_/A VGND VGND VPWR VPWR _35242_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19730_ _35452_/Q _35388_/Q _35324_/Q _35260_/Q _19554_/X _19555_/X VGND VGND VPWR
+ VPWR _19730_/X sky130_fd_sc_hd__mux4_1
X_28928_ _28928_/A VGND VGND VPWR VPWR _34775_/D sky130_fd_sc_hd__clkbuf_1
X_16942_ _35182_/Q _35118_/Q _35054_/Q _32174_/Q _16657_/X _16658_/X VGND VGND VPWR
+ VPWR _16942_/X sky130_fd_sc_hd__mux4_1
XFILLER_104_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19661_ _19655_/X _19660_/X _19451_/X VGND VGND VPWR VPWR _19671_/C sky130_fd_sc_hd__o21ba_1
XFILLER_238_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28859_ _34743_/Q _27137_/X _28871_/S VGND VGND VPWR VPWR _28860_/A sky130_fd_sc_hd__mux2_1
X_16873_ _34668_/Q _34604_/Q _34540_/Q _34476_/Q _16586_/X _16587_/X VGND VGND VPWR
+ VPWR _16873_/X sky130_fd_sc_hd__mux4_1
XFILLER_93_935 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18612_ _18612_/A _18612_/B _18612_/C _18612_/D VGND VGND VPWR VPWR _18613_/A sky130_fd_sc_hd__or4_1
XTAP_4050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19592_ _20298_/A VGND VGND VPWR VPWR _19592_/X sky130_fd_sc_hd__buf_8
X_31870_ _31870_/A VGND VGND VPWR VPWR _36139_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18543_ _18543_/A VGND VGND VPWR VPWR _32410_/D sky130_fd_sc_hd__clkbuf_4
XTAP_4094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30821_ _35643_/Q input31/X _30825_/S VGND VGND VPWR VPWR _30822_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_810 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33540_ _34182_/CLK _33540_/D VGND VGND VPWR VPWR _33540_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18474_ _18391_/X _18472_/X _18473_/X _18401_/X VGND VGND VPWR VPWR _18474_/X sky130_fd_sc_hd__a22o_1
X_30752_ _35610_/Q input45/X _30762_/S VGND VGND VPWR VPWR _30753_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_1015 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17425_ _17420_/X _17422_/X _17423_/X _17424_/X VGND VGND VPWR VPWR _17425_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33471_ _35453_/CLK _33471_/D VGND VGND VPWR VPWR _33471_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30683_ _30683_/A VGND VGND VPWR VPWR _35577_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35210_ _35210_/CLK _35210_/D VGND VGND VPWR VPWR _35210_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32422_ _36068_/CLK _32422_/D VGND VGND VPWR VPWR _32422_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36190_ _36205_/CLK _36190_/D VGND VGND VPWR VPWR _36190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17356_ _17864_/A VGND VGND VPWR VPWR _17356_/X sky130_fd_sc_hd__buf_4
XFILLER_144_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16307_ _16078_/X _16303_/X _16306_/X _16088_/X VGND VGND VPWR VPWR _16307_/X sky130_fd_sc_hd__a22o_1
X_35141_ _35718_/CLK _35141_/D VGND VGND VPWR VPWR _35141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32353_ _35875_/CLK _32353_/D VGND VGND VPWR VPWR _32353_/Q sky130_fd_sc_hd__dfxtp_1
X_17287_ _16998_/X _17285_/X _17286_/X _17001_/X VGND VGND VPWR VPWR _17287_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31304_ _31304_/A VGND VGND VPWR VPWR _35871_/D sky130_fd_sc_hd__clkbuf_1
X_19026_ _20236_/A VGND VGND VPWR VPWR _19026_/X sky130_fd_sc_hd__buf_4
X_16238_ _34394_/Q _36122_/Q _34266_/Q _34202_/Q _16170_/X _16171_/X VGND VGND VPWR
+ VPWR _16238_/X sky130_fd_sc_hd__mux4_1
X_35072_ _35715_/CLK _35072_/D VGND VGND VPWR VPWR _35072_/Q sky130_fd_sc_hd__dfxtp_1
X_32284_ _36053_/CLK _32284_/D VGND VGND VPWR VPWR _32284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34023_ _34149_/CLK _34023_/D VGND VGND VPWR VPWR _34023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31235_ _31235_/A VGND VGND VPWR VPWR _35838_/D sky130_fd_sc_hd__clkbuf_1
X_16169_ _16078_/X _16167_/X _16168_/X _16088_/X VGND VGND VPWR VPWR _16169_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31166_ _27667_/X _35806_/Q _31168_/S VGND VGND VPWR VPWR _31167_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19928_ _19924_/X _19927_/X _19785_/X VGND VGND VPWR VPWR _19954_/A sky130_fd_sc_hd__o21ba_1
X_30117_ _35309_/Q _29401_/X _30129_/S VGND VGND VPWR VPWR _30118_/A sky130_fd_sc_hd__mux2_1
X_31097_ _31145_/S VGND VGND VPWR VPWR _31116_/S sky130_fd_sc_hd__buf_4
X_35974_ _35974_/CLK _35974_/D VGND VGND VPWR VPWR _35974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30048_ _30048_/A VGND VGND VPWR VPWR _35276_/D sky130_fd_sc_hd__clkbuf_1
X_34925_ _35566_/CLK _34925_/D VGND VGND VPWR VPWR _34925_/Q sky130_fd_sc_hd__dfxtp_1
X_19859_ _20212_/A VGND VGND VPWR VPWR _19859_/X sky130_fd_sc_hd__buf_4
XFILLER_56_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_229_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_1388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22870_ _34709_/Q _34645_/Q _34581_/Q _34517_/Q _22598_/X _22599_/X VGND VGND VPWR
+ VPWR _22870_/X sky130_fd_sc_hd__mux4_1
X_34856_ _34920_/CLK _34856_/D VGND VGND VPWR VPWR _34856_/Q sky130_fd_sc_hd__dfxtp_1
X_33807_ _36113_/CLK _33807_/D VGND VGND VPWR VPWR _33807_/Q sky130_fd_sc_hd__dfxtp_1
X_21821_ _21598_/X _21819_/X _21820_/X _21601_/X VGND VGND VPWR VPWR _21821_/X sky130_fd_sc_hd__a22o_1
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34787_ _34918_/CLK _34787_/D VGND VGND VPWR VPWR _34787_/Q sky130_fd_sc_hd__dfxtp_1
X_31999_ _36207_/CLK _31999_/D VGND VGND VPWR VPWR _31999_/Q sky130_fd_sc_hd__dfxtp_1
X_24540_ _22906_/X _32796_/Q _24546_/S VGND VGND VPWR VPWR _24541_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_1426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33738_ _35210_/CLK _33738_/D VGND VGND VPWR VPWR _33738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21752_ _21747_/X _21750_/X _21751_/X VGND VGND VPWR VPWR _21767_/C sky130_fd_sc_hd__o21ba_1
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20703_ input76/X input75/X VGND VGND VPWR VPWR _22471_/A sky130_fd_sc_hd__or2b_4
X_24471_ _24471_/A VGND VGND VPWR VPWR _32763_/D sky130_fd_sc_hd__clkbuf_1
X_33669_ _34179_/CLK _33669_/D VGND VGND VPWR VPWR _33669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21683_ _34674_/Q _34610_/Q _34546_/Q _34482_/Q _21539_/X _21540_/X VGND VGND VPWR
+ VPWR _21683_/X sky130_fd_sc_hd__mux4_1
XFILLER_196_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26210_ _26210_/A VGND VGND VPWR VPWR _33554_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35408_ _35729_/CLK _35408_/D VGND VGND VPWR VPWR _35408_/Q sky130_fd_sc_hd__dfxtp_1
X_23422_ _32219_/Q _23420_/X _23451_/S VGND VGND VPWR VPWR _23423_/A sky130_fd_sc_hd__mux2_1
X_27190_ _27230_/S VGND VGND VPWR VPWR _27218_/S sky130_fd_sc_hd__buf_4
X_20634_ _22374_/A VGND VGND VPWR VPWR _22467_/A sky130_fd_sc_hd__buf_8
XFILLER_177_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26141_ _26141_/A VGND VGND VPWR VPWR _33521_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35339_ _35852_/CLK _35339_/D VGND VGND VPWR VPWR _35339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23353_ _32193_/Q _23280_/X _23359_/S VGND VGND VPWR VPWR _23354_/A sky130_fd_sc_hd__mux2_1
X_20565_ _18281_/X _20563_/X _20564_/X _18291_/X VGND VGND VPWR VPWR _20565_/X sky130_fd_sc_hd__a22o_1
XFILLER_126_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22304_ _22459_/A VGND VGND VPWR VPWR _22304_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_137_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26072_ _24982_/X _33489_/Q _26072_/S VGND VGND VPWR VPWR _26073_/A sky130_fd_sc_hd__mux2_1
X_23284_ _32167_/Q _23283_/X _23290_/S VGND VGND VPWR VPWR _23285_/A sky130_fd_sc_hd__mux2_1
X_20496_ _32659_/Q _32595_/Q _32531_/Q _35987_/Q _20282_/X _19177_/A VGND VGND VPWR
+ VPWR _20496_/X sky130_fd_sc_hd__mux4_1
X_29900_ _29900_/A VGND VGND VPWR VPWR _35206_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25023_ _25023_/A VGND VGND VPWR VPWR _32993_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22235_ _32898_/Q _32834_/Q _32770_/Q _32706_/Q _21946_/X _21947_/X VGND VGND VPWR
+ VPWR _22235_/X sky130_fd_sc_hd__mux4_1
XFILLER_69_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29831_ _29831_/A VGND VGND VPWR VPWR _35173_/D sky130_fd_sc_hd__clkbuf_1
X_22166_ _33152_/Q _36032_/Q _33024_/Q _32960_/Q _22015_/X _22016_/X VGND VGND VPWR
+ VPWR _22166_/X sky130_fd_sc_hd__mux4_1
XFILLER_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21117_ _33058_/Q _32034_/Q _35810_/Q _35746_/Q _20972_/X _20973_/X VGND VGND VPWR
+ VPWR _21117_/X sky130_fd_sc_hd__mux4_1
X_29762_ _35141_/Q _29475_/X _29766_/S VGND VGND VPWR VPWR _29763_/A sky130_fd_sc_hd__mux2_1
XTAP_6958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22097_ _22450_/A VGND VGND VPWR VPWR _22097_/X sky130_fd_sc_hd__buf_6
X_26974_ _26974_/A VGND VGND VPWR VPWR _33913_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28713_ _34675_/Q _27124_/X _28713_/S VGND VGND VPWR VPWR _28714_/A sky130_fd_sc_hd__mux2_1
X_25925_ _24964_/X _33419_/Q _25937_/S VGND VGND VPWR VPWR _25926_/A sky130_fd_sc_hd__mux2_1
X_21048_ _34656_/Q _34592_/Q _34528_/Q _34464_/Q _20833_/X _20834_/X VGND VGND VPWR
+ VPWR _21048_/X sky130_fd_sc_hd__mux4_1
X_29693_ _35108_/Q _29373_/X _29703_/S VGND VGND VPWR VPWR _29694_/A sky130_fd_sc_hd__mux2_1
XFILLER_232_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28644_ _27831_/X _34643_/Q _28648_/S VGND VGND VPWR VPWR _28645_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25856_ _24861_/X _33386_/Q _25874_/S VGND VGND VPWR VPWR _25857_/A sky130_fd_sc_hd__mux2_1
XFILLER_219_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24807_ _24806_/X _32920_/Q _24828_/S VGND VGND VPWR VPWR _24808_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_873 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28575_ _27729_/X _34610_/Q _28577_/S VGND VGND VPWR VPWR _28576_/A sky130_fd_sc_hd__mux2_1
X_25787_ _25787_/A VGND VGND VPWR VPWR _33353_/D sky130_fd_sc_hd__clkbuf_1
X_22999_ input30/X VGND VGND VPWR VPWR _22999_/X sky130_fd_sc_hd__buf_2
XFILLER_27_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27526_ _27637_/S VGND VGND VPWR VPWR _27545_/S sky130_fd_sc_hd__buf_6
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24738_ _22999_/X _32890_/Q _24744_/S VGND VGND VPWR VPWR _24739_/A sky130_fd_sc_hd__mux2_1
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24669_ _22897_/X _32857_/Q _24681_/S VGND VGND VPWR VPWR _24670_/A sky130_fd_sc_hd__mux2_1
X_27457_ _34111_/Q _27162_/X _27473_/S VGND VGND VPWR VPWR _27458_/A sky130_fd_sc_hd__mux2_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17210_ _17206_/X _17207_/X _17208_/X _17209_/X VGND VGND VPWR VPWR _17210_/X sky130_fd_sc_hd__a22o_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26408_ _26408_/A VGND VGND VPWR VPWR _33647_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18190_ _34195_/Q _34131_/Q _34067_/Q _34003_/Q _16049_/X _16050_/X VGND VGND VPWR
+ VPWR _18190_/X sky130_fd_sc_hd__mux4_1
X_27388_ _27388_/A VGND VGND VPWR VPWR _34078_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_559 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29127_ _34870_/Q _27134_/X _29141_/S VGND VGND VPWR VPWR _29128_/A sky130_fd_sc_hd__mux2_1
X_17141_ _17847_/A VGND VGND VPWR VPWR _17141_/X sky130_fd_sc_hd__clkbuf_4
X_26339_ _26339_/A VGND VGND VPWR VPWR _33615_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17072_ _17067_/X _17069_/X _17070_/X _17071_/X VGND VGND VPWR VPWR _17072_/X sky130_fd_sc_hd__a22o_1
X_29058_ _30202_/A _29797_/A VGND VGND VPWR VPWR _29191_/S sky130_fd_sc_hd__nor2_8
XFILLER_13_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16023_ _32598_/Q _32534_/Q _32470_/Q _35926_/Q _17866_/A _17717_/A VGND VGND VPWR
+ VPWR _16023_/X sky130_fd_sc_hd__mux4_1
XFILLER_13_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28009_ _28009_/A VGND VGND VPWR VPWR _34341_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31020_ _35737_/Q input34/X _31032_/S VGND VGND VPWR VPWR _31021_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_848 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17974_ _17974_/A VGND VGND VPWR VPWR _32011_/D sky130_fd_sc_hd__clkbuf_4
X_19713_ _20066_/A VGND VGND VPWR VPWR _19713_/X sky130_fd_sc_hd__buf_4
X_16925_ _33134_/Q _36014_/Q _33006_/Q _32942_/Q _16709_/X _16710_/X VGND VGND VPWR
+ VPWR _16925_/X sky130_fd_sc_hd__mux4_1
X_32971_ _36044_/CLK _32971_/D VGND VGND VPWR VPWR _32971_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34710_ _34904_/CLK _34710_/D VGND VGND VPWR VPWR _34710_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_293_CLK clkbuf_6_56__f_CLK/X VGND VGND VPWR VPWR _35970_/CLK sky130_fd_sc_hd__clkbuf_16
X_31922_ _31922_/A VGND VGND VPWR VPWR _36164_/D sky130_fd_sc_hd__clkbuf_1
X_19644_ _19359_/X _19642_/X _19643_/X _19365_/X VGND VGND VPWR VPWR _19644_/X sky130_fd_sc_hd__a22o_1
X_35690_ _35690_/CLK _35690_/D VGND VGND VPWR VPWR _35690_/Q sky130_fd_sc_hd__dfxtp_1
X_16856_ _17915_/A VGND VGND VPWR VPWR _16856_/X sky130_fd_sc_hd__buf_4
XFILLER_38_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34641_ _34705_/CLK _34641_/D VGND VGND VPWR VPWR _34641_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19575_ _19571_/X _19574_/X _19432_/X VGND VGND VPWR VPWR _19601_/A sky130_fd_sc_hd__o21ba_1
XFILLER_37_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31853_ _31853_/A VGND VGND VPWR VPWR _36131_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_884 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16787_ _17846_/A VGND VGND VPWR VPWR _16787_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_225_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18526_ _35674_/Q _32180_/Q _35546_/Q _35482_/Q _18349_/X _18350_/X VGND VGND VPWR
+ VPWR _18526_/X sky130_fd_sc_hd__mux4_1
X_30804_ _35635_/Q input22/X _30804_/S VGND VGND VPWR VPWR _30805_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34572_ _36173_/CLK _34572_/D VGND VGND VPWR VPWR _34572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31784_ _36099_/Q input40/X _31792_/S VGND VGND VPWR VPWR _31785_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33523_ _34098_/CLK _33523_/D VGND VGND VPWR VPWR _33523_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_233_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_221_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18457_ _32856_/Q _32792_/Q _32728_/Q _32664_/Q _18337_/X _18339_/X VGND VGND VPWR
+ VPWR _18457_/X sky130_fd_sc_hd__mux4_1
X_30735_ _30735_/A VGND VGND VPWR VPWR _35602_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36242_ _36242_/CLK _36242_/D VGND VGND VPWR VPWR _36242_/Q sky130_fd_sc_hd__dfxtp_1
X_17408_ _33404_/Q _33340_/Q _33276_/Q _33212_/Q _17127_/X _17128_/X VGND VGND VPWR
+ VPWR _17408_/X sky130_fd_sc_hd__mux4_1
X_33454_ _35630_/CLK _33454_/D VGND VGND VPWR VPWR _33454_/Q sky130_fd_sc_hd__dfxtp_1
X_18388_ _19456_/A VGND VGND VPWR VPWR _18388_/X sky130_fd_sc_hd__buf_4
XFILLER_21_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30666_ _30666_/A VGND VGND VPWR VPWR _35569_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32405_ _35989_/CLK _32405_/D VGND VGND VPWR VPWR _32405_/Q sky130_fd_sc_hd__dfxtp_1
X_36173_ _36173_/CLK _36173_/D VGND VGND VPWR VPWR _36173_/Q sky130_fd_sc_hd__dfxtp_1
X_17339_ _33914_/Q _33850_/Q _33786_/Q _36090_/Q _17024_/X _17025_/X VGND VGND VPWR
+ VPWR _17339_/X sky130_fd_sc_hd__mux4_1
X_33385_ _35624_/CLK _33385_/D VGND VGND VPWR VPWR _33385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30597_ _35537_/Q _29512_/X _30597_/S VGND VGND VPWR VPWR _30598_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35124_ _35124_/CLK _35124_/D VGND VGND VPWR VPWR _35124_/Q sky130_fd_sc_hd__dfxtp_1
X_32336_ _35921_/CLK _32336_/D VGND VGND VPWR VPWR _32336_/Q sky130_fd_sc_hd__dfxtp_1
X_20350_ _32910_/Q _32846_/Q _32782_/Q _32718_/Q _18284_/X _18287_/X VGND VGND VPWR
+ VPWR _20350_/X sky130_fd_sc_hd__mux4_1
XFILLER_88_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19009_ _20206_/A VGND VGND VPWR VPWR _19009_/X sky130_fd_sc_hd__buf_4
XFILLER_162_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35055_ _35183_/CLK _35055_/D VGND VGND VPWR VPWR _35055_/Q sky130_fd_sc_hd__dfxtp_1
X_20281_ _20277_/X _20280_/X _20138_/X VGND VGND VPWR VPWR _20307_/A sky130_fd_sc_hd__o21ba_2
X_32267_ _35147_/CLK _32267_/D VGND VGND VPWR VPWR _32267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34006_ _34135_/CLK _34006_/D VGND VGND VPWR VPWR _34006_/Q sky130_fd_sc_hd__dfxtp_1
X_22020_ _22512_/A VGND VGND VPWR VPWR _22020_/X sky130_fd_sc_hd__clkbuf_4
X_31218_ _31218_/A VGND VGND VPWR VPWR _35830_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32198_ _35377_/CLK _32198_/D VGND VGND VPWR VPWR _32198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31149_ _31281_/S VGND VGND VPWR VPWR _31168_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_130_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23971_ _23073_/X _32530_/Q _23977_/S VGND VGND VPWR VPWR _23972_/A sky130_fd_sc_hd__mux2_1
XTAP_4819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35957_ _36021_/CLK _35957_/D VGND VGND VPWR VPWR _35957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_284_CLK clkbuf_6_58__f_CLK/X VGND VGND VPWR VPWR _35711_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_96_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25710_ _24846_/X _33317_/Q _25718_/S VGND VGND VPWR VPWR _25711_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_1057 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22922_ input3/X VGND VGND VPWR VPWR _22922_/X sky130_fd_sc_hd__buf_2
X_34908_ _34911_/CLK _34908_/D VGND VGND VPWR VPWR _34908_/Q sky130_fd_sc_hd__dfxtp_1
X_26690_ _33779_/Q _23384_/X _26690_/S VGND VGND VPWR VPWR _26691_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35888_ _35952_/CLK _35888_/D VGND VGND VPWR VPWR _35888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_244_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22853_ _33941_/Q _33877_/Q _33813_/Q _36117_/Q _20662_/X _20664_/X VGND VGND VPWR
+ VPWR _22853_/X sky130_fd_sc_hd__mux4_1
X_25641_ _25641_/A VGND VGND VPWR VPWR _33284_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34839_ _34904_/CLK _34839_/D VGND VGND VPWR VPWR _34839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_232_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21804_ _22510_/A VGND VGND VPWR VPWR _21804_/X sky130_fd_sc_hd__buf_6
X_28360_ _27810_/X _34508_/Q _28370_/S VGND VGND VPWR VPWR _28361_/A sky130_fd_sc_hd__mux2_1
X_25572_ _25572_/A VGND VGND VPWR VPWR _33251_/D sky130_fd_sc_hd__clkbuf_1
X_22784_ _34962_/Q _34898_/Q _34834_/Q _34770_/Q _20683_/X _20685_/X VGND VGND VPWR
+ VPWR _22784_/X sky130_fd_sc_hd__mux4_1
XFILLER_231_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24523_ _24523_/A VGND VGND VPWR VPWR _32788_/D sky130_fd_sc_hd__clkbuf_1
X_27311_ _34042_/Q _27146_/X _27317_/S VGND VGND VPWR VPWR _27312_/A sky130_fd_sc_hd__mux2_1
XFILLER_197_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21735_ _33140_/Q _36020_/Q _33012_/Q _32948_/Q _21662_/X _21663_/X VGND VGND VPWR
+ VPWR _21735_/X sky130_fd_sc_hd__mux4_1
XFILLER_243_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28291_ _27708_/X _34475_/Q _28307_/S VGND VGND VPWR VPWR _28292_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27242_ _34009_/Q _27044_/X _27254_/S VGND VGND VPWR VPWR _27243_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24454_ _24454_/A VGND VGND VPWR VPWR _32755_/D sky130_fd_sc_hd__clkbuf_1
X_21666_ _21659_/X _21661_/X _21664_/X _21665_/X VGND VGND VPWR VPWR _21666_/X sky130_fd_sc_hd__a22o_1
XFILLER_197_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23405_ input29/X VGND VGND VPWR VPWR _23405_/X sky130_fd_sc_hd__buf_4
X_27173_ _27173_/A VGND VGND VPWR VPWR _33986_/D sky130_fd_sc_hd__clkbuf_1
X_20617_ _22365_/A VGND VGND VPWR VPWR _22505_/A sky130_fd_sc_hd__buf_12
XFILLER_177_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24385_ _23076_/X _32723_/Q _24389_/S VGND VGND VPWR VPWR _24386_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21597_ _21591_/X _21596_/X _21387_/X _21388_/X VGND VGND VPWR VPWR _21618_/B sky130_fd_sc_hd__o211a_1
XFILLER_240_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26124_ _26124_/A VGND VGND VPWR VPWR _33513_/D sky130_fd_sc_hd__clkbuf_1
X_23336_ _23336_/A VGND VGND VPWR VPWR _32185_/D sky130_fd_sc_hd__clkbuf_1
X_20548_ _20548_/A VGND VGND VPWR VPWR _32468_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_126_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26055_ _26055_/A VGND VGND VPWR VPWR _33480_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_748 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23267_ _23267_/A VGND VGND VPWR VPWR _32161_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20479_ _20475_/X _20478_/X _20157_/A VGND VGND VPWR VPWR _20487_/C sky130_fd_sc_hd__o21ba_1
XFILLER_238_1352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25006_ _25006_/A VGND VGND VPWR VPWR _32985_/D sky130_fd_sc_hd__clkbuf_1
X_22218_ _22111_/X _22216_/X _22217_/X _22116_/X VGND VGND VPWR VPWR _22218_/X sky130_fd_sc_hd__a22o_1
XTAP_6700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23198_ _23198_/A VGND VGND VPWR VPWR _32136_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_238_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29814_ _29814_/A VGND VGND VPWR VPWR _35165_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22149_ _22145_/X _22148_/X _22118_/X VGND VGND VPWR VPWR _22150_/D sky130_fd_sc_hd__o21ba_1
XFILLER_121_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29745_ _35133_/Q _29450_/X _29745_/S VGND VGND VPWR VPWR _29746_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26957_ _26957_/A VGND VGND VPWR VPWR _33905_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_275_CLK clkbuf_6_59__f_CLK/X VGND VGND VPWR VPWR _36099_/CLK sky130_fd_sc_hd__clkbuf_16
X_16710_ _17907_/A VGND VGND VPWR VPWR _16710_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_235_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25908_ _24939_/X _33411_/Q _25916_/S VGND VGND VPWR VPWR _25909_/A sky130_fd_sc_hd__mux2_1
X_17690_ _17552_/X _17688_/X _17689_/X _17557_/X VGND VGND VPWR VPWR _17690_/X sky130_fd_sc_hd__a22o_1
X_29676_ _35100_/Q _29348_/X _29682_/S VGND VGND VPWR VPWR _29677_/A sky130_fd_sc_hd__mux2_1
X_26888_ _33873_/Q _23484_/X _26888_/S VGND VGND VPWR VPWR _26889_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_1299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28627_ _28627_/A VGND VGND VPWR VPWR _34634_/D sky130_fd_sc_hd__clkbuf_1
X_16641_ _17834_/A VGND VGND VPWR VPWR _16641_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_235_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25839_ _24837_/X _33378_/Q _25853_/S VGND VGND VPWR VPWR _25840_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19360_ _20066_/A VGND VGND VPWR VPWR _19360_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_204_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28558_ _28648_/S VGND VGND VPWR VPWR _28577_/S sky130_fd_sc_hd__buf_4
XFILLER_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16572_ _33124_/Q _36004_/Q _32996_/Q _32932_/Q _16356_/X _16357_/X VGND VGND VPWR
+ VPWR _16572_/X sky130_fd_sc_hd__mux4_1
XFILLER_27_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_779 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18311_ _20261_/A VGND VGND VPWR VPWR _18311_/X sky130_fd_sc_hd__buf_4
XFILLER_231_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27509_ _27509_/A VGND VGND VPWR VPWR _34135_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19291_ _19006_/X _19289_/X _19290_/X _19012_/X VGND VGND VPWR VPWR _19291_/X sky130_fd_sc_hd__a22o_1
X_28489_ _27801_/X _34569_/Q _28505_/S VGND VGND VPWR VPWR _28490_/A sky130_fd_sc_hd__mux2_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18242_ _16048_/X _18240_/X _18241_/X _16058_/X VGND VGND VPWR VPWR _18242_/X sky130_fd_sc_hd__a22o_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30520_ _35500_/Q _29398_/X _30534_/S VGND VGND VPWR VPWR _30521_/A sky130_fd_sc_hd__mux2_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18173_ _35730_/Q _32241_/Q _35602_/Q _35538_/Q _15993_/X _15995_/X VGND VGND VPWR
+ VPWR _18173_/X sky130_fd_sc_hd__mux4_1
X_30451_ _30451_/A VGND VGND VPWR VPWR _35467_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_1226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17124_ _33652_/Q _33588_/Q _33524_/Q _33460_/Q _16847_/X _16848_/X VGND VGND VPWR
+ VPWR _17124_/X sky130_fd_sc_hd__mux4_1
XFILLER_190_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33170_ _36051_/CLK _33170_/D VGND VGND VPWR VPWR _33170_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_1387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30382_ _30382_/A VGND VGND VPWR VPWR _35434_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32121_ _32889_/CLK _32121_/D VGND VGND VPWR VPWR _32121_/Q sky130_fd_sc_hd__dfxtp_1
X_17055_ _33394_/Q _33330_/Q _33266_/Q _33202_/Q _16774_/X _16775_/X VGND VGND VPWR
+ VPWR _17055_/X sky130_fd_sc_hd__mux4_1
X_16006_ _17777_/A VGND VGND VPWR VPWR _17915_/A sky130_fd_sc_hd__buf_12
X_32052_ _35698_/CLK _32052_/D VGND VGND VPWR VPWR _32052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31003_ _31003_/A VGND VGND VPWR VPWR _35729_/D sky130_fd_sc_hd__clkbuf_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35811_ _35812_/CLK _35811_/D VGND VGND VPWR VPWR _35811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_215_1160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17957_ _35723_/Q _32234_/Q _35595_/Q _35531_/Q _17670_/X _17671_/X VGND VGND VPWR
+ VPWR _17957_/X sky130_fd_sc_hd__mux4_1
XFILLER_113_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_874 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_266_CLK clkbuf_6_62__f_CLK/X VGND VGND VPWR VPWR _34815_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_22_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_721 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35742_ _35807_/CLK _35742_/D VGND VGND VPWR VPWR _35742_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16908_ _35181_/Q _35117_/Q _35053_/Q _32173_/Q _16657_/X _16658_/X VGND VGND VPWR
+ VPWR _16908_/X sky130_fd_sc_hd__mux4_1
X_32954_ _35451_/CLK _32954_/D VGND VGND VPWR VPWR _32954_/Q sky130_fd_sc_hd__dfxtp_1
X_17888_ _17884_/X _17887_/X _17846_/X _17847_/X VGND VGND VPWR VPWR _17903_/B sky130_fd_sc_hd__o211a_1
XFILLER_22_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31905_ _31905_/A VGND VGND VPWR VPWR _36156_/D sky130_fd_sc_hd__clkbuf_1
X_19627_ _35193_/Q _35129_/Q _35065_/Q _32249_/Q _19310_/X _19311_/X VGND VGND VPWR
+ VPWR _19627_/X sky130_fd_sc_hd__mux4_1
XFILLER_226_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35673_ _35673_/CLK _35673_/D VGND VGND VPWR VPWR _35673_/Q sky130_fd_sc_hd__dfxtp_1
X_16839_ _16800_/X _16837_/X _16838_/X _16803_/X VGND VGND VPWR VPWR _16839_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32885_ _32885_/CLK _32885_/D VGND VGND VPWR VPWR _32885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34624_ _34690_/CLK _34624_/D VGND VGND VPWR VPWR _34624_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31836_ _31836_/A VGND VGND VPWR VPWR _36123_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19558_ _19303_/X _19556_/X _19557_/X _19306_/X VGND VGND VPWR VPWR _19558_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18509_ _18509_/A VGND VGND VPWR VPWR _32409_/D sky130_fd_sc_hd__clkbuf_4
X_34555_ _34685_/CLK _34555_/D VGND VGND VPWR VPWR _34555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31767_ _36091_/Q input31/X _31771_/S VGND VGND VPWR VPWR _31768_/A sky130_fd_sc_hd__mux2_1
X_19489_ _19485_/X _19488_/X _19451_/X VGND VGND VPWR VPWR _19497_/C sky130_fd_sc_hd__o21ba_1
X_21520_ _33902_/Q _33838_/Q _33774_/Q _36078_/Q _21271_/X _21272_/X VGND VGND VPWR
+ VPWR _21520_/X sky130_fd_sc_hd__mux4_1
X_33506_ _33573_/CLK _33506_/D VGND VGND VPWR VPWR _33506_/Q sky130_fd_sc_hd__dfxtp_1
X_30718_ _35594_/Q _29491_/X _30732_/S VGND VGND VPWR VPWR _30719_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34486_ _36024_/CLK _34486_/D VGND VGND VPWR VPWR _34486_/Q sky130_fd_sc_hd__dfxtp_1
X_31698_ _36058_/Q input45/X _31708_/S VGND VGND VPWR VPWR _31699_/A sky130_fd_sc_hd__mux2_1
X_36225_ _36229_/CLK _36225_/D VGND VGND VPWR VPWR _36225_/Q sky130_fd_sc_hd__dfxtp_1
X_33437_ _36205_/CLK _33437_/D VGND VGND VPWR VPWR _33437_/Q sky130_fd_sc_hd__dfxtp_1
X_21451_ _22510_/A VGND VGND VPWR VPWR _21451_/X sky130_fd_sc_hd__clkbuf_4
X_30649_ _30649_/A VGND VGND VPWR VPWR _35561_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20402_ _33424_/Q _33360_/Q _33296_/Q _33232_/Q _20133_/X _20134_/X VGND VGND VPWR
+ VPWR _20402_/X sky130_fd_sc_hd__mux4_2
XFILLER_193_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36156_ _36157_/CLK _36156_/D VGND VGND VPWR VPWR _36156_/Q sky130_fd_sc_hd__dfxtp_1
X_24170_ _32622_/Q _23305_/X _24180_/S VGND VGND VPWR VPWR _24171_/A sky130_fd_sc_hd__mux2_1
X_33368_ _36057_/CLK _33368_/D VGND VGND VPWR VPWR _33368_/Q sky130_fd_sc_hd__dfxtp_1
X_21382_ _33130_/Q _36010_/Q _33002_/Q _32938_/Q _21309_/X _21310_/X VGND VGND VPWR
+ VPWR _21382_/X sky130_fd_sc_hd__mux4_1
X_35107_ _36210_/CLK _35107_/D VGND VGND VPWR VPWR _35107_/Q sky130_fd_sc_hd__dfxtp_1
X_23121_ _22931_/X _32100_/Q _23131_/S VGND VGND VPWR VPWR _23122_/A sky130_fd_sc_hd__mux2_1
X_20333_ _34445_/Q _36173_/Q _34317_/Q _34253_/Q _20235_/X _20236_/X VGND VGND VPWR
+ VPWR _20333_/X sky130_fd_sc_hd__mux4_1
X_32319_ _32895_/CLK _32319_/D VGND VGND VPWR VPWR _32319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36087_ _36087_/CLK _36087_/D VGND VGND VPWR VPWR _36087_/Q sky130_fd_sc_hd__dfxtp_1
X_33299_ _36180_/CLK _33299_/D VGND VGND VPWR VPWR _33299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35038_ _36223_/CLK _35038_/D VGND VGND VPWR VPWR _35038_/Q sky130_fd_sc_hd__dfxtp_1
X_23052_ input49/X VGND VGND VPWR VPWR _23052_/X sky130_fd_sc_hd__buf_2
X_20264_ _20009_/X _20262_/X _20263_/X _20012_/X VGND VGND VPWR VPWR _20264_/X sky130_fd_sc_hd__a22o_1
XFILLER_162_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22003_ _22003_/A _22003_/B _22003_/C _22003_/D VGND VGND VPWR VPWR _22004_/A sky130_fd_sc_hd__or4_4
XTAP_6029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27860_ _27670_/X _34271_/Q _27860_/S VGND VGND VPWR VPWR _27861_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20195_ _20191_/X _20194_/X _20157_/X VGND VGND VPWR VPWR _20203_/C sky130_fd_sc_hd__o21ba_1
XTAP_5317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26811_ _33836_/Q _23299_/X _26825_/S VGND VGND VPWR VPWR _26812_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27791_ input43/X VGND VGND VPWR VPWR _27791_/X sky130_fd_sc_hd__clkbuf_4
XTAP_4616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_257_CLK clkbuf_6_63__f_CLK/X VGND VGND VPWR VPWR _34942_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29530_ _29530_/A VGND VGND VPWR VPWR _35030_/D sky130_fd_sc_hd__clkbuf_1
X_26742_ _26742_/A VGND VGND VPWR VPWR _33803_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23954_ _23954_/A VGND VGND VPWR VPWR _32521_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22905_ _22905_/A VGND VGND VPWR VPWR _32027_/D sky130_fd_sc_hd__clkbuf_1
X_29461_ _35008_/Q _29460_/X _29482_/S VGND VGND VPWR VPWR _29462_/A sky130_fd_sc_hd__mux2_1
XTAP_3948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26673_ _26673_/A VGND VGND VPWR VPWR _33770_/D sky130_fd_sc_hd__clkbuf_1
X_23885_ _22946_/X _32489_/Q _23885_/S VGND VGND VPWR VPWR _23886_/A sky130_fd_sc_hd__mux2_1
XTAP_3959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1097 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28412_ _28412_/A VGND VGND VPWR VPWR _34532_/D sky130_fd_sc_hd__clkbuf_1
X_22836_ _35476_/Q _35412_/Q _35348_/Q _35284_/Q _22560_/X _22561_/X VGND VGND VPWR
+ VPWR _22836_/X sky130_fd_sc_hd__mux4_1
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25624_ _25624_/A VGND VGND VPWR VPWR _33276_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29392_ _29525_/S VGND VGND VPWR VPWR _29420_/S sky130_fd_sc_hd__buf_4
XFILLER_204_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28343_ _27785_/X _34500_/Q _28349_/S VGND VGND VPWR VPWR _28344_/A sky130_fd_sc_hd__mux2_1
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25555_ _25555_/A VGND VGND VPWR VPWR _33243_/D sky130_fd_sc_hd__clkbuf_1
X_22767_ _33170_/Q _36050_/Q _33042_/Q _32978_/Q _20632_/X _21761_/A VGND VGND VPWR
+ VPWR _22767_/X sky130_fd_sc_hd__mux4_1
XFILLER_25_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1075 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24506_ _23055_/X _32780_/Q _24516_/S VGND VGND VPWR VPWR _24507_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21718_ _34419_/Q _36147_/Q _34291_/Q _34227_/Q _21476_/X _21477_/X VGND VGND VPWR
+ VPWR _21718_/X sky130_fd_sc_hd__mux4_1
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25486_ _24914_/X _33211_/Q _25490_/S VGND VGND VPWR VPWR _25487_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28274_ _27683_/X _34467_/Q _28286_/S VGND VGND VPWR VPWR _28275_/A sky130_fd_sc_hd__mux2_1
X_22698_ _22698_/A VGND VGND VPWR VPWR _36239_/D sky130_fd_sc_hd__clkbuf_1
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27225_ _27225_/A VGND VGND VPWR VPWR _34003_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_240_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21649_ _21645_/X _21648_/X _21412_/X VGND VGND VPWR VPWR _21650_/D sky130_fd_sc_hd__o21ba_1
X_24437_ _22953_/X _32747_/Q _24453_/S VGND VGND VPWR VPWR _24438_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24368_ _24368_/A VGND VGND VPWR VPWR _32714_/D sky130_fd_sc_hd__clkbuf_1
X_27156_ _33981_/Q _27155_/X _27156_/S VGND VGND VPWR VPWR _27157_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23319_ _32177_/Q _23234_/X _23335_/S VGND VGND VPWR VPWR _23320_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26107_ _24834_/X _33505_/Q _26123_/S VGND VGND VPWR VPWR _26108_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27087_ input9/X VGND VGND VPWR VPWR _27087_/X sky130_fd_sc_hd__buf_4
XFILLER_197_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24299_ _24389_/S VGND VGND VPWR VPWR _24318_/S sky130_fd_sc_hd__buf_4
XFILLER_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26038_ _26038_/A VGND VGND VPWR VPWR _33472_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_496_CLK clkbuf_6_2__f_CLK/X VGND VGND VPWR VPWR _33697_/CLK sky130_fd_sc_hd__clkbuf_16
X_18860_ _18856_/X _18859_/X _18759_/X VGND VGND VPWR VPWR _18861_/D sky130_fd_sc_hd__o21ba_1
XTAP_6530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17811_ _32903_/Q _32839_/Q _32775_/Q _32711_/Q _17699_/X _17700_/X VGND VGND VPWR
+ VPWR _17811_/X sky130_fd_sc_hd__mux4_1
XFILLER_239_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18791_ _18791_/A _18791_/B _18791_/C _18791_/D VGND VGND VPWR VPWR _18792_/A sky130_fd_sc_hd__or4_2
XTAP_6585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27989_ _34332_/Q _27053_/X _27995_/S VGND VGND VPWR VPWR _27990_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_248_CLK clkbuf_6_61__f_CLK/X VGND VGND VPWR VPWR _34121_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_6596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17742_ _35717_/Q _32227_/Q _35589_/Q _35525_/Q _17670_/X _17671_/X VGND VGND VPWR
+ VPWR _17742_/X sky130_fd_sc_hd__mux4_1
X_29728_ _29728_/A VGND VGND VPWR VPWR _35124_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29659_ _29659_/A VGND VGND VPWR VPWR _35092_/D sky130_fd_sc_hd__clkbuf_1
X_17673_ _35651_/Q _35011_/Q _34371_/Q _33731_/Q _17497_/X _17498_/X VGND VGND VPWR
+ VPWR _17673_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19412_ _33075_/Q _32051_/Q _35827_/Q _35763_/Q _19378_/X _19379_/X VGND VGND VPWR
+ VPWR _19412_/X sky130_fd_sc_hd__mux4_1
X_16624_ _34917_/Q _34853_/Q _34789_/Q _34725_/Q _16454_/X _16455_/X VGND VGND VPWR
+ VPWR _16624_/X sky130_fd_sc_hd__mux4_1
XFILLER_235_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32670_ _35870_/CLK _32670_/D VGND VGND VPWR VPWR _32670_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19343_ _34673_/Q _34609_/Q _34545_/Q _34481_/Q _19239_/X _19240_/X VGND VGND VPWR
+ VPWR _19343_/X sky130_fd_sc_hd__mux4_1
X_31621_ _31621_/A VGND VGND VPWR VPWR _36021_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16555_ _35171_/Q _35107_/Q _35043_/Q _32163_/Q _16304_/X _16305_/X VGND VGND VPWR
+ VPWR _16555_/X sky130_fd_sc_hd__mux4_1
XFILLER_204_774 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_420_CLK clkbuf_6_33__f_CLK/X VGND VGND VPWR VPWR _34927_/CLK sky130_fd_sc_hd__clkbuf_16
X_34340_ _35620_/CLK _34340_/D VGND VGND VPWR VPWR _34340_/Q sky130_fd_sc_hd__dfxtp_1
X_31552_ _31552_/A VGND VGND VPWR VPWR _35989_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19274_ _35183_/Q _35119_/Q _35055_/Q _32176_/Q _18957_/X _18958_/X VGND VGND VPWR
+ VPWR _19274_/X sky130_fd_sc_hd__mux4_1
XFILLER_56_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16486_ _16447_/X _16484_/X _16485_/X _16450_/X VGND VGND VPWR VPWR _16486_/X sky130_fd_sc_hd__a22o_1
XFILLER_188_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18225_ _18221_/X _18224_/X _17838_/A VGND VGND VPWR VPWR _18247_/A sky130_fd_sc_hd__o21ba_1
X_30503_ _35492_/Q _29373_/X _30513_/S VGND VGND VPWR VPWR _30504_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34271_ _36127_/CLK _34271_/D VGND VGND VPWR VPWR _34271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_1170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31483_ _27735_/X _35956_/Q _31501_/S VGND VGND VPWR VPWR _31484_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36010_ _36010_/CLK _36010_/D VGND VGND VPWR VPWR _36010_/Q sky130_fd_sc_hd__dfxtp_1
X_33222_ _36102_/CLK _33222_/D VGND VGND VPWR VPWR _33222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18156_ _18152_/X _18155_/X _17871_/X VGND VGND VPWR VPWR _18157_/D sky130_fd_sc_hd__o21ba_1
XFILLER_175_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30434_ _30434_/A VGND VGND VPWR VPWR _35459_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17107_ _17103_/X _17106_/X _16787_/X _16788_/X VGND VGND VPWR VPWR _17122_/B sky130_fd_sc_hd__o211a_1
X_33153_ _36033_/CLK _33153_/D VGND VGND VPWR VPWR _33153_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18087_ _33103_/Q _32079_/Q _35855_/Q _35791_/Q _17784_/X _17785_/X VGND VGND VPWR
+ VPWR _18087_/X sky130_fd_sc_hd__mux4_1
X_30365_ _30365_/A VGND VGND VPWR VPWR _35426_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32104_ _32873_/CLK _32104_/D VGND VGND VPWR VPWR _32104_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_887 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17038_ _16998_/X _17036_/X _17037_/X _17001_/X VGND VGND VPWR VPWR _17038_/X sky130_fd_sc_hd__a22o_1
XFILLER_144_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33084_ _35453_/CLK _33084_/D VGND VGND VPWR VPWR _33084_/Q sky130_fd_sc_hd__dfxtp_1
X_30296_ _35394_/Q _29466_/X _30306_/S VGND VGND VPWR VPWR _30297_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_487_CLK _35560_/CLK VGND VGND VPWR VPWR _35690_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_113_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32035_ _35814_/CLK _32035_/D VGND VGND VPWR VPWR _32035_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_6_46__f_CLK clkbuf_5_23_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_46__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18989_ _18985_/X _18988_/X _18745_/X VGND VGND VPWR VPWR _18997_/C sky130_fd_sc_hd__o21ba_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_239_CLK clkbuf_6_60__f_CLK/X VGND VGND VPWR VPWR _36164_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33986_ _34945_/CLK _33986_/D VGND VGND VPWR VPWR _33986_/Q sky130_fd_sc_hd__dfxtp_1
X_35725_ _35727_/CLK _35725_/D VGND VGND VPWR VPWR _35725_/Q sky130_fd_sc_hd__dfxtp_1
X_20951_ _20747_/X _20949_/X _20950_/X _20750_/X VGND VGND VPWR VPWR _20951_/X sky130_fd_sc_hd__a22o_1
XFILLER_38_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32937_ _35755_/CLK _32937_/D VGND VGND VPWR VPWR _32937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_226_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_532 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23670_ _23670_/A VGND VGND VPWR VPWR _32325_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35656_ _35657_/CLK _35656_/D VGND VGND VPWR VPWR _35656_/Q sky130_fd_sc_hd__dfxtp_1
X_20882_ _20878_/X _20881_/X _20615_/X VGND VGND VPWR VPWR _20912_/A sky130_fd_sc_hd__o21ba_1
X_32868_ _32871_/CLK _32868_/D VGND VGND VPWR VPWR _32868_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22621_ _22373_/X _22619_/X _22620_/X _22377_/X VGND VGND VPWR VPWR _22621_/X sky130_fd_sc_hd__a22o_1
X_31819_ _36116_/Q input59/X _31821_/S VGND VGND VPWR VPWR _31820_/A sky130_fd_sc_hd__mux2_1
X_34607_ _36143_/CLK _34607_/D VGND VGND VPWR VPWR _34607_/Q sky130_fd_sc_hd__dfxtp_1
X_35587_ _35655_/CLK _35587_/D VGND VGND VPWR VPWR _35587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32799_ _35870_/CLK _32799_/D VGND VGND VPWR VPWR _32799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_411_CLK clkbuf_6_32__f_CLK/X VGND VGND VPWR VPWR _33393_/CLK sky130_fd_sc_hd__clkbuf_16
X_25340_ _25340_/A VGND VGND VPWR VPWR _33142_/D sky130_fd_sc_hd__clkbuf_1
X_22552_ _22365_/X _22550_/X _22551_/X _22371_/X VGND VGND VPWR VPWR _22552_/X sky130_fd_sc_hd__a22o_1
X_34538_ _35180_/CLK _34538_/D VGND VGND VPWR VPWR _34538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21503_ _35437_/Q _35373_/Q _35309_/Q _35245_/Q _21501_/X _21502_/X VGND VGND VPWR
+ VPWR _21503_/X sky130_fd_sc_hd__mux4_1
XFILLER_210_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25271_ _25403_/S VGND VGND VPWR VPWR _25290_/S sky130_fd_sc_hd__buf_6
X_22483_ _33161_/Q _36041_/Q _33033_/Q _32969_/Q _22368_/X _22369_/X VGND VGND VPWR
+ VPWR _22483_/X sky130_fd_sc_hd__mux4_1
X_34469_ _36136_/CLK _34469_/D VGND VGND VPWR VPWR _34469_/Q sky130_fd_sc_hd__dfxtp_1
X_27010_ _27010_/A VGND VGND VPWR VPWR _33930_/D sky130_fd_sc_hd__clkbuf_1
X_24222_ _32647_/Q _23450_/X _24222_/S VGND VGND VPWR VPWR _24223_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36208_ _36211_/CLK _36208_/D VGND VGND VPWR VPWR _36208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21434_ _33067_/Q _32043_/Q _35819_/Q _35755_/Q _21325_/X _21326_/X VGND VGND VPWR
+ VPWR _21434_/X sky130_fd_sc_hd__mux4_1
XFILLER_194_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36139_ _36140_/CLK _36139_/D VGND VGND VPWR VPWR _36139_/Q sky130_fd_sc_hd__dfxtp_1
X_24153_ _32614_/Q _23280_/X _24159_/S VGND VGND VPWR VPWR _24154_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_1434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21365_ _34409_/Q _36137_/Q _34281_/Q _34217_/Q _21123_/X _21124_/X VGND VGND VPWR
+ VPWR _21365_/X sky130_fd_sc_hd__mux4_1
XFILLER_206_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23104_ _22906_/X _32092_/Q _23110_/S VGND VGND VPWR VPWR _23105_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20316_ _32653_/Q _32589_/Q _32525_/Q _35981_/Q _20282_/X _20066_/X VGND VGND VPWR
+ VPWR _20316_/X sky130_fd_sc_hd__mux4_1
XFILLER_159_1478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24084_ _23039_/X _32583_/Q _24084_/S VGND VGND VPWR VPWR _24085_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28961_ _28961_/A VGND VGND VPWR VPWR _34791_/D sky130_fd_sc_hd__clkbuf_1
X_21296_ _21292_/X _21295_/X _21059_/X VGND VGND VPWR VPWR _21297_/D sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_478_CLK clkbuf_6_10__f_CLK/X VGND VGND VPWR VPWR _36076_/CLK sky130_fd_sc_hd__clkbuf_16
X_23035_ _23035_/A VGND VGND VPWR VPWR _32069_/D sky130_fd_sc_hd__clkbuf_1
X_27912_ _27912_/A VGND VGND VPWR VPWR _34295_/D sky130_fd_sc_hd__clkbuf_1
X_20247_ _33931_/Q _33867_/Q _33803_/Q _36107_/Q _20030_/X _20031_/X VGND VGND VPWR
+ VPWR _20247_/X sky130_fd_sc_hd__mux4_1
X_28892_ _34759_/Q _27186_/X _28892_/S VGND VGND VPWR VPWR _28893_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27843_ _27843_/A VGND VGND VPWR VPWR _34262_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20178_ _33417_/Q _33353_/Q _33289_/Q _33225_/Q _20133_/X _20134_/X VGND VGND VPWR
+ VPWR _20178_/X sky130_fd_sc_hd__mux4_1
XTAP_5136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27774_ _27773_/X _34240_/Q _27795_/S VGND VGND VPWR VPWR _27775_/A sky130_fd_sc_hd__mux2_1
XTAP_4435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24986_ _24985_/X _32978_/Q _24995_/S VGND VGND VPWR VPWR _24987_/A sky130_fd_sc_hd__mux2_1
XTAP_4446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29513_ _35025_/Q _29512_/X _29513_/S VGND VGND VPWR VPWR _29514_/A sky130_fd_sc_hd__mux2_1
XTAP_4457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26725_ _26725_/A VGND VGND VPWR VPWR _33795_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23937_ _23937_/A VGND VGND VPWR VPWR _32513_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29444_ input31/X VGND VGND VPWR VPWR _29444_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_166_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26656_ _26656_/A VGND VGND VPWR VPWR _33762_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23868_ _23868_/A VGND VGND VPWR VPWR _32480_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25607_ _24892_/X _33268_/Q _25625_/S VGND VGND VPWR VPWR _25608_/A sky130_fd_sc_hd__mux2_1
X_22819_ _33684_/Q _33620_/Q _33556_/Q _33492_/Q _20624_/X _20625_/X VGND VGND VPWR
+ VPWR _22819_/X sky130_fd_sc_hd__mux4_1
XFILLER_16_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29375_ _29375_/A VGND VGND VPWR VPWR _34980_/D sky130_fd_sc_hd__clkbuf_1
X_26587_ _24942_/X _33732_/Q _26593_/S VGND VGND VPWR VPWR _26588_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23799_ _23021_/X _32385_/Q _23811_/S VGND VGND VPWR VPWR _23800_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_402_CLK clkbuf_6_34__f_CLK/X VGND VGND VPWR VPWR _35699_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16340_ _34397_/Q _36125_/Q _34269_/Q _34205_/Q _16170_/X _16171_/X VGND VGND VPWR
+ VPWR _16340_/X sky130_fd_sc_hd__mux4_1
X_28326_ _27760_/X _34492_/Q _28328_/S VGND VGND VPWR VPWR _28327_/A sky130_fd_sc_hd__mux2_1
X_25538_ _24991_/X _33236_/Q _25540_/S VGND VGND VPWR VPWR _25539_/A sky130_fd_sc_hd__mux2_1
XFILLER_198_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_974 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_946 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16271_ _34907_/Q _34843_/Q _34779_/Q _34715_/Q _16096_/X _16098_/X VGND VGND VPWR
+ VPWR _16271_/X sky130_fd_sc_hd__mux4_1
X_28257_ _27658_/X _34459_/Q _28265_/S VGND VGND VPWR VPWR _28258_/A sky130_fd_sc_hd__mux2_1
X_25469_ _24889_/X _33203_/Q _25469_/S VGND VGND VPWR VPWR _25470_/A sky130_fd_sc_hd__mux2_1
X_18010_ _34189_/Q _34125_/Q _34061_/Q _33997_/Q _17799_/X _17800_/X VGND VGND VPWR
+ VPWR _18010_/X sky130_fd_sc_hd__mux4_1
XFILLER_139_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27208_ input52/X VGND VGND VPWR VPWR _27208_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_157_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28188_ _28188_/A VGND VGND VPWR VPWR _34426_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27139_ _27139_/A VGND VGND VPWR VPWR _33975_/D sky130_fd_sc_hd__clkbuf_1
X_19961_ _19859_/X _19959_/X _19960_/X _19862_/X VGND VGND VPWR VPWR _19961_/X sky130_fd_sc_hd__a22o_1
XFILLER_180_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30150_ _35325_/Q _29450_/X _30150_/S VGND VGND VPWR VPWR _30151_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18912_ _20100_/A VGND VGND VPWR VPWR _18912_/X sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_469_CLK clkbuf_6_11__f_CLK/X VGND VGND VPWR VPWR _35438_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_7050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19892_ _19852_/X _19890_/X _19891_/X _19857_/X VGND VGND VPWR VPWR _19892_/X sky130_fd_sc_hd__a22o_1
X_30081_ _35292_/Q _29348_/X _30087_/S VGND VGND VPWR VPWR _30082_/A sky130_fd_sc_hd__mux2_1
XTAP_7061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18843_ _18661_/X _18841_/X _18842_/X _18665_/X VGND VGND VPWR VPWR _18843_/X sky130_fd_sc_hd__a22o_1
XFILLER_67_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33840_ _33904_/CLK _33840_/D VGND VGND VPWR VPWR _33840_/Q sky130_fd_sc_hd__dfxtp_1
X_18774_ _32865_/Q _32801_/Q _32737_/Q _32673_/Q _18587_/X _18588_/X VGND VGND VPWR
+ VPWR _18774_/X sky130_fd_sc_hd__mux4_1
X_15986_ _16063_/A VGND VGND VPWR VPWR _17907_/A sky130_fd_sc_hd__buf_12
XTAP_5670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17725_ _17725_/A VGND VGND VPWR VPWR _32004_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_208_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33771_ _33895_/CLK _33771_/D VGND VGND VPWR VPWR _33771_/Q sky130_fd_sc_hd__dfxtp_1
X_30983_ _31010_/S VGND VGND VPWR VPWR _31002_/S sky130_fd_sc_hd__buf_4
XFILLER_180_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32722_ _35922_/CLK _32722_/D VGND VGND VPWR VPWR _32722_/Q sky130_fd_sc_hd__dfxtp_1
X_35510_ _35703_/CLK _35510_/D VGND VGND VPWR VPWR _35510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17656_ _33667_/Q _33603_/Q _33539_/Q _33475_/Q _17553_/X _17554_/X VGND VGND VPWR
+ VPWR _17656_/X sky130_fd_sc_hd__mux4_1
XFILLER_224_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35441_ _35764_/CLK _35441_/D VGND VGND VPWR VPWR _35441_/Q sky130_fd_sc_hd__dfxtp_1
X_16607_ _32101_/Q _32293_/Q _32357_/Q _35877_/Q _16574_/X _16362_/X VGND VGND VPWR
+ VPWR _16607_/X sky130_fd_sc_hd__mux4_1
X_32653_ _32655_/CLK _32653_/D VGND VGND VPWR VPWR _32653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17587_ _17581_/X _17586_/X _17518_/X VGND VGND VPWR VPWR _17588_/D sky130_fd_sc_hd__o21ba_1
XFILLER_23_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19326_ _33905_/Q _33841_/Q _33777_/Q _36081_/Q _19324_/X _19325_/X VGND VGND VPWR
+ VPWR _19326_/X sky130_fd_sc_hd__mux4_1
X_31604_ _31604_/A VGND VGND VPWR VPWR _36013_/D sky130_fd_sc_hd__clkbuf_1
X_35372_ _35691_/CLK _35372_/D VGND VGND VPWR VPWR _35372_/Q sky130_fd_sc_hd__dfxtp_1
X_16538_ _32611_/Q _32547_/Q _32483_/Q _35939_/Q _16217_/X _16354_/X VGND VGND VPWR
+ VPWR _16538_/X sky130_fd_sc_hd__mux4_1
X_32584_ _35976_/CLK _32584_/D VGND VGND VPWR VPWR _32584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34323_ _34963_/CLK _34323_/D VGND VGND VPWR VPWR _34323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31535_ _27813_/X _35981_/Q _31543_/S VGND VGND VPWR VPWR _31536_/A sky130_fd_sc_hd__mux2_1
X_19257_ _32623_/Q _32559_/Q _32495_/Q _35951_/Q _19223_/X _19007_/X VGND VGND VPWR
+ VPWR _19257_/X sky130_fd_sc_hd__mux4_1
X_16469_ _16465_/X _16468_/X _16426_/X VGND VGND VPWR VPWR _16491_/A sky130_fd_sc_hd__o21ba_1
XFILLER_148_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18208_ _16001_/X _18206_/X _18207_/X _16007_/X VGND VGND VPWR VPWR _18208_/X sky130_fd_sc_hd__a22o_1
X_34254_ _36176_/CLK _34254_/D VGND VGND VPWR VPWR _34254_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19188_ _33901_/Q _33837_/Q _33773_/Q _36077_/Q _18971_/X _18972_/X VGND VGND VPWR
+ VPWR _19188_/X sky130_fd_sc_hd__mux4_1
X_31466_ _27711_/X _35948_/Q _31480_/S VGND VGND VPWR VPWR _31467_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33205_ _34100_/CLK _33205_/D VGND VGND VPWR VPWR _33205_/Q sky130_fd_sc_hd__dfxtp_1
X_18139_ _32145_/Q _32337_/Q _32401_/Q _35921_/Q _17986_/X _17011_/A VGND VGND VPWR
+ VPWR _18139_/X sky130_fd_sc_hd__mux4_1
X_30417_ _30417_/A VGND VGND VPWR VPWR _35451_/D sky130_fd_sc_hd__clkbuf_1
X_34185_ _34185_/CLK _34185_/D VGND VGND VPWR VPWR _34185_/Q sky130_fd_sc_hd__dfxtp_1
X_31397_ _31397_/A VGND VGND VPWR VPWR _35915_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21150_ _35427_/Q _35363_/Q _35299_/Q _35235_/Q _21148_/X _21149_/X VGND VGND VPWR
+ VPWR _21150_/X sky130_fd_sc_hd__mux4_1
X_33136_ _36144_/CLK _33136_/D VGND VGND VPWR VPWR _33136_/Q sky130_fd_sc_hd__dfxtp_1
X_30348_ _30348_/A VGND VGND VPWR VPWR _35418_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20101_ _34183_/Q _34119_/Q _34055_/Q _33991_/Q _20099_/X _20100_/X VGND VGND VPWR
+ VPWR _20101_/X sky130_fd_sc_hd__mux4_1
XFILLER_208_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33067_ _35820_/CLK _33067_/D VGND VGND VPWR VPWR _33067_/Q sky130_fd_sc_hd__dfxtp_1
X_21081_ _33057_/Q _32033_/Q _35809_/Q _35745_/Q _20972_/X _20973_/X VGND VGND VPWR
+ VPWR _21081_/X sky130_fd_sc_hd__mux4_1
XFILLER_193_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30279_ _35386_/Q _29441_/X _30285_/S VGND VGND VPWR VPWR _30280_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20032_ _33925_/Q _33861_/Q _33797_/Q _36101_/Q _20030_/X _20031_/X VGND VGND VPWR
+ VPWR _20032_/X sky130_fd_sc_hd__mux4_1
X_32018_ _36207_/CLK _32018_/D VGND VGND VPWR VPWR _32018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24840_ input5/X VGND VGND VPWR VPWR _24840_/X sky130_fd_sc_hd__buf_4
XFILLER_37_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_979 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24771_ _24771_/A VGND VGND VPWR VPWR _32905_/D sky130_fd_sc_hd__clkbuf_1
X_21983_ _33147_/Q _36027_/Q _33019_/Q _32955_/Q _21662_/X _21663_/X VGND VGND VPWR
+ VPWR _21983_/X sky130_fd_sc_hd__mux4_1
XFILLER_27_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33969_ _35632_/CLK _33969_/D VGND VGND VPWR VPWR _33969_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26510_ _26510_/A VGND VGND VPWR VPWR _33695_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23722_ _23722_/A VGND VGND VPWR VPWR _32348_/D sky130_fd_sc_hd__clkbuf_1
X_20934_ _33053_/Q _32029_/Q _35805_/Q _35741_/Q _20667_/X _20669_/X VGND VGND VPWR
+ VPWR _20934_/X sky130_fd_sc_hd__mux4_1
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35708_ _35708_/CLK _35708_/D VGND VGND VPWR VPWR _35708_/Q sky130_fd_sc_hd__dfxtp_1
X_27490_ _34127_/Q _27211_/X _27494_/S VGND VGND VPWR VPWR _27491_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26441_ _33663_/Q _23426_/X _26457_/S VGND VGND VPWR VPWR _26442_/A sky130_fd_sc_hd__mux2_1
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20865_ _20660_/X _20863_/X _20864_/X _20672_/X VGND VGND VPWR VPWR _20865_/X sky130_fd_sc_hd__a22o_1
X_23653_ _23653_/A VGND VGND VPWR VPWR _32317_/D sky130_fd_sc_hd__clkbuf_1
X_35639_ _35768_/CLK _35639_/D VGND VGND VPWR VPWR _35639_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22604_ _34956_/Q _34892_/Q _34828_/Q _34764_/Q _22466_/X _22467_/X VGND VGND VPWR
+ VPWR _22604_/X sky130_fd_sc_hd__mux4_1
XFILLER_223_880 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29160_ _34886_/Q _27183_/X _29162_/S VGND VGND VPWR VPWR _29161_/A sky130_fd_sc_hd__mux2_1
X_23584_ _23584_/A VGND VGND VPWR VPWR _32284_/D sky130_fd_sc_hd__clkbuf_1
X_26372_ _26372_/A VGND VGND VPWR VPWR _33630_/D sky130_fd_sc_hd__clkbuf_1
X_20796_ _22451_/A VGND VGND VPWR VPWR _20796_/X sky130_fd_sc_hd__buf_4
X_28111_ _28243_/S VGND VGND VPWR VPWR _28130_/S sky130_fd_sc_hd__buf_4
X_22535_ _22535_/A VGND VGND VPWR VPWR _22535_/X sky130_fd_sc_hd__buf_6
XFILLER_179_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25323_ _25323_/A VGND VGND VPWR VPWR _33134_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29091_ _34853_/Q _27081_/X _29099_/S VGND VGND VPWR VPWR _29092_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28042_ _34357_/Q _27131_/X _28058_/S VGND VGND VPWR VPWR _28043_/A sky130_fd_sc_hd__mux2_1
X_22466_ _22466_/A VGND VGND VPWR VPWR _22466_/X sky130_fd_sc_hd__buf_4
X_25254_ _25254_/A VGND VGND VPWR VPWR _33102_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_241_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24205_ _24205_/A VGND VGND VPWR VPWR _32638_/D sky130_fd_sc_hd__clkbuf_1
X_21417_ _34155_/Q _34091_/Q _34027_/Q _33963_/Q _21340_/X _21341_/X VGND VGND VPWR
+ VPWR _21417_/X sky130_fd_sc_hd__mux4_1
XFILLER_33_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25185_ _25185_/A VGND VGND VPWR VPWR _33069_/D sky130_fd_sc_hd__clkbuf_1
X_22397_ _22397_/A VGND VGND VPWR VPWR _36230_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24136_ _32606_/Q _23255_/X _24138_/S VGND VGND VPWR VPWR _24137_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21348_ _32617_/Q _32553_/Q _32489_/Q _35945_/Q _21170_/X _21307_/X VGND VGND VPWR
+ VPWR _21348_/X sky130_fd_sc_hd__mux4_1
XFILLER_108_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29993_ _29993_/A VGND VGND VPWR VPWR _35250_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28944_ _28944_/A VGND VGND VPWR VPWR _34783_/D sky130_fd_sc_hd__clkbuf_1
X_24067_ _24067_/A VGND VGND VPWR VPWR _32574_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21279_ _32103_/Q _32295_/Q _32359_/Q _35879_/Q _21174_/X _20962_/X VGND VGND VPWR
+ VPWR _21279_/X sky130_fd_sc_hd__mux4_1
XFILLER_151_879 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23018_ input37/X VGND VGND VPWR VPWR _23018_/X sky130_fd_sc_hd__buf_2
XFILLER_110_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28875_ _28875_/A VGND VGND VPWR VPWR _34750_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_131_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27826_ _27825_/X _34257_/Q _27826_/S VGND VGND VPWR VPWR _27827_/A sky130_fd_sc_hd__mux2_1
XTAP_4210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27757_ input31/X VGND VGND VPWR VPWR _27757_/X sky130_fd_sc_hd__clkbuf_4
X_24969_ _24969_/A VGND VGND VPWR VPWR _32972_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17510_ _17506_/X _17507_/X _17508_/X _17509_/X VGND VGND VPWR VPWR _17510_/X sky130_fd_sc_hd__a22o_1
XTAP_4287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26708_ _26708_/A VGND VGND VPWR VPWR _33787_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_217_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18490_ _18330_/X _18488_/X _18489_/X _18341_/X VGND VGND VPWR VPWR _18490_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27688_ _27688_/A VGND VGND VPWR VPWR _34212_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_874 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29427_ _34997_/Q _29426_/X _29451_/S VGND VGND VPWR VPWR _29428_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17441_ _17158_/X _17439_/X _17440_/X _17163_/X VGND VGND VPWR VPWR _17441_/X sky130_fd_sc_hd__a22o_1
XFILLER_221_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26639_ _26639_/A VGND VGND VPWR VPWR _33754_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29358_ _34975_/Q _29357_/X _29358_/S VGND VGND VPWR VPWR _29359_/A sky130_fd_sc_hd__mux2_1
X_17372_ _17372_/A VGND VGND VPWR VPWR _31994_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19111_ _19105_/X _19106_/X _19109_/X _19110_/X VGND VGND VPWR VPWR _19111_/X sky130_fd_sc_hd__a22o_1
X_16323_ _32605_/Q _32541_/Q _32477_/Q _35933_/Q _16217_/X _17717_/A VGND VGND VPWR
+ VPWR _16323_/X sky130_fd_sc_hd__mux4_1
X_28309_ _28378_/S VGND VGND VPWR VPWR _28328_/S sky130_fd_sc_hd__buf_4
X_29289_ _34947_/Q _27174_/X _29297_/S VGND VGND VPWR VPWR _29290_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19042_ _34153_/Q _34089_/Q _34025_/Q _33961_/Q _19040_/X _19041_/X VGND VGND VPWR
+ VPWR _19042_/X sky130_fd_sc_hd__mux4_1
X_31320_ _27695_/X _35879_/Q _31324_/S VGND VGND VPWR VPWR _31321_/A sky130_fd_sc_hd__mux2_1
X_16254_ _32091_/Q _32283_/Q _32347_/Q _35867_/Q _16221_/X _17867_/A VGND VGND VPWR
+ VPWR _16254_/X sky130_fd_sc_hd__mux4_1
XFILLER_9_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31251_ _31251_/A VGND VGND VPWR VPWR _35846_/D sky130_fd_sc_hd__clkbuf_1
X_16185_ _32601_/Q _32537_/Q _32473_/Q _35929_/Q _17866_/A _17717_/A VGND VGND VPWR
+ VPWR _16185_/X sky130_fd_sc_hd__mux4_1
Xoutput207 _36240_/Q VGND VGND VPWR VPWR D2[58] sky130_fd_sc_hd__buf_2
X_30202_ _30202_/A _30877_/A VGND VGND VPWR VPWR _30335_/S sky130_fd_sc_hd__nor2_8
Xoutput218 _32406_/Q VGND VGND VPWR VPWR D3[0] sky130_fd_sc_hd__buf_2
Xoutput229 _32407_/Q VGND VGND VPWR VPWR D3[1] sky130_fd_sc_hd__buf_2
X_31182_ _31182_/A VGND VGND VPWR VPWR _35813_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_1247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30133_ _30133_/A VGND VGND VPWR VPWR _35316_/D sky130_fd_sc_hd__clkbuf_1
X_19944_ _19940_/X _19943_/X _19804_/X VGND VGND VPWR VPWR _19954_/C sky130_fd_sc_hd__o21ba_1
XFILLER_99_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35990_ _35990_/CLK _35990_/D VGND VGND VPWR VPWR _35990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30064_ _30064_/A VGND VGND VPWR VPWR _35284_/D sky130_fd_sc_hd__clkbuf_1
X_34941_ _34941_/CLK _34941_/D VGND VGND VPWR VPWR _34941_/Q sky130_fd_sc_hd__dfxtp_1
X_19875_ _35456_/Q _35392_/Q _35328_/Q _35264_/Q _19554_/X _19555_/X VGND VGND VPWR
+ VPWR _19875_/X sky130_fd_sc_hd__mux4_1
XFILLER_214_1247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18826_ _34914_/Q _34850_/Q _34786_/Q _34722_/Q _18754_/X _18755_/X VGND VGND VPWR
+ VPWR _18826_/X sky130_fd_sc_hd__mux4_1
XTAP_6190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34872_ _35833_/CLK _34872_/D VGND VGND VPWR VPWR _34872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33823_ _36129_/CLK _33823_/D VGND VGND VPWR VPWR _33823_/Q sky130_fd_sc_hd__dfxtp_1
X_18757_ _19463_/A VGND VGND VPWR VPWR _18757_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_82_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17708_ _17704_/X _17705_/X _17706_/X _17707_/X VGND VGND VPWR VPWR _17708_/X sky130_fd_sc_hd__a22o_1
XFILLER_224_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33754_ _33818_/CLK _33754_/D VGND VGND VPWR VPWR _33754_/Q sky130_fd_sc_hd__dfxtp_1
X_30966_ _30966_/A VGND VGND VPWR VPWR _35711_/D sky130_fd_sc_hd__clkbuf_1
X_18688_ _20261_/A VGND VGND VPWR VPWR _18688_/X sky130_fd_sc_hd__buf_4
XFILLER_97_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32705_ _35902_/CLK _32705_/D VGND VGND VPWR VPWR _32705_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17639_ _35650_/Q _35010_/Q _34370_/Q _33730_/Q _17497_/X _17498_/X VGND VGND VPWR
+ VPWR _17639_/X sky130_fd_sc_hd__mux4_1
XFILLER_58_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33685_ _33685_/CLK _33685_/D VGND VGND VPWR VPWR _33685_/Q sky130_fd_sc_hd__dfxtp_1
X_30897_ _35679_/Q input64/X _30897_/S VGND VGND VPWR VPWR _30898_/A sky130_fd_sc_hd__mux2_1
XFILLER_224_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20650_ _22400_/A VGND VGND VPWR VPWR _20650_/X sky130_fd_sc_hd__buf_6
X_32636_ _35965_/CLK _32636_/D VGND VGND VPWR VPWR _32636_/Q sky130_fd_sc_hd__dfxtp_1
X_35424_ _36005_/CLK _35424_/D VGND VGND VPWR VPWR _35424_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19309_ _34672_/Q _34608_/Q _34544_/Q _34480_/Q _19239_/X _19240_/X VGND VGND VPWR
+ VPWR _19309_/X sky130_fd_sc_hd__mux4_1
X_35355_ _36059_/CLK _35355_/D VGND VGND VPWR VPWR _35355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20581_ _22459_/A VGND VGND VPWR VPWR _20581_/X sky130_fd_sc_hd__clkbuf_4
X_32567_ _35961_/CLK _32567_/D VGND VGND VPWR VPWR _32567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22320_ _34436_/Q _36164_/Q _34308_/Q _34244_/Q _22182_/X _22183_/X VGND VGND VPWR
+ VPWR _22320_/X sky130_fd_sc_hd__mux4_1
XFILLER_176_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34306_ _36163_/CLK _34306_/D VGND VGND VPWR VPWR _34306_/Q sky130_fd_sc_hd__dfxtp_1
X_31518_ _27788_/X _35973_/Q _31522_/S VGND VGND VPWR VPWR _31519_/A sky130_fd_sc_hd__mux2_1
X_35286_ _36118_/CLK _35286_/D VGND VGND VPWR VPWR _35286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32498_ _35955_/CLK _32498_/D VGND VGND VPWR VPWR _32498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22251_ _34946_/Q _34882_/Q _34818_/Q _34754_/Q _22113_/X _22114_/X VGND VGND VPWR
+ VPWR _22251_/X sky130_fd_sc_hd__mux4_1
XFILLER_192_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34237_ _36157_/CLK _34237_/D VGND VGND VPWR VPWR _34237_/Q sky130_fd_sc_hd__dfxtp_1
X_31449_ _27686_/X _35940_/Q _31459_/S VGND VGND VPWR VPWR _31450_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21202_ _21100_/X _21200_/X _21201_/X _21103_/X VGND VGND VPWR VPWR _21202_/X sky130_fd_sc_hd__a22o_1
XFILLER_155_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22182_ _22535_/A VGND VGND VPWR VPWR _22182_/X sky130_fd_sc_hd__buf_6
XFILLER_173_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34168_ _35320_/CLK _34168_/D VGND VGND VPWR VPWR _34168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33119_ _33119_/CLK _33119_/D VGND VGND VPWR VPWR _33119_/Q sky130_fd_sc_hd__dfxtp_1
X_21133_ _21093_/X _21131_/X _21132_/X _21098_/X VGND VGND VPWR VPWR _21133_/X sky130_fd_sc_hd__a22o_1
X_26990_ _33921_/Q _23432_/X _27002_/S VGND VGND VPWR VPWR _26991_/A sky130_fd_sc_hd__mux2_1
X_34099_ _34099_/CLK _34099_/D VGND VGND VPWR VPWR _34099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25941_ _24988_/X _33427_/Q _25945_/S VGND VGND VPWR VPWR _25942_/A sky130_fd_sc_hd__mux2_1
X_21064_ _34145_/Q _34081_/Q _34017_/Q _33953_/Q _20987_/X _20988_/X VGND VGND VPWR
+ VPWR _21064_/X sky130_fd_sc_hd__mux4_1
XFILLER_87_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20015_ _34692_/Q _34628_/Q _34564_/Q _34500_/Q _19945_/X _19946_/X VGND VGND VPWR
+ VPWR _20015_/X sky130_fd_sc_hd__mux4_1
X_28660_ _28660_/A VGND VGND VPWR VPWR _34649_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_246_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25872_ _24886_/X _33394_/Q _25874_/S VGND VGND VPWR VPWR _25873_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27611_ _34184_/Q _27189_/X _27629_/S VGND VGND VPWR VPWR _27612_/A sky130_fd_sc_hd__mux2_1
X_24823_ _24823_/A VGND VGND VPWR VPWR _32925_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28591_ _28591_/A VGND VGND VPWR VPWR _34617_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27542_ _27542_/A VGND VGND VPWR VPWR _34151_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24754_ _24754_/A VGND VGND VPWR VPWR _32897_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21966_ _21753_/X _21962_/X _21965_/X _21756_/X VGND VGND VPWR VPWR _21966_/X sky130_fd_sc_hd__a22o_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23705_ _27232_/B _25132_/A VGND VGND VPWR VPWR _28786_/B sky130_fd_sc_hd__nand2_4
XFILLER_15_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27473_ _34119_/Q _27186_/X _27473_/S VGND VGND VPWR VPWR _27474_/A sky130_fd_sc_hd__mux2_1
X_20917_ _33373_/Q _33309_/Q _33245_/Q _33181_/Q _20602_/X _20603_/X VGND VGND VPWR
+ VPWR _20917_/X sky130_fd_sc_hd__mux4_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24685_ _24685_/A VGND VGND VPWR VPWR _32864_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21897_ _34424_/Q _36152_/Q _34296_/Q _34232_/Q _21829_/X _21830_/X VGND VGND VPWR
+ VPWR _21897_/X sky130_fd_sc_hd__mux4_1
XFILLER_214_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29212_ _29212_/A VGND VGND VPWR VPWR _34910_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26424_ _33655_/Q _23399_/X _26436_/S VGND VGND VPWR VPWR _26425_/A sky130_fd_sc_hd__mux2_1
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20848_ _33883_/Q _33819_/Q _33755_/Q _36059_/Q _20712_/X _20713_/X VGND VGND VPWR
+ VPWR _20848_/X sky130_fd_sc_hd__mux4_1
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23636_ _22984_/X _32309_/Q _23652_/S VGND VGND VPWR VPWR _23637_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29143_ _29191_/S VGND VGND VPWR VPWR _29162_/S sky130_fd_sc_hd__buf_4
XFILLER_161_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26355_ _33622_/Q _23225_/X _26373_/S VGND VGND VPWR VPWR _26356_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_1146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20779_ _34137_/Q _34073_/Q _34009_/Q _33945_/Q _20609_/X _20611_/X VGND VGND VPWR
+ VPWR _20779_/X sky130_fd_sc_hd__mux4_1
X_23567_ _25132_/A input83/X input89/X _27232_/B VGND VGND VPWR VPWR _23568_/A sky130_fd_sc_hd__and4b_1
XFILLER_168_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25306_ _25306_/A VGND VGND VPWR VPWR _33126_/D sky130_fd_sc_hd__clkbuf_1
X_29074_ _34845_/Q _27056_/X _29078_/S VGND VGND VPWR VPWR _29075_/A sky130_fd_sc_hd__mux2_1
X_22518_ _32650_/Q _32586_/Q _32522_/Q _35978_/Q _22229_/X _22366_/X VGND VGND VPWR
+ VPWR _22518_/X sky130_fd_sc_hd__mux4_1
XFILLER_127_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23498_ input60/X VGND VGND VPWR VPWR _23498_/X sky130_fd_sc_hd__clkbuf_4
X_26286_ _24899_/X _33590_/Q _26300_/S VGND VGND VPWR VPWR _26287_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28025_ _34349_/Q _27106_/X _28037_/S VGND VGND VPWR VPWR _28026_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22449_ _35720_/Q _32230_/Q _35592_/Q _35528_/Q _22270_/X _22271_/X VGND VGND VPWR
+ VPWR _22449_/X sky130_fd_sc_hd__mux4_1
X_25237_ _25237_/A VGND VGND VPWR VPWR _33094_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25168_ _25168_/A VGND VGND VPWR VPWR _33061_/D sky130_fd_sc_hd__clkbuf_1
X_24119_ _24251_/S VGND VGND VPWR VPWR _24138_/S sky130_fd_sc_hd__buf_6
X_25099_ _24948_/X _33030_/Q _25101_/S VGND VGND VPWR VPWR _25100_/A sky130_fd_sc_hd__mux2_1
X_17990_ _17985_/X _17989_/X _17846_/X _17847_/X VGND VGND VPWR VPWR _18007_/B sky130_fd_sc_hd__o211a_1
X_29976_ _35242_/Q _29391_/X _29994_/S VGND VGND VPWR VPWR _29977_/A sky130_fd_sc_hd__mux2_1
X_28927_ _34775_/Q _27038_/X _28943_/S VGND VGND VPWR VPWR _28928_/A sky130_fd_sc_hd__mux2_1
X_16941_ _34670_/Q _34606_/Q _34542_/Q _34478_/Q _16939_/X _16940_/X VGND VGND VPWR
+ VPWR _16941_/X sky130_fd_sc_hd__mux4_1
XFILLER_172_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19660_ _19656_/X _19657_/X _19658_/X _19659_/X VGND VGND VPWR VPWR _19660_/X sky130_fd_sc_hd__a22o_1
XFILLER_237_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16872_ _16868_/X _16871_/X _16798_/X VGND VGND VPWR VPWR _16882_/C sky130_fd_sc_hd__o21ba_1
X_28858_ _28858_/A VGND VGND VPWR VPWR _34742_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18611_ _18607_/X _18610_/X _18404_/X VGND VGND VPWR VPWR _18612_/D sky130_fd_sc_hd__o21ba_1
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27809_ _27809_/A VGND VGND VPWR VPWR _34251_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19591_ _19587_/X _19590_/X _19451_/X VGND VGND VPWR VPWR _19601_/C sky130_fd_sc_hd__o21ba_1
XFILLER_93_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28789_ _28921_/S VGND VGND VPWR VPWR _28808_/S sky130_fd_sc_hd__buf_4
XFILLER_225_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_994 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18542_ _18542_/A _18542_/B _18542_/C _18542_/D VGND VGND VPWR VPWR _18543_/A sky130_fd_sc_hd__or4_1
XTAP_4084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30820_ _30820_/A VGND VGND VPWR VPWR _35642_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_234_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18473_ _34904_/Q _34840_/Q _34776_/Q _34712_/Q _18396_/X _18398_/X VGND VGND VPWR
+ VPWR _18473_/X sky130_fd_sc_hd__mux4_1
X_30751_ _30751_/A VGND VGND VPWR VPWR _35609_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1027 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17424_ _17915_/A VGND VGND VPWR VPWR _17424_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33470_ _35453_/CLK _33470_/D VGND VGND VPWR VPWR _33470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30682_ _35577_/Q _29438_/X _30690_/S VGND VGND VPWR VPWR _30683_/A sky130_fd_sc_hd__mux2_1
XFILLER_92_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32421_ _33828_/CLK _32421_/D VGND VGND VPWR VPWR _32421_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17355_ _17351_/X _17352_/X _17353_/X _17354_/X VGND VGND VPWR VPWR _17355_/X sky130_fd_sc_hd__a22o_1
XFILLER_140_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16306_ _35164_/Q _35100_/Q _35036_/Q _32156_/Q _16304_/X _16305_/X VGND VGND VPWR
+ VPWR _16306_/X sky130_fd_sc_hd__mux4_1
X_35140_ _35717_/CLK _35140_/D VGND VGND VPWR VPWR _35140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32352_ _32804_/CLK _32352_/D VGND VGND VPWR VPWR _32352_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17286_ _35640_/Q _35000_/Q _34360_/Q _33720_/Q _17144_/X _17145_/X VGND VGND VPWR
+ VPWR _17286_/X sky130_fd_sc_hd__mux4_1
XFILLER_201_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31303_ _27670_/X _35871_/Q _31303_/S VGND VGND VPWR VPWR _31304_/A sky130_fd_sc_hd__mux2_1
X_19025_ _20235_/A VGND VGND VPWR VPWR _19025_/X sky130_fd_sc_hd__buf_6
X_16237_ _16078_/X _16235_/X _16236_/X _16088_/X VGND VGND VPWR VPWR _16237_/X sky130_fd_sc_hd__a22o_1
X_35071_ _35071_/CLK _35071_/D VGND VGND VPWR VPWR _35071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32283_ _35860_/CLK _32283_/D VGND VGND VPWR VPWR _32283_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34022_ _34790_/CLK _34022_/D VGND VGND VPWR VPWR _34022_/Q sky130_fd_sc_hd__dfxtp_1
X_31234_ _27766_/X _35838_/Q _31252_/S VGND VGND VPWR VPWR _31235_/A sky130_fd_sc_hd__mux2_1
X_16168_ _35160_/Q _35096_/Q _35032_/Q _32152_/Q _16083_/X _16085_/X VGND VGND VPWR
+ VPWR _16168_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31165_ _31165_/A VGND VGND VPWR VPWR _35805_/D sky130_fd_sc_hd__clkbuf_1
X_16099_ _34902_/Q _34838_/Q _34774_/Q _34710_/Q _16096_/X _16098_/X VGND VGND VPWR
+ VPWR _16099_/X sky130_fd_sc_hd__mux4_1
XFILLER_138_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30116_ _30116_/A VGND VGND VPWR VPWR _35308_/D sky130_fd_sc_hd__clkbuf_1
X_19927_ _19859_/X _19925_/X _19926_/X _19862_/X VGND VGND VPWR VPWR _19927_/X sky130_fd_sc_hd__a22o_1
XFILLER_190_1350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35973_ _35973_/CLK _35973_/D VGND VGND VPWR VPWR _35973_/Q sky130_fd_sc_hd__dfxtp_1
X_31096_ _31096_/A VGND VGND VPWR VPWR _35773_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_229_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30047_ _35276_/Q _29497_/X _30057_/S VGND VGND VPWR VPWR _30048_/A sky130_fd_sc_hd__mux2_1
X_34924_ _34924_/CLK _34924_/D VGND VGND VPWR VPWR _34924_/Q sky130_fd_sc_hd__dfxtp_1
X_19858_ _19852_/X _19855_/X _19856_/X _19857_/X VGND VGND VPWR VPWR _19858_/X sky130_fd_sc_hd__a22o_1
XFILLER_151_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18809_ _32098_/Q _32290_/Q _32354_/Q _35874_/Q _18521_/X _18662_/X VGND VGND VPWR
+ VPWR _18809_/X sky130_fd_sc_hd__mux4_1
XFILLER_216_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34855_ _34921_/CLK _34855_/D VGND VGND VPWR VPWR _34855_/Q sky130_fd_sc_hd__dfxtp_1
X_19789_ _19712_/X _19787_/X _19788_/X _19718_/X VGND VGND VPWR VPWR _19789_/X sky130_fd_sc_hd__a22o_1
XFILLER_186_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33806_ _33934_/CLK _33806_/D VGND VGND VPWR VPWR _33806_/Q sky130_fd_sc_hd__dfxtp_1
X_21820_ _35638_/Q _34998_/Q _34358_/Q _33718_/Q _21744_/X _21745_/X VGND VGND VPWR
+ VPWR _21820_/X sky130_fd_sc_hd__mux4_1
XFILLER_110_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31998_ _36207_/CLK _31998_/D VGND VGND VPWR VPWR _31998_/Q sky130_fd_sc_hd__dfxtp_1
X_34786_ _34914_/CLK _34786_/D VGND VGND VPWR VPWR _34786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21751_ _22457_/A VGND VGND VPWR VPWR _21751_/X sky130_fd_sc_hd__buf_4
X_33737_ _35658_/CLK _33737_/D VGND VGND VPWR VPWR _33737_/Q sky130_fd_sc_hd__dfxtp_1
X_30949_ _30949_/A VGND VGND VPWR VPWR _35703_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20702_ _20691_/X _20695_/X _20699_/X _20701_/X VGND VGND VPWR VPWR _20702_/X sky130_fd_sc_hd__a22o_1
XFILLER_51_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21682_ _21676_/X _21681_/X _21398_/X VGND VGND VPWR VPWR _21690_/C sky130_fd_sc_hd__o21ba_1
X_24470_ _23002_/X _32763_/Q _24474_/S VGND VGND VPWR VPWR _24471_/A sky130_fd_sc_hd__mux2_1
X_33668_ _34182_/CLK _33668_/D VGND VGND VPWR VPWR _33668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35407_ _35471_/CLK _35407_/D VGND VGND VPWR VPWR _35407_/Q sky130_fd_sc_hd__dfxtp_1
X_20633_ _20663_/A VGND VGND VPWR VPWR _22374_/A sky130_fd_sc_hd__clkbuf_16
X_23421_ _23499_/S VGND VGND VPWR VPWR _23451_/S sky130_fd_sc_hd__buf_6
X_32619_ _36010_/CLK _32619_/D VGND VGND VPWR VPWR _32619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33599_ _34174_/CLK _33599_/D VGND VGND VPWR VPWR _33599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26140_ _24883_/X _33521_/Q _26144_/S VGND VGND VPWR VPWR _26141_/A sky130_fd_sc_hd__mux2_1
X_23352_ _23352_/A VGND VGND VPWR VPWR _32192_/D sky130_fd_sc_hd__clkbuf_1
X_20564_ _35669_/Q _35029_/Q _34389_/Q _33749_/Q _18412_/X _18413_/X VGND VGND VPWR
+ VPWR _20564_/X sky130_fd_sc_hd__mux4_1
X_35338_ _35849_/CLK _35338_/D VGND VGND VPWR VPWR _35338_/Q sky130_fd_sc_hd__dfxtp_1
X_22303_ _22297_/X _22302_/X _22093_/X _22094_/X VGND VGND VPWR VPWR _22324_/B sky130_fd_sc_hd__o211a_1
X_26071_ _26071_/A VGND VGND VPWR VPWR _33488_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23283_ input9/X VGND VGND VPWR VPWR _23283_/X sky130_fd_sc_hd__buf_4
X_20495_ _20491_/X _20494_/X _20138_/A VGND VGND VPWR VPWR _20517_/A sky130_fd_sc_hd__o21ba_1
X_35269_ _35845_/CLK _35269_/D VGND VGND VPWR VPWR _35269_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_5_23_0_CLK clkbuf_2_2_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_23_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_180_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22234_ _32130_/Q _32322_/Q _32386_/Q _35906_/Q _22233_/X _22021_/X VGND VGND VPWR
+ VPWR _22234_/X sky130_fd_sc_hd__mux4_1
X_25022_ _24834_/X _32993_/Q _25038_/S VGND VGND VPWR VPWR _25023_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_1193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29830_ _35173_/Q _29376_/X _29838_/S VGND VGND VPWR VPWR _29831_/A sky130_fd_sc_hd__mux2_1
X_22165_ _32640_/Q _32576_/Q _32512_/Q _35968_/Q _21876_/X _22013_/X VGND VGND VPWR
+ VPWR _22165_/X sky130_fd_sc_hd__mux4_1
XTAP_6904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21116_ _35426_/Q _35362_/Q _35298_/Q _35234_/Q _20795_/X _20796_/X VGND VGND VPWR
+ VPWR _21116_/X sky130_fd_sc_hd__mux4_1
XTAP_6937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29761_ _29761_/A VGND VGND VPWR VPWR _35140_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22096_ _35710_/Q _32219_/Q _35582_/Q _35518_/Q _21917_/X _21918_/X VGND VGND VPWR
+ VPWR _22096_/X sky130_fd_sc_hd__mux4_1
XFILLER_132_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26973_ _33913_/Q _23405_/X _26981_/S VGND VGND VPWR VPWR _26974_/A sky130_fd_sc_hd__mux2_1
XTAP_6959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28712_ _28712_/A VGND VGND VPWR VPWR _34674_/D sky130_fd_sc_hd__clkbuf_1
X_25924_ _25924_/A VGND VGND VPWR VPWR _33418_/D sky130_fd_sc_hd__clkbuf_1
X_21047_ _21753_/A VGND VGND VPWR VPWR _21047_/X sky130_fd_sc_hd__buf_4
X_29692_ _29692_/A VGND VGND VPWR VPWR _35107_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28643_ _28643_/A VGND VGND VPWR VPWR _34642_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25855_ _25945_/S VGND VGND VPWR VPWR _25874_/S sky130_fd_sc_hd__buf_4
XFILLER_247_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_1043 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24806_ input23/X VGND VGND VPWR VPWR _24806_/X sky130_fd_sc_hd__clkbuf_4
X_28574_ _28574_/A VGND VGND VPWR VPWR _34609_/D sky130_fd_sc_hd__clkbuf_1
X_25786_ _24958_/X _33353_/Q _25802_/S VGND VGND VPWR VPWR _25787_/A sky130_fd_sc_hd__mux2_1
XFILLER_216_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22998_ _22998_/A VGND VGND VPWR VPWR _32057_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_885 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27525_ _27525_/A VGND VGND VPWR VPWR _34143_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24737_ _24737_/A VGND VGND VPWR VPWR _32889_/D sky130_fd_sc_hd__clkbuf_1
X_21949_ _21667_/X _21945_/X _21948_/X _21671_/X VGND VGND VPWR VPWR _21949_/X sky130_fd_sc_hd__a22o_1
XFILLER_199_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27456_ _27456_/A VGND VGND VPWR VPWR _34110_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24668_ _24668_/A VGND VGND VPWR VPWR _32856_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26407_ _33647_/Q _23316_/X _26415_/S VGND VGND VPWR VPWR _26408_/A sky130_fd_sc_hd__mux2_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23619_ _22959_/X _32301_/Q _23631_/S VGND VGND VPWR VPWR _23620_/A sky130_fd_sc_hd__mux2_1
X_27387_ _34078_/Q _27059_/X _27389_/S VGND VGND VPWR VPWR _27388_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24599_ _22993_/X _32824_/Q _24609_/S VGND VGND VPWR VPWR _24600_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29126_ _29126_/A VGND VGND VPWR VPWR _34869_/D sky130_fd_sc_hd__clkbuf_1
X_17140_ _17846_/A VGND VGND VPWR VPWR _17140_/X sky130_fd_sc_hd__clkbuf_4
X_26338_ _24976_/X _33615_/Q _26342_/S VGND VGND VPWR VPWR _26339_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29057_ _29057_/A VGND VGND VPWR VPWR _34837_/D sky130_fd_sc_hd__clkbuf_1
X_17071_ _17915_/A VGND VGND VPWR VPWR _17071_/X sky130_fd_sc_hd__clkbuf_4
X_26269_ _24874_/X _33582_/Q _26279_/S VGND VGND VPWR VPWR _26270_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16022_ _17766_/A VGND VGND VPWR VPWR _17717_/A sky130_fd_sc_hd__buf_8
X_28008_ _34341_/Q _27081_/X _28016_/S VGND VGND VPWR VPWR _28009_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17973_ _17973_/A _17973_/B _17973_/C _17973_/D VGND VGND VPWR VPWR _17974_/A sky130_fd_sc_hd__or4_2
XFILLER_123_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29959_ _35234_/Q _29367_/X _29973_/S VGND VGND VPWR VPWR _29960_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16924_ _32622_/Q _32558_/Q _32494_/Q _35950_/Q _16923_/X _16707_/X VGND VGND VPWR
+ VPWR _16924_/X sky130_fd_sc_hd__mux4_1
X_19712_ _20205_/A VGND VGND VPWR VPWR _19712_/X sky130_fd_sc_hd__clkbuf_4
X_32970_ _36042_/CLK _32970_/D VGND VGND VPWR VPWR _32970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_242_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31921_ _23441_/X _36164_/Q _31927_/S VGND VGND VPWR VPWR _31922_/A sky130_fd_sc_hd__mux2_1
X_16855_ _33900_/Q _33836_/Q _33772_/Q _36076_/Q _16671_/X _16672_/X VGND VGND VPWR
+ VPWR _16855_/X sky130_fd_sc_hd__mux4_1
X_19643_ _33146_/Q _36026_/Q _33018_/Q _32954_/Q _19362_/X _19363_/X VGND VGND VPWR
+ VPWR _19643_/X sky130_fd_sc_hd__mux4_1
XFILLER_238_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34640_ _35217_/CLK _34640_/D VGND VGND VPWR VPWR _34640_/Q sky130_fd_sc_hd__dfxtp_1
X_19574_ _19506_/X _19572_/X _19573_/X _19509_/X VGND VGND VPWR VPWR _19574_/X sky130_fd_sc_hd__a22o_1
X_31852_ _23271_/X _36131_/Q _31864_/S VGND VGND VPWR VPWR _31853_/A sky130_fd_sc_hd__mux2_1
X_16786_ _16714_/X _16784_/X _16785_/X _16718_/X VGND VGND VPWR VPWR _16786_/X sky130_fd_sc_hd__a22o_1
XFILLER_225_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18525_ _18520_/X _18524_/X _18344_/X _18346_/X VGND VGND VPWR VPWR _18542_/B sky130_fd_sc_hd__o211a_1
X_30803_ _30803_/A VGND VGND VPWR VPWR _35634_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34571_ _35208_/CLK _34571_/D VGND VGND VPWR VPWR _34571_/Q sky130_fd_sc_hd__dfxtp_1
X_31783_ _31783_/A VGND VGND VPWR VPWR _36098_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18456_ _32088_/Q _32280_/Q _32344_/Q _35864_/Q _18332_/X _20167_/A VGND VGND VPWR
+ VPWR _18456_/X sky130_fd_sc_hd__mux4_1
X_30734_ _35602_/Q _29515_/X _30740_/S VGND VGND VPWR VPWR _30735_/A sky130_fd_sc_hd__mux2_1
X_33522_ _34098_/CLK _33522_/D VGND VGND VPWR VPWR _33522_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17407_ _17199_/X _17405_/X _17406_/X _17204_/X VGND VGND VPWR VPWR _17407_/X sky130_fd_sc_hd__a22o_1
XFILLER_60_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36241_ _36242_/CLK _36241_/D VGND VGND VPWR VPWR _36241_/Q sky130_fd_sc_hd__dfxtp_1
X_33453_ _36077_/CLK _33453_/D VGND VGND VPWR VPWR _33453_/Q sky130_fd_sc_hd__dfxtp_1
X_18387_ _20071_/A VGND VGND VPWR VPWR _19456_/A sky130_fd_sc_hd__clkbuf_16
X_30665_ _35569_/Q _29413_/X _30669_/S VGND VGND VPWR VPWR _30666_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32404_ _35989_/CLK _32404_/D VGND VGND VPWR VPWR _32404_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17338_ _33402_/Q _33338_/Q _33274_/Q _33210_/Q _17127_/X _17128_/X VGND VGND VPWR
+ VPWR _17338_/X sky130_fd_sc_hd__mux4_1
XFILLER_53_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36172_ _36173_/CLK _36172_/D VGND VGND VPWR VPWR _36172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33384_ _36072_/CLK _33384_/D VGND VGND VPWR VPWR _33384_/Q sky130_fd_sc_hd__dfxtp_1
X_30596_ _30596_/A VGND VGND VPWR VPWR _35536_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32335_ _32879_/CLK _32335_/D VGND VGND VPWR VPWR _32335_/Q sky130_fd_sc_hd__dfxtp_1
X_35123_ _35187_/CLK _35123_/D VGND VGND VPWR VPWR _35123_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17269_ _33656_/Q _33592_/Q _33528_/Q _33464_/Q _17200_/X _17201_/X VGND VGND VPWR
+ VPWR _17269_/X sky130_fd_sc_hd__mux4_1
XFILLER_220_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19008_ _32616_/Q _32552_/Q _32488_/Q _35944_/Q _18870_/X _19007_/X VGND VGND VPWR
+ VPWR _19008_/X sky130_fd_sc_hd__mux4_1
XFILLER_146_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35054_ _35183_/CLK _35054_/D VGND VGND VPWR VPWR _35054_/Q sky130_fd_sc_hd__dfxtp_1
X_20280_ _20212_/X _20278_/X _20279_/X _20215_/X VGND VGND VPWR VPWR _20280_/X sky130_fd_sc_hd__a22o_1
X_32266_ _35212_/CLK _32266_/D VGND VGND VPWR VPWR _32266_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34005_ _34773_/CLK _34005_/D VGND VGND VPWR VPWR _34005_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31217_ _27742_/X _35830_/Q _31231_/S VGND VGND VPWR VPWR _31218_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32197_ _35690_/CLK _32197_/D VGND VGND VPWR VPWR _32197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31148_ _31148_/A VGND VGND VPWR VPWR _31281_/S sky130_fd_sc_hd__buf_8
XFILLER_115_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23970_ _23970_/A VGND VGND VPWR VPWR _32529_/D sky130_fd_sc_hd__clkbuf_1
X_31079_ _35765_/Q input25/X _31095_/S VGND VGND VPWR VPWR _31080_/A sky130_fd_sc_hd__mux2_1
X_35956_ _35956_/CLK _35956_/D VGND VGND VPWR VPWR _35956_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34907_ _34907_/CLK _34907_/D VGND VGND VPWR VPWR _34907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_217_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22921_ _22921_/A VGND VGND VPWR VPWR _32032_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_217_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1069 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35887_ _35951_/CLK _35887_/D VGND VGND VPWR VPWR _35887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25640_ _24942_/X _33284_/Q _25646_/S VGND VGND VPWR VPWR _25641_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34838_ _34904_/CLK _34838_/D VGND VGND VPWR VPWR _34838_/Q sky130_fd_sc_hd__dfxtp_1
X_22852_ _33429_/Q _33365_/Q _33301_/Q _33237_/Q _20637_/X _20639_/X VGND VGND VPWR
+ VPWR _22852_/X sky130_fd_sc_hd__mux4_1
XFILLER_244_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21803_ _34166_/Q _34102_/Q _34038_/Q _33974_/Q _21693_/X _21694_/X VGND VGND VPWR
+ VPWR _21803_/X sky130_fd_sc_hd__mux4_1
X_25571_ _24840_/X _33251_/Q _25583_/S VGND VGND VPWR VPWR _25572_/A sky130_fd_sc_hd__mux2_1
X_34769_ _34897_/CLK _34769_/D VGND VGND VPWR VPWR _34769_/Q sky130_fd_sc_hd__dfxtp_1
X_22783_ _34450_/Q _36178_/Q _34322_/Q _34258_/Q _22535_/X _22536_/X VGND VGND VPWR
+ VPWR _22783_/X sky130_fd_sc_hd__mux4_1
X_27310_ _27310_/A VGND VGND VPWR VPWR _34041_/D sky130_fd_sc_hd__clkbuf_1
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24522_ _23079_/X _32788_/Q _24524_/S VGND VGND VPWR VPWR _24523_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_22 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28290_ _28290_/A VGND VGND VPWR VPWR _34474_/D sky130_fd_sc_hd__clkbuf_1
X_21734_ _32628_/Q _32564_/Q _32500_/Q _35956_/Q _21523_/X _21660_/X VGND VGND VPWR
+ VPWR _21734_/X sky130_fd_sc_hd__mux4_1
XFILLER_169_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27241_ _27241_/A VGND VGND VPWR VPWR _34008_/D sky130_fd_sc_hd__clkbuf_1
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24453_ _22977_/X _32755_/Q _24453_/S VGND VGND VPWR VPWR _24454_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21665_ _22510_/A VGND VGND VPWR VPWR _21665_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_240_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23404_ _23404_/A VGND VGND VPWR VPWR _32213_/D sky130_fd_sc_hd__clkbuf_1
X_27172_ _33986_/Q _27171_/X _27187_/S VGND VGND VPWR VPWR _27173_/A sky130_fd_sc_hd__mux2_1
X_20616_ _20597_/X _20613_/X _20615_/X VGND VGND VPWR VPWR _20706_/A sky130_fd_sc_hd__o21ba_1
X_24384_ _24384_/A VGND VGND VPWR VPWR _32722_/D sky130_fd_sc_hd__clkbuf_1
X_21596_ _21314_/X _21592_/X _21595_/X _21318_/X VGND VGND VPWR VPWR _21596_/X sky130_fd_sc_hd__a22o_1
XFILLER_193_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26123_ _24858_/X _33513_/Q _26123_/S VGND VGND VPWR VPWR _26124_/A sky130_fd_sc_hd__mux2_1
X_20547_ _20547_/A _20547_/B _20547_/C _20547_/D VGND VGND VPWR VPWR _20548_/A sky130_fd_sc_hd__or4_1
X_23335_ _32185_/Q _23258_/X _23335_/S VGND VGND VPWR VPWR _23336_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_874 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26054_ _24954_/X _33480_/Q _26072_/S VGND VGND VPWR VPWR _26055_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20478_ _18301_/X _20476_/X _20477_/X _18307_/X VGND VGND VPWR VPWR _20478_/X sky130_fd_sc_hd__a22o_1
X_23266_ _32161_/Q _23265_/X _23290_/S VGND VGND VPWR VPWR _23267_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25005_ _24809_/X _32985_/Q _25017_/S VGND VGND VPWR VPWR _25006_/A sky130_fd_sc_hd__mux2_1
X_22217_ _34945_/Q _34881_/Q _34817_/Q _34753_/Q _22113_/X _22114_/X VGND VGND VPWR
+ VPWR _22217_/X sky130_fd_sc_hd__mux4_1
XFILLER_238_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23197_ _23042_/X _32136_/Q _23215_/S VGND VGND VPWR VPWR _23198_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22148_ _22111_/X _22146_/X _22147_/X _22116_/X VGND VGND VPWR VPWR _22148_/X sky130_fd_sc_hd__a22o_1
X_29813_ _35165_/Q _29351_/X _29817_/S VGND VGND VPWR VPWR _29814_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22079_ _21799_/X _22077_/X _22078_/X _21804_/X VGND VGND VPWR VPWR _22079_/X sky130_fd_sc_hd__a22o_1
X_26956_ _33905_/Q _23364_/X _26960_/S VGND VGND VPWR VPWR _26957_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29744_ _29744_/A VGND VGND VPWR VPWR _35132_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25907_ _25907_/A VGND VGND VPWR VPWR _33410_/D sky130_fd_sc_hd__clkbuf_1
X_29675_ _29675_/A VGND VGND VPWR VPWR _35099_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26887_ _26887_/A VGND VGND VPWR VPWR _33872_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28626_ _27804_/X _34634_/Q _28640_/S VGND VGND VPWR VPWR _28627_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16640_ _17833_/A VGND VGND VPWR VPWR _16640_/X sky130_fd_sc_hd__buf_4
X_25838_ _25838_/A VGND VGND VPWR VPWR _33377_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28557_ _28557_/A VGND VGND VPWR VPWR _34601_/D sky130_fd_sc_hd__clkbuf_1
X_16571_ _32612_/Q _32548_/Q _32484_/Q _35940_/Q _16570_/X _16354_/X VGND VGND VPWR
+ VPWR _16571_/X sky130_fd_sc_hd__mux4_1
XFILLER_245_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25769_ _24933_/X _33345_/Q _25781_/S VGND VGND VPWR VPWR _25770_/A sky130_fd_sc_hd__mux2_1
X_18310_ _18363_/A VGND VGND VPWR VPWR _20261_/A sky130_fd_sc_hd__buf_12
X_27508_ _34135_/Q _27038_/X _27524_/S VGND VGND VPWR VPWR _27509_/A sky130_fd_sc_hd__mux2_1
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19290_ _33136_/Q _36016_/Q _33008_/Q _32944_/Q _19009_/X _19010_/X VGND VGND VPWR
+ VPWR _19290_/X sky130_fd_sc_hd__mux4_1
X_28488_ _28488_/A VGND VGND VPWR VPWR _34568_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_245_1379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18241_ _35220_/Q _35156_/Q _35092_/Q _32276_/Q _16092_/X _16094_/X VGND VGND VPWR
+ VPWR _18241_/X sky130_fd_sc_hd__mux4_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27439_ _27439_/A VGND VGND VPWR VPWR _34102_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30450_ _35467_/Q _29494_/X _30462_/S VGND VGND VPWR VPWR _30451_/A sky130_fd_sc_hd__mux2_1
X_18172_ _18168_/X _18171_/X _17846_/A _17847_/A VGND VGND VPWR VPWR _18187_/B sky130_fd_sc_hd__o211a_1
XFILLER_168_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29109_ _29109_/A VGND VGND VPWR VPWR _34861_/D sky130_fd_sc_hd__clkbuf_1
X_17123_ _17123_/A VGND VGND VPWR VPWR _31987_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30381_ _35434_/Q _29391_/X _30399_/S VGND VGND VPWR VPWR _30382_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32120_ _32889_/CLK _32120_/D VGND VGND VPWR VPWR _32120_/Q sky130_fd_sc_hd__dfxtp_1
X_17054_ _16846_/X _17052_/X _17053_/X _16851_/X VGND VGND VPWR VPWR _17054_/X sky130_fd_sc_hd__a22o_1
XFILLER_87_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16005_ input68/X input67/X VGND VGND VPWR VPWR _17777_/A sky130_fd_sc_hd__nor2b_4
X_32051_ _36019_/CLK _32051_/D VGND VGND VPWR VPWR _32051_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31002_ _35729_/Q input55/X _31002_/S VGND VGND VPWR VPWR _31003_/A sky130_fd_sc_hd__mux2_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35810_ _35810_/CLK _35810_/D VGND VGND VPWR VPWR _35810_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17956_ _17952_/X _17955_/X _17846_/X _17847_/X VGND VGND VPWR VPWR _17973_/B sky130_fd_sc_hd__o211a_1
XFILLER_112_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_936 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35741_ _35805_/CLK _35741_/D VGND VGND VPWR VPWR _35741_/Q sky130_fd_sc_hd__dfxtp_1
X_16907_ _34669_/Q _34605_/Q _34541_/Q _34477_/Q _16586_/X _16587_/X VGND VGND VPWR
+ VPWR _16907_/X sky130_fd_sc_hd__mux4_1
XFILLER_239_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17887_ _17773_/X _17885_/X _17886_/X _17777_/X VGND VGND VPWR VPWR _17887_/X sky130_fd_sc_hd__a22o_1
X_32953_ _35191_/CLK _32953_/D VGND VGND VPWR VPWR _32953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31904_ _23414_/X _36156_/Q _31906_/S VGND VGND VPWR VPWR _31905_/A sky130_fd_sc_hd__mux2_1
X_19626_ _34681_/Q _34617_/Q _34553_/Q _34489_/Q _19592_/X _19593_/X VGND VGND VPWR
+ VPWR _19626_/X sky130_fd_sc_hd__mux4_1
X_35672_ _35800_/CLK _35672_/D VGND VGND VPWR VPWR _35672_/Q sky130_fd_sc_hd__dfxtp_1
X_16838_ _35179_/Q _35115_/Q _35051_/Q _32171_/Q _16657_/X _16658_/X VGND VGND VPWR
+ VPWR _16838_/X sky130_fd_sc_hd__mux4_1
XFILLER_4_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32884_ _32903_/CLK _32884_/D VGND VGND VPWR VPWR _32884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34623_ _35071_/CLK _34623_/D VGND VGND VPWR VPWR _34623_/Q sky130_fd_sc_hd__dfxtp_1
X_31835_ _23246_/X _36123_/Q _31843_/S VGND VGND VPWR VPWR _31836_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19557_ _33079_/Q _32055_/Q _35831_/Q _35767_/Q _19378_/X _19379_/X VGND VGND VPWR
+ VPWR _19557_/X sky130_fd_sc_hd__mux4_1
X_16769_ _16769_/A _16769_/B _16769_/C _16769_/D VGND VGND VPWR VPWR _16770_/A sky130_fd_sc_hd__or4_2
XFILLER_241_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18508_ _18508_/A _18508_/B _18508_/C _18508_/D VGND VGND VPWR VPWR _18509_/A sky130_fd_sc_hd__or4_1
X_31766_ _31766_/A VGND VGND VPWR VPWR _36090_/D sky130_fd_sc_hd__clkbuf_1
X_34554_ _35193_/CLK _34554_/D VGND VGND VPWR VPWR _34554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19488_ _19303_/X _19486_/X _19487_/X _19306_/X VGND VGND VPWR VPWR _19488_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30717_ _30717_/A VGND VGND VPWR VPWR _35593_/D sky130_fd_sc_hd__clkbuf_1
X_33505_ _34593_/CLK _33505_/D VGND VGND VPWR VPWR _33505_/Q sky130_fd_sc_hd__dfxtp_1
X_18439_ _18439_/A VGND VGND VPWR VPWR _32407_/D sky130_fd_sc_hd__buf_4
XFILLER_33_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31697_ _31697_/A VGND VGND VPWR VPWR _36057_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34485_ _34485_/CLK _34485_/D VGND VGND VPWR VPWR _34485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36224_ _36229_/CLK _36224_/D VGND VGND VPWR VPWR _36224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21450_ _34156_/Q _34092_/Q _34028_/Q _33964_/Q _21340_/X _21341_/X VGND VGND VPWR
+ VPWR _21450_/X sky130_fd_sc_hd__mux4_1
XFILLER_222_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33436_ _36211_/CLK _33436_/D VGND VGND VPWR VPWR _33436_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30648_ _35561_/Q _29388_/X _30648_/S VGND VGND VPWR VPWR _30649_/A sky130_fd_sc_hd__mux2_1
X_20401_ _20205_/X _20399_/X _20400_/X _20210_/X VGND VGND VPWR VPWR _20401_/X sky130_fd_sc_hd__a22o_1
XFILLER_222_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33367_ _36055_/CLK _33367_/D VGND VGND VPWR VPWR _33367_/Q sky130_fd_sc_hd__dfxtp_1
X_36155_ _36157_/CLK _36155_/D VGND VGND VPWR VPWR _36155_/Q sky130_fd_sc_hd__dfxtp_1
X_21381_ _32618_/Q _32554_/Q _32490_/Q _35946_/Q _21170_/X _21307_/X VGND VGND VPWR
+ VPWR _21381_/X sky130_fd_sc_hd__mux4_1
X_30579_ _35528_/Q _29484_/X _30597_/S VGND VGND VPWR VPWR _30580_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20332_ _20159_/X _20330_/X _20331_/X _20162_/X VGND VGND VPWR VPWR _20332_/X sky130_fd_sc_hd__a22o_1
X_35106_ _36210_/CLK _35106_/D VGND VGND VPWR VPWR _35106_/Q sky130_fd_sc_hd__dfxtp_1
X_23120_ _23120_/A VGND VGND VPWR VPWR _32099_/D sky130_fd_sc_hd__clkbuf_1
X_32318_ _35902_/CLK _32318_/D VGND VGND VPWR VPWR _32318_/Q sky130_fd_sc_hd__dfxtp_1
X_33298_ _36179_/CLK _33298_/D VGND VGND VPWR VPWR _33298_/Q sky130_fd_sc_hd__dfxtp_1
X_36086_ _36087_/CLK _36086_/D VGND VGND VPWR VPWR _36086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23051_ _23051_/A VGND VGND VPWR VPWR _32074_/D sky130_fd_sc_hd__clkbuf_1
X_35037_ _36219_/CLK _35037_/D VGND VGND VPWR VPWR _35037_/Q sky130_fd_sc_hd__dfxtp_1
X_20263_ _33099_/Q _32075_/Q _35851_/Q _35787_/Q _20084_/X _20085_/X VGND VGND VPWR
+ VPWR _20263_/X sky130_fd_sc_hd__mux4_1
X_32249_ _35191_/CLK _32249_/D VGND VGND VPWR VPWR _32249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22002_ _21998_/X _22001_/X _21765_/X VGND VGND VPWR VPWR _22003_/D sky130_fd_sc_hd__o21ba_1
XTAP_6019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20194_ _20009_/X _20192_/X _20193_/X _20012_/X VGND VGND VPWR VPWR _20194_/X sky130_fd_sc_hd__a22o_1
XFILLER_142_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26810_ _26810_/A VGND VGND VPWR VPWR _33835_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27790_ _27790_/A VGND VGND VPWR VPWR _34245_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26741_ _33803_/Q _23466_/X _26753_/S VGND VGND VPWR VPWR _26742_/A sky130_fd_sc_hd__mux2_1
XTAP_4628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23953_ _23046_/X _32521_/Q _23969_/S VGND VGND VPWR VPWR _23954_/A sky130_fd_sc_hd__mux2_1
X_35939_ _35939_/CLK _35939_/D VGND VGND VPWR VPWR _35939_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22904_ _22903_/X _32027_/Q _22916_/S VGND VGND VPWR VPWR _22905_/A sky130_fd_sc_hd__mux2_1
X_29460_ input37/X VGND VGND VPWR VPWR _29460_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26672_ _33770_/Q _23292_/X _26690_/S VGND VGND VPWR VPWR _26673_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_1024 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23884_ _23884_/A VGND VGND VPWR VPWR _32488_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28411_ _27686_/X _34532_/Q _28421_/S VGND VGND VPWR VPWR _28412_/A sky130_fd_sc_hd__mux2_1
X_25623_ _24917_/X _33276_/Q _25625_/S VGND VGND VPWR VPWR _25624_/A sky130_fd_sc_hd__mux2_1
XFILLER_232_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22835_ _20581_/X _22833_/X _22834_/X _20591_/X VGND VGND VPWR VPWR _22835_/X sky130_fd_sc_hd__a22o_1
X_29391_ input13/X VGND VGND VPWR VPWR _29391_/X sky130_fd_sc_hd__buf_2
XFILLER_112_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28342_ _28342_/A VGND VGND VPWR VPWR _34499_/D sky130_fd_sc_hd__clkbuf_1
X_25554_ _24815_/X _33243_/Q _25562_/S VGND VGND VPWR VPWR _25555_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22766_ _32658_/Q _32594_/Q _32530_/Q _35986_/Q _22582_/X _21477_/A VGND VGND VPWR
+ VPWR _22766_/X sky130_fd_sc_hd__mux4_1
XFILLER_53_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_212_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24505_ _24505_/A VGND VGND VPWR VPWR _32779_/D sky130_fd_sc_hd__clkbuf_1
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21717_ _21400_/X _21715_/X _21716_/X _21403_/X VGND VGND VPWR VPWR _21717_/X sky130_fd_sc_hd__a22o_1
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28273_ _28273_/A VGND VGND VPWR VPWR _34466_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_227_1087 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25485_ _25485_/A VGND VGND VPWR VPWR _33210_/D sky130_fd_sc_hd__clkbuf_1
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22697_ _22697_/A _22697_/B _22697_/C _22697_/D VGND VGND VPWR VPWR _22698_/A sky130_fd_sc_hd__or4_4
XFILLER_201_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_244_1390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27224_ _34003_/Q _27223_/X _27230_/S VGND VGND VPWR VPWR _27225_/A sky130_fd_sc_hd__mux2_1
XFILLER_197_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24436_ _24436_/A VGND VGND VPWR VPWR _32746_/D sky130_fd_sc_hd__clkbuf_1
X_21648_ _21405_/X _21646_/X _21647_/X _21410_/X VGND VGND VPWR VPWR _21648_/X sky130_fd_sc_hd__a22o_1
XFILLER_123_1030 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27155_ input33/X VGND VGND VPWR VPWR _27155_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_240_1287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_193_CLK clkbuf_6_49__f_CLK/X VGND VGND VPWR VPWR _36042_/CLK sky130_fd_sc_hd__clkbuf_16
X_24367_ _23049_/X _32714_/Q _24381_/S VGND VGND VPWR VPWR _24368_/A sky130_fd_sc_hd__mux2_1
X_21579_ _21575_/X _21578_/X _21412_/X VGND VGND VPWR VPWR _21580_/D sky130_fd_sc_hd__o21ba_1
XFILLER_197_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26106_ _26106_/A VGND VGND VPWR VPWR _33504_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23318_ _23318_/A VGND VGND VPWR VPWR _32176_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27086_ _27086_/A VGND VGND VPWR VPWR _33958_/D sky130_fd_sc_hd__clkbuf_1
X_24298_ _24298_/A VGND VGND VPWR VPWR _32681_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26037_ _24930_/X _33472_/Q _26051_/S VGND VGND VPWR VPWR _26038_/A sky130_fd_sc_hd__mux2_1
X_23249_ input61/X VGND VGND VPWR VPWR _23249_/X sky130_fd_sc_hd__buf_4
XFILLER_49_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17810_ _32135_/Q _32327_/Q _32391_/Q _35911_/Q _17633_/X _17774_/X VGND VGND VPWR
+ VPWR _17810_/X sky130_fd_sc_hd__mux4_1
XFILLER_122_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18790_ _18786_/X _18789_/X _18759_/X VGND VGND VPWR VPWR _18791_/D sky130_fd_sc_hd__o21ba_1
XTAP_5830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27988_ _27988_/A VGND VGND VPWR VPWR _34331_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17741_ _17737_/X _17740_/X _17493_/X _17494_/X VGND VGND VPWR VPWR _17756_/B sky130_fd_sc_hd__o211a_1
XFILLER_248_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26939_ _33897_/Q _23289_/X _26939_/S VGND VGND VPWR VPWR _26940_/A sky130_fd_sc_hd__mux2_1
X_29727_ _35124_/Q _29422_/X _29745_/S VGND VGND VPWR VPWR _29728_/A sky130_fd_sc_hd__mux2_1
XTAP_5874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17672_ _35715_/Q _32225_/Q _35587_/Q _35523_/Q _17670_/X _17671_/X VGND VGND VPWR
+ VPWR _17672_/X sky130_fd_sc_hd__mux4_1
XFILLER_48_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29658_ _35092_/Q _29521_/X _29660_/S VGND VGND VPWR VPWR _29659_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19411_ _35443_/Q _35379_/Q _35315_/Q _35251_/Q _19201_/X _19202_/X VGND VGND VPWR
+ VPWR _19411_/X sky130_fd_sc_hd__mux4_1
X_16623_ _34405_/Q _36133_/Q _34277_/Q _34213_/Q _16523_/X _16524_/X VGND VGND VPWR
+ VPWR _16623_/X sky130_fd_sc_hd__mux4_1
X_28609_ _27779_/X _34626_/Q _28619_/S VGND VGND VPWR VPWR _28610_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_1108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29589_ _35059_/Q _29419_/X _29589_/S VGND VGND VPWR VPWR _29590_/A sky130_fd_sc_hd__mux2_1
XFILLER_245_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31620_ _27739_/X _36021_/Q _31636_/S VGND VGND VPWR VPWR _31621_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19342_ _19338_/X _19341_/X _19098_/X VGND VGND VPWR VPWR _19350_/C sky130_fd_sc_hd__o21ba_1
XFILLER_91_1305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16554_ _34659_/Q _34595_/Q _34531_/Q _34467_/Q _16233_/X _16234_/X VGND VGND VPWR
+ VPWR _16554_/X sky130_fd_sc_hd__mux4_1
XFILLER_204_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31551_ _27837_/X _35989_/Q _31551_/S VGND VGND VPWR VPWR _31552_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_1417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19273_ _34671_/Q _34607_/Q _34543_/Q _34479_/Q _19239_/X _19240_/X VGND VGND VPWR
+ VPWR _19273_/X sky130_fd_sc_hd__mux4_1
XFILLER_91_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16485_ _35169_/Q _35105_/Q _35041_/Q _32161_/Q _16304_/X _16305_/X VGND VGND VPWR
+ VPWR _16485_/X sky130_fd_sc_hd__mux4_1
X_18224_ _16030_/X _18222_/X _18223_/X _16041_/X VGND VGND VPWR VPWR _18224_/X sky130_fd_sc_hd__a22o_1
X_30502_ _30502_/A VGND VGND VPWR VPWR _35491_/D sky130_fd_sc_hd__clkbuf_1
X_34270_ _36235_/CLK _34270_/D VGND VGND VPWR VPWR _34270_/Q sky130_fd_sc_hd__dfxtp_1
X_31482_ _31551_/S VGND VGND VPWR VPWR _31501_/S sky130_fd_sc_hd__buf_4
XFILLER_129_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33221_ _34177_/CLK _33221_/D VGND VGND VPWR VPWR _33221_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18155_ _17864_/X _18153_/X _18154_/X _17869_/X VGND VGND VPWR VPWR _18155_/X sky130_fd_sc_hd__a22o_1
XFILLER_191_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30433_ _35459_/Q _29469_/X _30441_/S VGND VGND VPWR VPWR _30434_/A sky130_fd_sc_hd__mux2_1
XFILLER_200_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_184_CLK clkbuf_6_27__f_CLK/X VGND VGND VPWR VPWR _35859_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_15_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_671 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17106_ _17067_/X _17104_/X _17105_/X _17071_/X VGND VGND VPWR VPWR _17106_/X sky130_fd_sc_hd__a22o_1
X_33152_ _36030_/CLK _33152_/D VGND VGND VPWR VPWR _33152_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18086_ _35471_/Q _35407_/Q _35343_/Q _35279_/Q _17960_/X _17961_/X VGND VGND VPWR
+ VPWR _18086_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30364_ _35426_/Q _29367_/X _30378_/S VGND VGND VPWR VPWR _30365_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32103_ _35947_/CLK _32103_/D VGND VGND VPWR VPWR _32103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17037_ _35633_/Q _34993_/Q _34353_/Q _33713_/Q _16791_/X _16792_/X VGND VGND VPWR
+ VPWR _17037_/X sky130_fd_sc_hd__mux4_1
X_33083_ _35835_/CLK _33083_/D VGND VGND VPWR VPWR _33083_/Q sky130_fd_sc_hd__dfxtp_1
X_30295_ _30295_/A VGND VGND VPWR VPWR _35393_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32034_ _35812_/CLK _32034_/D VGND VGND VPWR VPWR _32034_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18988_ _18950_/X _18986_/X _18987_/X _18953_/X VGND VGND VPWR VPWR _18988_/X sky130_fd_sc_hd__a22o_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17939_ _17864_/X _17937_/X _17938_/X _17869_/X VGND VGND VPWR VPWR _17939_/X sky130_fd_sc_hd__a22o_1
XFILLER_6_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33985_ _34177_/CLK _33985_/D VGND VGND VPWR VPWR _33985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35724_ _35724_/CLK _35724_/D VGND VGND VPWR VPWR _35724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20950_ _33886_/Q _33822_/Q _33758_/Q _36062_/Q _20918_/X _20919_/X VGND VGND VPWR
+ VPWR _20950_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32936_ _35755_/CLK _32936_/D VGND VGND VPWR VPWR _32936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19609_ _19605_/X _19608_/X _19432_/X VGND VGND VPWR VPWR _19633_/A sky130_fd_sc_hd__o21ba_1
XFILLER_54_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35655_ _35655_/CLK _35655_/D VGND VGND VPWR VPWR _35655_/Q sky130_fd_sc_hd__dfxtp_1
X_20881_ _20747_/X _20879_/X _20880_/X _20750_/X VGND VGND VPWR VPWR _20881_/X sky130_fd_sc_hd__a22o_1
X_32867_ _32871_/CLK _32867_/D VGND VGND VPWR VPWR _32867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22620_ _32909_/Q _32845_/Q _32781_/Q _32717_/Q _22299_/X _22300_/X VGND VGND VPWR
+ VPWR _22620_/X sky130_fd_sc_hd__mux4_1
X_34606_ _36142_/CLK _34606_/D VGND VGND VPWR VPWR _34606_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31818_ _31818_/A VGND VGND VPWR VPWR _36115_/D sky130_fd_sc_hd__clkbuf_1
X_35586_ _35841_/CLK _35586_/D VGND VGND VPWR VPWR _35586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32798_ _35870_/CLK _32798_/D VGND VGND VPWR VPWR _32798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22551_ _33163_/Q _36043_/Q _33035_/Q _32971_/Q _22368_/X _22369_/X VGND VGND VPWR
+ VPWR _22551_/X sky130_fd_sc_hd__mux4_1
XFILLER_22_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34537_ _34913_/CLK _34537_/D VGND VGND VPWR VPWR _34537_/Q sky130_fd_sc_hd__dfxtp_1
X_31749_ _31749_/A VGND VGND VPWR VPWR _36082_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_179_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21502_ _22561_/A VGND VGND VPWR VPWR _21502_/X sky130_fd_sc_hd__buf_4
X_25270_ _25270_/A VGND VGND VPWR VPWR _25403_/S sky130_fd_sc_hd__buf_8
X_22482_ _32649_/Q _32585_/Q _32521_/Q _35977_/Q _22229_/X _22366_/X VGND VGND VPWR
+ VPWR _22482_/X sky130_fd_sc_hd__mux4_1
XFILLER_21_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34468_ _36136_/CLK _34468_/D VGND VGND VPWR VPWR _34468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24221_ _24221_/A VGND VGND VPWR VPWR _32646_/D sky130_fd_sc_hd__clkbuf_1
X_36207_ _36207_/CLK _36207_/D VGND VGND VPWR VPWR _36207_/Q sky130_fd_sc_hd__dfxtp_1
X_33419_ _33420_/CLK _33419_/D VGND VGND VPWR VPWR _33419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21433_ _35435_/Q _35371_/Q _35307_/Q _35243_/Q _21148_/X _21149_/X VGND VGND VPWR
+ VPWR _21433_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_175_CLK clkbuf_leaf_77_CLK/A VGND VGND VPWR VPWR _35668_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_120_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34399_ _36125_/CLK _34399_/D VGND VGND VPWR VPWR _34399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_1440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21364_ _21047_/X _21362_/X _21363_/X _21050_/X VGND VGND VPWR VPWR _21364_/X sky130_fd_sc_hd__a22o_1
X_36138_ _36140_/CLK _36138_/D VGND VGND VPWR VPWR _36138_/Q sky130_fd_sc_hd__dfxtp_1
X_24152_ _24152_/A VGND VGND VPWR VPWR _32613_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20315_ _20311_/X _20314_/X _20138_/X VGND VGND VPWR VPWR _20337_/A sky130_fd_sc_hd__o21ba_1
X_23103_ _23103_/A VGND VGND VPWR VPWR _32091_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24083_ _24083_/A VGND VGND VPWR VPWR _32582_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36069_ _36070_/CLK _36069_/D VGND VGND VPWR VPWR _36069_/Q sky130_fd_sc_hd__dfxtp_1
X_28960_ _34791_/Q _27087_/X _28964_/S VGND VGND VPWR VPWR _28961_/A sky130_fd_sc_hd__mux2_1
X_21295_ _21052_/X _21293_/X _21294_/X _21057_/X VGND VGND VPWR VPWR _21295_/X sky130_fd_sc_hd__a22o_1
XFILLER_116_782 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20246_ _33419_/Q _33355_/Q _33291_/Q _33227_/Q _20133_/X _20134_/X VGND VGND VPWR
+ VPWR _20246_/X sky130_fd_sc_hd__mux4_1
X_23034_ _23033_/X _32069_/Q _23040_/S VGND VGND VPWR VPWR _23035_/A sky130_fd_sc_hd__mux2_1
X_27911_ _27745_/X _34295_/Q _27923_/S VGND VGND VPWR VPWR _27912_/A sky130_fd_sc_hd__mux2_1
X_28891_ _28891_/A VGND VGND VPWR VPWR _34758_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_235_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27842_ _27639_/X _34262_/Q _27860_/S VGND VGND VPWR VPWR _27843_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20177_ _19852_/X _20175_/X _20176_/X _19857_/X VGND VGND VPWR VPWR _20177_/X sky130_fd_sc_hd__a22o_1
XTAP_5115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27773_ input37/X VGND VGND VPWR VPWR _27773_/X sky130_fd_sc_hd__clkbuf_4
X_24985_ input57/X VGND VGND VPWR VPWR _24985_/X sky130_fd_sc_hd__clkbuf_4
XTAP_4425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29512_ input55/X VGND VGND VPWR VPWR _29512_/X sky130_fd_sc_hd__clkbuf_4
X_26724_ _33795_/Q _23438_/X _26732_/S VGND VGND VPWR VPWR _26725_/A sky130_fd_sc_hd__mux2_1
XTAP_4458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23936_ _23021_/X _32513_/Q _23948_/S VGND VGND VPWR VPWR _23937_/A sky130_fd_sc_hd__mux2_1
XTAP_3724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_218_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_245_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_244_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29443_ _29443_/A VGND VGND VPWR VPWR _35002_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_229_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26655_ _33762_/Q _23268_/X _26669_/S VGND VGND VPWR VPWR _26656_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23867_ _22918_/X _32480_/Q _23885_/S VGND VGND VPWR VPWR _23868_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25606_ _25675_/S VGND VGND VPWR VPWR _25625_/S sky130_fd_sc_hd__buf_4
XFILLER_246_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22818_ _22818_/A VGND VGND VPWR VPWR _36243_/D sky130_fd_sc_hd__clkbuf_1
X_29374_ _34980_/Q _29373_/X _29389_/S VGND VGND VPWR VPWR _29375_/A sky130_fd_sc_hd__mux2_1
X_26586_ _26586_/A VGND VGND VPWR VPWR _33731_/D sky130_fd_sc_hd__clkbuf_1
X_23798_ _23798_/A VGND VGND VPWR VPWR _32384_/D sky130_fd_sc_hd__clkbuf_1
X_28325_ _28325_/A VGND VGND VPWR VPWR _34491_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_246_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25537_ _25537_/A VGND VGND VPWR VPWR _33235_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_213_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22749_ _22745_/X _22748_/X _22457_/X VGND VGND VPWR VPWR _22757_/C sky130_fd_sc_hd__o21ba_1
XFILLER_186_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16270_ _34395_/Q _36123_/Q _34267_/Q _34203_/Q _16170_/X _16171_/X VGND VGND VPWR
+ VPWR _16270_/X sky130_fd_sc_hd__mux4_1
X_28256_ _28256_/A VGND VGND VPWR VPWR _34458_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25468_ _25468_/A VGND VGND VPWR VPWR _33202_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27207_ _27207_/A VGND VGND VPWR VPWR _33997_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_52__f_CLK clkbuf_5_26_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_52__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_8_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24419_ _24419_/A VGND VGND VPWR VPWR _32738_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_166_CLK clkbuf_6_30__f_CLK/X VGND VGND VPWR VPWR _35731_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_16_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28187_ _27754_/X _34426_/Q _28193_/S VGND VGND VPWR VPWR _28188_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25399_ _33171_/Q _23492_/X _25403_/S VGND VGND VPWR VPWR _25400_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27138_ _33975_/Q _27137_/X _27156_/S VGND VGND VPWR VPWR _27139_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19960_ _33923_/Q _33859_/Q _33795_/Q _36099_/Q _19677_/X _19678_/X VGND VGND VPWR
+ VPWR _19960_/X sky130_fd_sc_hd__mux4_1
XFILLER_141_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27069_ input3/X VGND VGND VPWR VPWR _27069_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_10_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18911_ _20099_/A VGND VGND VPWR VPWR _18911_/X sky130_fd_sc_hd__buf_4
XTAP_7040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30080_ _30080_/A VGND VGND VPWR VPWR _35291_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19891_ _34177_/Q _34113_/Q _34049_/Q _33985_/Q _19746_/X _19747_/X VGND VGND VPWR
+ VPWR _19891_/X sky130_fd_sc_hd__mux4_1
XFILLER_180_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18842_ _32867_/Q _32803_/Q _32739_/Q _32675_/Q _18587_/X _18588_/X VGND VGND VPWR
+ VPWR _18842_/X sky130_fd_sc_hd__mux4_1
XTAP_7095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15985_ input66/X VGND VGND VPWR VPWR _16063_/A sky130_fd_sc_hd__clkbuf_16
XTAP_6394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18773_ _32097_/Q _32289_/Q _32353_/Q _35873_/Q _18521_/X _18662_/X VGND VGND VPWR
+ VPWR _18773_/X sky130_fd_sc_hd__mux4_1
XTAP_5660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17724_ _17724_/A _17724_/B _17724_/C _17724_/D VGND VGND VPWR VPWR _17725_/A sky130_fd_sc_hd__or4_4
XFILLER_23_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30982_ _30982_/A VGND VGND VPWR VPWR _35719_/D sky130_fd_sc_hd__clkbuf_1
X_33770_ _33895_/CLK _33770_/D VGND VGND VPWR VPWR _33770_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32721_ _32913_/CLK _32721_/D VGND VGND VPWR VPWR _32721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17655_ _17655_/A VGND VGND VPWR VPWR _32002_/D sky130_fd_sc_hd__buf_4
XFILLER_21_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35440_ _35764_/CLK _35440_/D VGND VGND VPWR VPWR _35440_/Q sky130_fd_sc_hd__dfxtp_1
X_16606_ _16353_/X _16604_/X _16605_/X _16359_/X VGND VGND VPWR VPWR _16606_/X sky130_fd_sc_hd__a22o_1
X_17586_ _17511_/X _17584_/X _17585_/X _17516_/X VGND VGND VPWR VPWR _17586_/X sky130_fd_sc_hd__a22o_1
X_32652_ _36044_/CLK _32652_/D VGND VGND VPWR VPWR _32652_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16537_ _16533_/X _16536_/X _16426_/X VGND VGND VPWR VPWR _16561_/A sky130_fd_sc_hd__o21ba_1
X_19325_ _20151_/A VGND VGND VPWR VPWR _19325_/X sky130_fd_sc_hd__clkbuf_4
X_31603_ _27714_/X _36013_/Q _31615_/S VGND VGND VPWR VPWR _31604_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32583_ _35974_/CLK _32583_/D VGND VGND VPWR VPWR _32583_/Q sky130_fd_sc_hd__dfxtp_1
X_35371_ _35433_/CLK _35371_/D VGND VGND VPWR VPWR _35371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34322_ _36180_/CLK _34322_/D VGND VGND VPWR VPWR _34322_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31534_ _31534_/A VGND VGND VPWR VPWR _35980_/D sky130_fd_sc_hd__clkbuf_1
X_19256_ _19252_/X _19255_/X _19079_/X VGND VGND VPWR VPWR _19280_/A sky130_fd_sc_hd__o21ba_1
X_16468_ _16147_/X _16466_/X _16467_/X _16150_/X VGND VGND VPWR VPWR _16468_/X sky130_fd_sc_hd__a22o_1
X_18207_ _33107_/Q _32083_/Q _35859_/Q _35795_/Q _16079_/X _16080_/X VGND VGND VPWR
+ VPWR _18207_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_157_CLK clkbuf_6_31__f_CLK/X VGND VGND VPWR VPWR _34961_/CLK sky130_fd_sc_hd__clkbuf_16
X_34253_ _34956_/CLK _34253_/D VGND VGND VPWR VPWR _34253_/Q sky130_fd_sc_hd__dfxtp_1
X_19187_ _33389_/Q _33325_/Q _33261_/Q _33197_/Q _19074_/X _19075_/X VGND VGND VPWR
+ VPWR _19187_/X sky130_fd_sc_hd__mux4_1
X_31465_ _31465_/A VGND VGND VPWR VPWR _35947_/D sky130_fd_sc_hd__clkbuf_1
X_16399_ _32863_/Q _32799_/Q _32735_/Q _32671_/Q _16287_/X _16288_/X VGND VGND VPWR
+ VPWR _16399_/X sky130_fd_sc_hd__mux4_1
XFILLER_191_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18138_ _17153_/A _18136_/X _18137_/X _17156_/A VGND VGND VPWR VPWR _18138_/X sky130_fd_sc_hd__a22o_1
X_33204_ _34100_/CLK _33204_/D VGND VGND VPWR VPWR _33204_/Q sky130_fd_sc_hd__dfxtp_1
X_30416_ _35451_/Q _29444_/X _30420_/S VGND VGND VPWR VPWR _30417_/A sky130_fd_sc_hd__mux2_1
X_34184_ _34185_/CLK _34184_/D VGND VGND VPWR VPWR _34184_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31396_ _27807_/X _35915_/Q _31408_/S VGND VGND VPWR VPWR _31397_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_866 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18069_ _33679_/Q _33615_/Q _33551_/Q _33487_/Q _17906_/X _17907_/X VGND VGND VPWR
+ VPWR _18069_/X sky130_fd_sc_hd__mux4_1
X_30347_ _35418_/Q _29342_/X _30357_/S VGND VGND VPWR VPWR _30348_/A sky130_fd_sc_hd__mux2_1
X_33135_ _36144_/CLK _33135_/D VGND VGND VPWR VPWR _33135_/Q sky130_fd_sc_hd__dfxtp_1
X_20100_ _20100_/A VGND VGND VPWR VPWR _20100_/X sky130_fd_sc_hd__buf_4
X_33066_ _35753_/CLK _33066_/D VGND VGND VPWR VPWR _33066_/Q sky130_fd_sc_hd__dfxtp_1
X_21080_ _35425_/Q _35361_/Q _35297_/Q _35233_/Q _20795_/X _20796_/X VGND VGND VPWR
+ VPWR _21080_/X sky130_fd_sc_hd__mux4_1
XFILLER_208_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30278_ _30278_/A VGND VGND VPWR VPWR _35385_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20031_ _20151_/A VGND VGND VPWR VPWR _20031_/X sky130_fd_sc_hd__buf_4
X_32017_ _36207_/CLK _32017_/D VGND VGND VPWR VPWR _32017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_861 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24770_ _23046_/X _32905_/Q _24786_/S VGND VGND VPWR VPWR _24771_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33968_ _34035_/CLK _33968_/D VGND VGND VPWR VPWR _33968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21982_ _32635_/Q _32571_/Q _32507_/Q _35963_/Q _21876_/X _21660_/X VGND VGND VPWR
+ VPWR _21982_/X sky130_fd_sc_hd__mux4_1
XFILLER_67_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_226_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23721_ _22906_/X _32348_/Q _23727_/S VGND VGND VPWR VPWR _23722_/A sky130_fd_sc_hd__mux2_1
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35707_ _35709_/CLK _35707_/D VGND VGND VPWR VPWR _35707_/Q sky130_fd_sc_hd__dfxtp_1
X_32919_ _35993_/CLK _32919_/D VGND VGND VPWR VPWR _32919_/Q sky130_fd_sc_hd__dfxtp_1
X_20933_ _35421_/Q _35357_/Q _35293_/Q _35229_/Q _20795_/X _20796_/X VGND VGND VPWR
+ VPWR _20933_/X sky130_fd_sc_hd__mux4_1
X_33899_ _34091_/CLK _33899_/D VGND VGND VPWR VPWR _33899_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26440_ _26440_/A VGND VGND VPWR VPWR _33662_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23652_ _23008_/X _32317_/Q _23652_/S VGND VGND VPWR VPWR _23653_/A sky130_fd_sc_hd__mux2_1
X_35638_ _35703_/CLK _35638_/D VGND VGND VPWR VPWR _35638_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20864_ _33051_/Q _32027_/Q _35803_/Q _35739_/Q _20667_/X _20669_/X VGND VGND VPWR
+ VPWR _20864_/X sky130_fd_sc_hd__mux4_1
XFILLER_241_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_931 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22603_ _34444_/Q _36172_/Q _34316_/Q _34252_/Q _22535_/X _22536_/X VGND VGND VPWR
+ VPWR _22603_/X sky130_fd_sc_hd__mux4_1
X_26371_ _33630_/Q _23255_/X _26373_/S VGND VGND VPWR VPWR _26372_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23583_ _22906_/X _32284_/Q _23589_/S VGND VGND VPWR VPWR _23584_/A sky130_fd_sc_hd__mux2_1
X_35569_ _35697_/CLK _35569_/D VGND VGND VPWR VPWR _35569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_396_CLK clkbuf_6_41__f_CLK/X VGND VGND VPWR VPWR _35830_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_223_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20795_ _22450_/A VGND VGND VPWR VPWR _20795_/X sky130_fd_sc_hd__buf_6
XFILLER_222_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28110_ _28110_/A _31823_/B VGND VGND VPWR VPWR _28243_/S sky130_fd_sc_hd__nand2_8
XFILLER_139_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25322_ _33134_/Q _23305_/X _25332_/S VGND VGND VPWR VPWR _25323_/A sky130_fd_sc_hd__mux2_1
X_22534_ _22459_/X _22532_/X _22533_/X _22462_/X VGND VGND VPWR VPWR _22534_/X sky130_fd_sc_hd__a22o_1
X_29090_ _29090_/A VGND VGND VPWR VPWR _34852_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28041_ _28041_/A VGND VGND VPWR VPWR _34356_/D sky130_fd_sc_hd__clkbuf_1
X_25253_ _33102_/Q _23475_/X _25259_/S VGND VGND VPWR VPWR _25254_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_148_CLK clkbuf_6_29__f_CLK/X VGND VGND VPWR VPWR _33685_/CLK sky130_fd_sc_hd__clkbuf_16
X_22465_ _34440_/Q _36168_/Q _34312_/Q _34248_/Q _22182_/X _22183_/X VGND VGND VPWR
+ VPWR _22465_/X sky130_fd_sc_hd__mux4_1
XFILLER_154_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24204_ _32638_/Q _23420_/X _24222_/S VGND VGND VPWR VPWR _24205_/A sky130_fd_sc_hd__mux2_1
X_21416_ _33643_/Q _33579_/Q _33515_/Q _33451_/Q _21094_/X _21095_/X VGND VGND VPWR
+ VPWR _21416_/X sky130_fd_sc_hd__mux4_1
X_25184_ _33069_/Q _23302_/X _25196_/S VGND VGND VPWR VPWR _25185_/A sky130_fd_sc_hd__mux2_1
XFILLER_198_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22396_ _22396_/A _22396_/B _22396_/C _22396_/D VGND VGND VPWR VPWR _22397_/A sky130_fd_sc_hd__or4_4
X_24135_ _24135_/A VGND VGND VPWR VPWR _32605_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21347_ _21343_/X _21346_/X _21026_/X VGND VGND VPWR VPWR _21369_/A sky130_fd_sc_hd__o21ba_1
XFILLER_108_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29992_ _35250_/Q _29416_/X _29994_/S VGND VGND VPWR VPWR _29993_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28943_ _34783_/Q _27062_/X _28943_/S VGND VGND VPWR VPWR _28944_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24066_ _23011_/X _32574_/Q _24084_/S VGND VGND VPWR VPWR _24067_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21278_ _20953_/X _21276_/X _21277_/X _20959_/X VGND VGND VPWR VPWR _21278_/X sky130_fd_sc_hd__a22o_1
X_23017_ _23017_/A VGND VGND VPWR VPWR _32063_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20229_ _33098_/Q _32074_/Q _35850_/Q _35786_/Q _20084_/X _20085_/X VGND VGND VPWR
+ VPWR _20229_/X sky130_fd_sc_hd__mux4_1
XFILLER_150_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_320_CLK clkbuf_6_37__f_CLK/X VGND VGND VPWR VPWR _32818_/CLK sky130_fd_sc_hd__clkbuf_16
X_28874_ _34750_/Q _27158_/X _28892_/S VGND VGND VPWR VPWR _28875_/A sky130_fd_sc_hd__mux2_1
XFILLER_235_1186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27825_ input55/X VGND VGND VPWR VPWR _27825_/X sky130_fd_sc_hd__clkbuf_4
XTAP_4211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24968_ _24967_/X _32972_/Q _24983_/S VGND VGND VPWR VPWR _24969_/A sky130_fd_sc_hd__mux2_1
XTAP_4255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27756_ _27756_/A VGND VGND VPWR VPWR _34234_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26707_ _33787_/Q _23411_/X _26711_/S VGND VGND VPWR VPWR _26708_/A sky130_fd_sc_hd__mux2_1
X_23919_ _22996_/X _32505_/Q _23927_/S VGND VGND VPWR VPWR _23920_/A sky130_fd_sc_hd__mux2_1
XTAP_4299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27687_ _27686_/X _34212_/Q _27702_/S VGND VGND VPWR VPWR _27688_/A sky130_fd_sc_hd__mux2_1
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24899_ input26/X VGND VGND VPWR VPWR _24899_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17440_ _34940_/Q _34876_/Q _34812_/Q _34748_/Q _17160_/X _17161_/X VGND VGND VPWR
+ VPWR _17440_/X sky130_fd_sc_hd__mux4_1
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26638_ _33754_/Q _23243_/X _26648_/S VGND VGND VPWR VPWR _26639_/A sky130_fd_sc_hd__mux2_1
XTAP_3598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29426_ input25/X VGND VGND VPWR VPWR _29426_/X sky130_fd_sc_hd__buf_2
XFILLER_73_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_818 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17371_ _17371_/A _17371_/B _17371_/C _17371_/D VGND VGND VPWR VPWR _17372_/A sky130_fd_sc_hd__or4_4
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29357_ input64/X VGND VGND VPWR VPWR _29357_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_387_CLK clkbuf_6_40__f_CLK/X VGND VGND VPWR VPWR _33850_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_60_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26569_ _26569_/A VGND VGND VPWR VPWR _33723_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16322_ _16316_/X _16321_/X _16015_/X VGND VGND VPWR VPWR _16344_/A sky130_fd_sc_hd__o21ba_1
X_19110_ _19463_/A VGND VGND VPWR VPWR _19110_/X sky130_fd_sc_hd__buf_2
XFILLER_159_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28308_ _28308_/A VGND VGND VPWR VPWR _34483_/D sky130_fd_sc_hd__clkbuf_1
X_29288_ _29288_/A VGND VGND VPWR VPWR _34946_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_203_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19041_ _20261_/A VGND VGND VPWR VPWR _19041_/X sky130_fd_sc_hd__buf_4
XFILLER_13_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28239_ _27831_/X _34451_/Q _28243_/S VGND VGND VPWR VPWR _28240_/A sky130_fd_sc_hd__mux2_1
X_16253_ _16018_/X _16251_/X _16252_/X _16027_/X VGND VGND VPWR VPWR _16253_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_139_CLK clkbuf_6_22__f_CLK/X VGND VGND VPWR VPWR _35992_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_16_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31250_ _27791_/X _35846_/Q _31252_/S VGND VGND VPWR VPWR _31251_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16184_ _16180_/X _16183_/X _16015_/X VGND VGND VPWR VPWR _16208_/A sky130_fd_sc_hd__o21ba_1
XFILLER_86_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30201_ _30201_/A VGND VGND VPWR VPWR _35349_/D sky130_fd_sc_hd__clkbuf_1
Xoutput208 _36241_/Q VGND VGND VPWR VPWR D2[59] sky130_fd_sc_hd__buf_2
XFILLER_103_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31181_ _27689_/X _35813_/Q _31189_/S VGND VGND VPWR VPWR _31182_/A sky130_fd_sc_hd__mux2_1
Xoutput219 _32416_/Q VGND VGND VPWR VPWR D3[10] sky130_fd_sc_hd__buf_2
XFILLER_86_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30132_ _35316_/Q _29422_/X _30150_/S VGND VGND VPWR VPWR _30133_/A sky130_fd_sc_hd__mux2_1
X_19943_ _19656_/X _19941_/X _19942_/X _19659_/X VGND VGND VPWR VPWR _19943_/X sky130_fd_sc_hd__a22o_1
X_30063_ _35284_/Q _29521_/X _30065_/S VGND VGND VPWR VPWR _30064_/A sky130_fd_sc_hd__mux2_1
X_34940_ _36157_/CLK _34940_/D VGND VGND VPWR VPWR _34940_/Q sky130_fd_sc_hd__dfxtp_1
X_19874_ _19651_/X _19872_/X _19873_/X _19654_/X VGND VGND VPWR VPWR _19874_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_311_CLK clkbuf_6_50__f_CLK/X VGND VGND VPWR VPWR _35976_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_214_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18825_ _34402_/Q _36130_/Q _34274_/Q _34210_/Q _18823_/X _18824_/X VGND VGND VPWR
+ VPWR _18825_/X sky130_fd_sc_hd__mux4_1
XFILLER_228_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34871_ _35192_/CLK _34871_/D VGND VGND VPWR VPWR _34871_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33822_ _36207_/CLK _33822_/D VGND VGND VPWR VPWR _33822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_1254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18756_ _34912_/Q _34848_/Q _34784_/Q _34720_/Q _18754_/X _18755_/X VGND VGND VPWR
+ VPWR _18756_/X sky130_fd_sc_hd__mux4_1
XTAP_5490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17707_ _17862_/A VGND VGND VPWR VPWR _17707_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_1461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33753_ _33753_/CLK _33753_/D VGND VGND VPWR VPWR _33753_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30965_ _35711_/Q input36/X _30981_/S VGND VGND VPWR VPWR _30966_/A sky130_fd_sc_hd__mux2_1
X_18687_ _20260_/A VGND VGND VPWR VPWR _18687_/X sky130_fd_sc_hd__buf_6
XFILLER_184_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32704_ _32896_/CLK _32704_/D VGND VGND VPWR VPWR _32704_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17638_ _35714_/Q _32224_/Q _35586_/Q _35522_/Q _17317_/X _17318_/X VGND VGND VPWR
+ VPWR _17638_/X sky130_fd_sc_hd__mux4_1
XFILLER_97_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33684_ _33685_/CLK _33684_/D VGND VGND VPWR VPWR _33684_/Q sky130_fd_sc_hd__dfxtp_1
X_30896_ _30896_/A VGND VGND VPWR VPWR _35678_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35423_ _35677_/CLK _35423_/D VGND VGND VPWR VPWR _35423_/Q sky130_fd_sc_hd__dfxtp_1
X_32635_ _35835_/CLK _32635_/D VGND VGND VPWR VPWR _32635_/Q sky130_fd_sc_hd__dfxtp_1
X_17569_ _32896_/Q _32832_/Q _32768_/Q _32704_/Q _17346_/X _17347_/X VGND VGND VPWR
+ VPWR _17569_/X sky130_fd_sc_hd__mux4_1
XFILLER_17_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_378_CLK clkbuf_6_42__f_CLK/X VGND VGND VPWR VPWR _35320_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_182_1060 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19308_ _19302_/X _19307_/X _19098_/X VGND VGND VPWR VPWR _19318_/C sky130_fd_sc_hd__o21ba_1
X_35354_ _35802_/CLK _35354_/D VGND VGND VPWR VPWR _35354_/Q sky130_fd_sc_hd__dfxtp_1
X_20580_ _22365_/A VGND VGND VPWR VPWR _22459_/A sky130_fd_sc_hd__buf_12
XFILLER_182_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32566_ _36023_/CLK _32566_/D VGND VGND VPWR VPWR _32566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34305_ _34690_/CLK _34305_/D VGND VGND VPWR VPWR _34305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_1186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31517_ _31517_/A VGND VGND VPWR VPWR _35972_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19239_ _20298_/A VGND VGND VPWR VPWR _19239_/X sky130_fd_sc_hd__buf_6
X_35285_ _36055_/CLK _35285_/D VGND VGND VPWR VPWR _35285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_939 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32497_ _36017_/CLK _32497_/D VGND VGND VPWR VPWR _32497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22250_ _34434_/Q _36162_/Q _34306_/Q _34242_/Q _22182_/X _22183_/X VGND VGND VPWR
+ VPWR _22250_/X sky130_fd_sc_hd__mux4_1
X_34236_ _35644_/CLK _34236_/D VGND VGND VPWR VPWR _34236_/Q sky130_fd_sc_hd__dfxtp_1
X_31448_ _31448_/A VGND VGND VPWR VPWR _35939_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21201_ _33893_/Q _33829_/Q _33765_/Q _36069_/Q _20918_/X _20919_/X VGND VGND VPWR
+ VPWR _21201_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22181_ _22106_/X _22179_/X _22180_/X _22109_/X VGND VGND VPWR VPWR _22181_/X sky130_fd_sc_hd__a22o_1
XFILLER_219_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31379_ _27782_/X _35907_/Q _31387_/S VGND VGND VPWR VPWR _31380_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34167_ _35704_/CLK _34167_/D VGND VGND VPWR VPWR _34167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_219_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33118_ _33119_/CLK _33118_/D VGND VGND VPWR VPWR _33118_/Q sky130_fd_sc_hd__dfxtp_1
X_21132_ _34147_/Q _34083_/Q _34019_/Q _33955_/Q _20987_/X _20988_/X VGND VGND VPWR
+ VPWR _21132_/X sky130_fd_sc_hd__mux4_1
X_34098_ _34098_/CLK _34098_/D VGND VGND VPWR VPWR _34098_/Q sky130_fd_sc_hd__dfxtp_1
X_25940_ _25940_/A VGND VGND VPWR VPWR _33426_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21063_ _33633_/Q _33569_/Q _33505_/Q _33441_/Q _20741_/X _20742_/X VGND VGND VPWR
+ VPWR _21063_/X sky130_fd_sc_hd__mux4_1
X_33049_ _35801_/CLK _33049_/D VGND VGND VPWR VPWR _33049_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_302_CLK clkbuf_6_51__f_CLK/X VGND VGND VPWR VPWR _35525_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_235_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20014_ _20008_/X _20013_/X _19804_/X VGND VGND VPWR VPWR _20024_/C sky130_fd_sc_hd__o21ba_1
XFILLER_141_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25871_ _25871_/A VGND VGND VPWR VPWR _33393_/D sky130_fd_sc_hd__clkbuf_1
X_27610_ _27637_/S VGND VGND VPWR VPWR _27629_/S sky130_fd_sc_hd__buf_4
X_24822_ _24821_/X _32925_/Q _24828_/S VGND VGND VPWR VPWR _24823_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28590_ _27751_/X _34617_/Q _28598_/S VGND VGND VPWR VPWR _28591_/A sky130_fd_sc_hd__mux2_1
XFILLER_246_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27541_ _34151_/Q _27087_/X _27545_/S VGND VGND VPWR VPWR _27542_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24753_ _23021_/X _32897_/Q _24765_/S VGND VGND VPWR VPWR _24754_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21965_ _35194_/Q _35130_/Q _35066_/Q _32250_/Q _21963_/X _21964_/X VGND VGND VPWR
+ VPWR _21965_/X sky130_fd_sc_hd__mux4_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23704_ input83/X input89/X VGND VGND VPWR VPWR _27232_/A sky130_fd_sc_hd__or2b_2
XFILLER_27_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27472_ _27472_/A VGND VGND VPWR VPWR _34118_/D sky130_fd_sc_hd__clkbuf_1
X_20916_ _20740_/X _20914_/X _20915_/X _20745_/X VGND VGND VPWR VPWR _20916_/X sky130_fd_sc_hd__a22o_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24684_ _22918_/X _32864_/Q _24702_/S VGND VGND VPWR VPWR _24685_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_226_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21896_ _21753_/X _21894_/X _21895_/X _21756_/X VGND VGND VPWR VPWR _21896_/X sky130_fd_sc_hd__a22o_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29211_ _34910_/Q _27059_/X _29213_/S VGND VGND VPWR VPWR _29212_/A sky130_fd_sc_hd__mux2_1
XFILLER_202_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26423_ _26423_/A VGND VGND VPWR VPWR _33654_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23635_ _23635_/A VGND VGND VPWR VPWR _32308_/D sky130_fd_sc_hd__clkbuf_1
X_20847_ _33371_/Q _33307_/Q _33243_/Q _33179_/Q _20602_/X _20603_/X VGND VGND VPWR
+ VPWR _20847_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_369_CLK clkbuf_6_43__f_CLK/X VGND VGND VPWR VPWR _35769_/CLK sky130_fd_sc_hd__clkbuf_16
X_29142_ _29142_/A VGND VGND VPWR VPWR _34877_/D sky130_fd_sc_hd__clkbuf_1
X_26354_ _26486_/S VGND VGND VPWR VPWR _26373_/S sky130_fd_sc_hd__buf_6
X_23566_ _23566_/A VGND VGND VPWR VPWR _32277_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20778_ _33625_/Q _33561_/Q _33497_/Q _33433_/Q _20741_/X _20742_/X VGND VGND VPWR
+ VPWR _20778_/X sky130_fd_sc_hd__mux4_1
XFILLER_196_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25305_ _33126_/Q _23280_/X _25311_/S VGND VGND VPWR VPWR _25306_/A sky130_fd_sc_hd__mux2_1
X_29073_ _29073_/A VGND VGND VPWR VPWR _34844_/D sky130_fd_sc_hd__clkbuf_1
X_22517_ _22511_/X _22516_/X _22438_/X VGND VGND VPWR VPWR _22541_/A sky130_fd_sc_hd__o21ba_1
XFILLER_128_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26285_ _26285_/A VGND VGND VPWR VPWR _33589_/D sky130_fd_sc_hd__clkbuf_1
X_23497_ _23497_/A VGND VGND VPWR VPWR _32244_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28024_ _28024_/A VGND VGND VPWR VPWR _34348_/D sky130_fd_sc_hd__clkbuf_1
X_25236_ _33094_/Q _23447_/X _25238_/S VGND VGND VPWR VPWR _25237_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22448_ _22442_/X _22445_/X _22446_/X _22447_/X VGND VGND VPWR VPWR _22473_/B sky130_fd_sc_hd__o211a_2
XFILLER_171_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25167_ _33061_/Q _23277_/X _25175_/S VGND VGND VPWR VPWR _25168_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_1448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22379_ _22372_/X _22378_/X _22093_/X _22094_/X VGND VGND VPWR VPWR _22396_/B sky130_fd_sc_hd__o211a_1
XFILLER_163_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24118_ _24118_/A _30877_/B VGND VGND VPWR VPWR _24251_/S sky130_fd_sc_hd__nor2_8
XFILLER_151_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25098_ _25098_/A VGND VGND VPWR VPWR _33029_/D sky130_fd_sc_hd__clkbuf_1
X_29975_ _30065_/S VGND VGND VPWR VPWR _29994_/S sky130_fd_sc_hd__buf_6
XFILLER_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28926_ _28926_/A VGND VGND VPWR VPWR _34774_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16940_ _17999_/A VGND VGND VPWR VPWR _16940_/X sky130_fd_sc_hd__clkbuf_4
X_24049_ _22987_/X _32566_/Q _24063_/S VGND VGND VPWR VPWR _24050_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16871_ _16650_/X _16869_/X _16870_/X _16653_/X VGND VGND VPWR VPWR _16871_/X sky130_fd_sc_hd__a22o_1
X_28857_ _34742_/Q _27134_/X _28871_/S VGND VGND VPWR VPWR _28858_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18610_ _18391_/X _18608_/X _18609_/X _18401_/X VGND VGND VPWR VPWR _18610_/X sky130_fd_sc_hd__a22o_1
X_27808_ _27807_/X _34251_/Q _27826_/S VGND VGND VPWR VPWR _27809_/A sky130_fd_sc_hd__mux2_1
XTAP_4030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19590_ _19303_/X _19588_/X _19589_/X _19306_/X VGND VGND VPWR VPWR _19590_/X sky130_fd_sc_hd__a22o_1
X_28788_ _29797_/A _31688_/A VGND VGND VPWR VPWR _28921_/S sky130_fd_sc_hd__nor2_8
XTAP_4052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18541_ _18537_/X _18540_/X _18404_/X VGND VGND VPWR VPWR _18542_/D sky130_fd_sc_hd__o21ba_1
XTAP_4074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1030 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27739_ input25/X VGND VGND VPWR VPWR _27739_/X sky130_fd_sc_hd__buf_2
XTAP_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18472_ _34392_/Q _36120_/Q _34264_/Q _34200_/Q _18470_/X _18471_/X VGND VGND VPWR
+ VPWR _18472_/X sky130_fd_sc_hd__mux4_1
X_30750_ _35609_/Q input34/X _30762_/S VGND VGND VPWR VPWR _30751_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29409_ _29409_/A VGND VGND VPWR VPWR _34991_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17423_ _32892_/Q _32828_/Q _32764_/Q _32700_/Q _17346_/X _17347_/X VGND VGND VPWR
+ VPWR _17423_/X sky130_fd_sc_hd__mux4_1
XFILLER_205_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30681_ _30681_/A VGND VGND VPWR VPWR _35576_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32420_ _33828_/CLK _32420_/D VGND VGND VPWR VPWR _32420_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17354_ _17862_/A VGND VGND VPWR VPWR _17354_/X sky130_fd_sc_hd__buf_6
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16305_ _17011_/A VGND VGND VPWR VPWR _16305_/X sky130_fd_sc_hd__buf_6
XFILLER_159_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32351_ _35871_/CLK _32351_/D VGND VGND VPWR VPWR _32351_/Q sky130_fd_sc_hd__dfxtp_1
X_17285_ _35704_/Q _32213_/Q _35576_/Q _35512_/Q _16964_/X _16965_/X VGND VGND VPWR
+ VPWR _17285_/X sky130_fd_sc_hd__mux4_1
XFILLER_146_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16236_ _35162_/Q _35098_/Q _35034_/Q _32154_/Q _16083_/X _16085_/X VGND VGND VPWR
+ VPWR _16236_/X sky130_fd_sc_hd__mux4_1
X_31302_ _31302_/A VGND VGND VPWR VPWR _35870_/D sky130_fd_sc_hd__clkbuf_1
X_19024_ _35432_/Q _35368_/Q _35304_/Q _35240_/Q _18848_/X _18849_/X VGND VGND VPWR
+ VPWR _19024_/X sky130_fd_sc_hd__mux4_1
XFILLER_70_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35070_ _36100_/CLK _35070_/D VGND VGND VPWR VPWR _35070_/Q sky130_fd_sc_hd__dfxtp_1
X_32282_ _35995_/CLK _32282_/D VGND VGND VPWR VPWR _32282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31233_ _31281_/S VGND VGND VPWR VPWR _31252_/S sky130_fd_sc_hd__clkbuf_8
X_34021_ _34149_/CLK _34021_/D VGND VGND VPWR VPWR _34021_/Q sky130_fd_sc_hd__dfxtp_1
X_16167_ _34648_/Q _34584_/Q _34520_/Q _34456_/Q _16079_/X _16080_/X VGND VGND VPWR
+ VPWR _16167_/X sky130_fd_sc_hd__mux4_1
XFILLER_173_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31164_ _27664_/X _35805_/Q _31168_/S VGND VGND VPWR VPWR _31165_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16098_ _17161_/A VGND VGND VPWR VPWR _16098_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_29_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30115_ _35308_/Q _29398_/X _30129_/S VGND VGND VPWR VPWR _30116_/A sky130_fd_sc_hd__mux2_1
X_19926_ _33922_/Q _33858_/Q _33794_/Q _36098_/Q _19677_/X _19678_/X VGND VGND VPWR
+ VPWR _19926_/X sky130_fd_sc_hd__mux4_1
X_35972_ _35973_/CLK _35972_/D VGND VGND VPWR VPWR _35972_/Q sky130_fd_sc_hd__dfxtp_1
X_31095_ _35773_/Q input33/X _31095_/S VGND VGND VPWR VPWR _31096_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_214_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30046_ _30046_/A VGND VGND VPWR VPWR _35275_/D sky130_fd_sc_hd__clkbuf_1
X_34923_ _34924_/CLK _34923_/D VGND VGND VPWR VPWR _34923_/Q sky130_fd_sc_hd__dfxtp_1
X_19857_ _20210_/A VGND VGND VPWR VPWR _19857_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_190_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18808_ _18653_/X _18806_/X _18807_/X _18659_/X VGND VGND VPWR VPWR _18808_/X sky130_fd_sc_hd__a22o_1
XFILLER_18_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34854_ _34920_/CLK _34854_/D VGND VGND VPWR VPWR _34854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19788_ _33150_/Q _36030_/Q _33022_/Q _32958_/Q _19715_/X _19716_/X VGND VGND VPWR
+ VPWR _19788_/X sky130_fd_sc_hd__mux4_1
XFILLER_110_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33805_ _36109_/CLK _33805_/D VGND VGND VPWR VPWR _33805_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18739_ _20299_/A VGND VGND VPWR VPWR _18739_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_83_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1084 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34785_ _34915_/CLK _34785_/D VGND VGND VPWR VPWR _34785_/Q sky130_fd_sc_hd__dfxtp_1
X_31997_ _34405_/CLK _31997_/D VGND VGND VPWR VPWR _31997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33736_ _35724_/CLK _33736_/D VGND VGND VPWR VPWR _33736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_1291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21750_ _21603_/X _21748_/X _21749_/X _21606_/X VGND VGND VPWR VPWR _21750_/X sky130_fd_sc_hd__a22o_1
X_30948_ _35703_/Q input27/X _30960_/S VGND VGND VPWR VPWR _30949_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20701_ _21763_/A VGND VGND VPWR VPWR _20701_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_58_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_1008 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_558 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33667_ _34942_/CLK _33667_/D VGND VGND VPWR VPWR _33667_/Q sky130_fd_sc_hd__dfxtp_1
X_21681_ _21603_/X _21677_/X _21680_/X _21606_/X VGND VGND VPWR VPWR _21681_/X sky130_fd_sc_hd__a22o_1
X_30879_ _35670_/Q input1/X _30897_/S VGND VGND VPWR VPWR _30880_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35406_ _35855_/CLK _35406_/D VGND VGND VPWR VPWR _35406_/Q sky130_fd_sc_hd__dfxtp_1
X_23420_ input35/X VGND VGND VPWR VPWR _23420_/X sky130_fd_sc_hd__buf_4
X_20632_ _22586_/A VGND VGND VPWR VPWR _20632_/X sky130_fd_sc_hd__buf_6
X_32618_ _36010_/CLK _32618_/D VGND VGND VPWR VPWR _32618_/Q sky130_fd_sc_hd__dfxtp_1
X_33598_ _34174_/CLK _33598_/D VGND VGND VPWR VPWR _33598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35337_ _35466_/CLK _35337_/D VGND VGND VPWR VPWR _35337_/Q sky130_fd_sc_hd__dfxtp_1
X_23351_ _32192_/Q _23277_/X _23359_/S VGND VGND VPWR VPWR _23352_/A sky130_fd_sc_hd__mux2_1
X_20563_ _35733_/Q _32245_/Q _35605_/Q _35541_/Q _18293_/X _18295_/X VGND VGND VPWR
+ VPWR _20563_/X sky130_fd_sc_hd__mux4_1
X_32549_ _35943_/CLK _32549_/D VGND VGND VPWR VPWR _32549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22302_ _22020_/X _22298_/X _22301_/X _22024_/X VGND VGND VPWR VPWR _22302_/X sky130_fd_sc_hd__a22o_1
XFILLER_109_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26070_ _24979_/X _33488_/Q _26072_/S VGND VGND VPWR VPWR _26071_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35268_ _35843_/CLK _35268_/D VGND VGND VPWR VPWR _35268_/Q sky130_fd_sc_hd__dfxtp_1
X_23282_ _23282_/A VGND VGND VPWR VPWR _32166_/D sky130_fd_sc_hd__clkbuf_1
X_20494_ _20212_/X _20492_/X _20493_/X _20215_/X VGND VGND VPWR VPWR _20494_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25021_ _25021_/A VGND VGND VPWR VPWR _32992_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22233_ _22586_/A VGND VGND VPWR VPWR _22233_/X sky130_fd_sc_hd__buf_6
X_34219_ _36141_/CLK _34219_/D VGND VGND VPWR VPWR _34219_/Q sky130_fd_sc_hd__dfxtp_1
X_35199_ _36101_/CLK _35199_/D VGND VGND VPWR VPWR _35199_/Q sky130_fd_sc_hd__dfxtp_1
X_22164_ _22158_/X _22163_/X _22085_/X VGND VGND VPWR VPWR _22188_/A sky130_fd_sc_hd__o21ba_1
XFILLER_246_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21115_ _20892_/X _21113_/X _21114_/X _20895_/X VGND VGND VPWR VPWR _21115_/X sky130_fd_sc_hd__a22o_1
XTAP_6938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29760_ _35140_/Q _29472_/X _29766_/S VGND VGND VPWR VPWR _29761_/A sky130_fd_sc_hd__mux2_1
X_22095_ _22089_/X _22092_/X _22093_/X _22094_/X VGND VGND VPWR VPWR _22120_/B sky130_fd_sc_hd__o211a_1
X_26972_ _26972_/A VGND VGND VPWR VPWR _33912_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28711_ _34674_/Q _27121_/X _28713_/S VGND VGND VPWR VPWR _28712_/A sky130_fd_sc_hd__mux2_1
X_25923_ _24961_/X _33418_/Q _25937_/S VGND VGND VPWR VPWR _25924_/A sky130_fd_sc_hd__mux2_1
X_21046_ _21041_/X _21044_/X _21045_/X VGND VGND VPWR VPWR _21061_/C sky130_fd_sc_hd__o21ba_1
X_29691_ _35107_/Q _29370_/X _29703_/S VGND VGND VPWR VPWR _29692_/A sky130_fd_sc_hd__mux2_1
XFILLER_219_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28642_ _27828_/X _34642_/Q _28648_/S VGND VGND VPWR VPWR _28643_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25854_ _25854_/A VGND VGND VPWR VPWR _33385_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24805_ _24805_/A VGND VGND VPWR VPWR _32919_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_228_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25785_ _25785_/A VGND VGND VPWR VPWR _33352_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_189_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28573_ _27726_/X _34609_/Q _28577_/S VGND VGND VPWR VPWR _28574_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22997_ _22996_/X _32057_/Q _23009_/S VGND VGND VPWR VPWR _22998_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_1214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27524_ _34143_/Q _27062_/X _27524_/S VGND VGND VPWR VPWR _27525_/A sky130_fd_sc_hd__mux2_1
X_24736_ _22996_/X _32889_/Q _24744_/S VGND VGND VPWR VPWR _24737_/A sky130_fd_sc_hd__mux2_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21948_ _32890_/Q _32826_/Q _32762_/Q _32698_/Q _21946_/X _21947_/X VGND VGND VPWR
+ VPWR _21948_/X sky130_fd_sc_hd__mux4_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27455_ _34110_/Q _27158_/X _27473_/S VGND VGND VPWR VPWR _27456_/A sky130_fd_sc_hd__mux2_1
XFILLER_242_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24667_ _22894_/X _32856_/Q _24681_/S VGND VGND VPWR VPWR _24668_/A sky130_fd_sc_hd__mux2_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21879_ _21659_/X _21877_/X _21878_/X _21665_/X VGND VGND VPWR VPWR _21879_/X sky130_fd_sc_hd__a22o_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26406_ _26406_/A VGND VGND VPWR VPWR _33646_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23618_ _23618_/A VGND VGND VPWR VPWR _32300_/D sky130_fd_sc_hd__clkbuf_1
X_27386_ _27386_/A VGND VGND VPWR VPWR _34077_/D sky130_fd_sc_hd__clkbuf_1
X_24598_ _24598_/A VGND VGND VPWR VPWR _32823_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26337_ _26337_/A VGND VGND VPWR VPWR _33614_/D sky130_fd_sc_hd__clkbuf_1
X_29125_ _34869_/Q _27131_/X _29141_/S VGND VGND VPWR VPWR _29126_/A sky130_fd_sc_hd__mux2_1
X_23549_ _32269_/Q _23472_/X _23557_/S VGND VGND VPWR VPWR _23550_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29056_ _34837_/Q _27229_/X _29056_/S VGND VGND VPWR VPWR _29057_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17070_ _32882_/Q _32818_/Q _32754_/Q _32690_/Q _16993_/X _16994_/X VGND VGND VPWR
+ VPWR _17070_/X sky130_fd_sc_hd__mux4_1
XFILLER_155_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26268_ _26268_/A VGND VGND VPWR VPWR _33581_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16021_ _16063_/A VGND VGND VPWR VPWR _17766_/A sky130_fd_sc_hd__buf_12
X_25219_ _25267_/S VGND VGND VPWR VPWR _25238_/S sky130_fd_sc_hd__buf_4
X_28007_ _28007_/A VGND VGND VPWR VPWR _34340_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26199_ _24970_/X _33549_/Q _26207_/S VGND VGND VPWR VPWR _26200_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_780 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_70_CLK clkbuf_leaf_73_CLK/A VGND VGND VPWR VPWR _35871_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_178_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17972_ _17968_/X _17971_/X _17871_/X VGND VGND VPWR VPWR _17973_/D sky130_fd_sc_hd__o21ba_1
XFILLER_124_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29958_ _29958_/A VGND VGND VPWR VPWR _35233_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19711_ _19707_/X _19710_/X _19432_/X VGND VGND VPWR VPWR _19743_/A sky130_fd_sc_hd__o21ba_1
X_28909_ _34767_/Q _27211_/X _28913_/S VGND VGND VPWR VPWR _28910_/A sky130_fd_sc_hd__mux2_1
X_16923_ _17982_/A VGND VGND VPWR VPWR _16923_/X sky130_fd_sc_hd__buf_6
XFILLER_242_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29889_ _35201_/Q _29463_/X _29901_/S VGND VGND VPWR VPWR _29890_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_1043 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31920_ _31920_/A VGND VGND VPWR VPWR _36163_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19642_ _32634_/Q _32570_/Q _32506_/Q _35962_/Q _19576_/X _19360_/X VGND VGND VPWR
+ VPWR _19642_/X sky130_fd_sc_hd__mux4_1
X_16854_ _33388_/Q _33324_/Q _33260_/Q _33196_/Q _16774_/X _16775_/X VGND VGND VPWR
+ VPWR _16854_/X sky130_fd_sc_hd__mux4_1
XFILLER_226_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19573_ _33912_/Q _33848_/Q _33784_/Q _36088_/Q _19324_/X _19325_/X VGND VGND VPWR
+ VPWR _19573_/X sky130_fd_sc_hd__mux4_1
X_31851_ _31851_/A VGND VGND VPWR VPWR _36130_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16785_ _32874_/Q _32810_/Q _32746_/Q _32682_/Q _16640_/X _16641_/X VGND VGND VPWR
+ VPWR _16785_/X sky130_fd_sc_hd__mux4_1
XFILLER_59_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18524_ _18330_/X _18522_/X _18523_/X _18341_/X VGND VGND VPWR VPWR _18524_/X sky130_fd_sc_hd__a22o_1
X_30802_ _35634_/Q input21/X _30804_/S VGND VGND VPWR VPWR _30803_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34570_ _35208_/CLK _34570_/D VGND VGND VPWR VPWR _34570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31782_ _36098_/Q input39/X _31792_/S VGND VGND VPWR VPWR _31783_/A sky130_fd_sc_hd__mux2_1
XTAP_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33521_ _33904_/CLK _33521_/D VGND VGND VPWR VPWR _33521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18455_ _18318_/X _18453_/X _18454_/X _18327_/X VGND VGND VPWR VPWR _18455_/X sky130_fd_sc_hd__a22o_1
X_30733_ _30733_/A VGND VGND VPWR VPWR _35601_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_968 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_1459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36240_ _36242_/CLK _36240_/D VGND VGND VPWR VPWR _36240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17406_ _34172_/Q _34108_/Q _34044_/Q _33980_/Q _17093_/X _17094_/X VGND VGND VPWR
+ VPWR _17406_/X sky130_fd_sc_hd__mux4_1
XFILLER_226_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33452_ _34093_/CLK _33452_/D VGND VGND VPWR VPWR _33452_/Q sky130_fd_sc_hd__dfxtp_1
X_18386_ _35158_/Q _35094_/Q _35030_/Q _32150_/Q _18383_/X _18385_/X VGND VGND VPWR
+ VPWR _18386_/X sky130_fd_sc_hd__mux4_1
X_30664_ _30664_/A VGND VGND VPWR VPWR _35568_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32403_ _35922_/CLK _32403_/D VGND VGND VPWR VPWR _32403_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36171_ _36171_/CLK _36171_/D VGND VGND VPWR VPWR _36171_/Q sky130_fd_sc_hd__dfxtp_1
X_17337_ _17199_/X _17335_/X _17336_/X _17204_/X VGND VGND VPWR VPWR _17337_/X sky130_fd_sc_hd__a22o_1
X_30595_ _35536_/Q _29509_/X _30597_/S VGND VGND VPWR VPWR _30596_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33383_ _36072_/CLK _33383_/D VGND VGND VPWR VPWR _33383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_1088 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35122_ _35828_/CLK _35122_/D VGND VGND VPWR VPWR _35122_/Q sky130_fd_sc_hd__dfxtp_1
X_32334_ _35921_/CLK _32334_/D VGND VGND VPWR VPWR _32334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17268_ _17268_/A VGND VGND VPWR VPWR _31991_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19007_ _20066_/A VGND VGND VPWR VPWR _19007_/X sky130_fd_sc_hd__clkbuf_4
X_16219_ _33114_/Q _35994_/Q _32986_/Q _32922_/Q _16024_/X _16025_/X VGND VGND VPWR
+ VPWR _16219_/X sky130_fd_sc_hd__mux4_1
XFILLER_134_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35053_ _35181_/CLK _35053_/D VGND VGND VPWR VPWR _35053_/Q sky130_fd_sc_hd__dfxtp_1
X_32265_ _35210_/CLK _32265_/D VGND VGND VPWR VPWR _32265_/Q sky130_fd_sc_hd__dfxtp_1
X_17199_ _17905_/A VGND VGND VPWR VPWR _17199_/X sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_505_CLK clkbuf_leaf_2_CLK/A VGND VGND VPWR VPWR _33827_/CLK sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_61_CLK clkbuf_leaf_61_CLK/A VGND VGND VPWR VPWR _32913_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_155_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34004_ _34773_/CLK _34004_/D VGND VGND VPWR VPWR _34004_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31216_ _31216_/A VGND VGND VPWR VPWR _35829_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32196_ _35691_/CLK _32196_/D VGND VGND VPWR VPWR _32196_/Q sky130_fd_sc_hd__dfxtp_1
X_31147_ _31147_/A _31147_/B VGND VGND VPWR VPWR _31148_/A sky130_fd_sc_hd__or2_1
XFILLER_9_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19909_ _35457_/Q _35393_/Q _35329_/Q _35265_/Q _19907_/X _19908_/X VGND VGND VPWR
+ VPWR _19909_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_6_29__f_CLK clkbuf_5_14_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_29__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_190_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31078_ _31078_/A VGND VGND VPWR VPWR _35764_/D sky130_fd_sc_hd__clkbuf_1
X_35955_ _35955_/CLK _35955_/D VGND VGND VPWR VPWR _35955_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34906_ _34911_/CLK _34906_/D VGND VGND VPWR VPWR _34906_/Q sky130_fd_sc_hd__dfxtp_1
X_30029_ _30029_/A VGND VGND VPWR VPWR _35267_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22920_ _22918_/X _32032_/Q _22947_/S VGND VGND VPWR VPWR _22921_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35886_ _35951_/CLK _35886_/D VGND VGND VPWR VPWR _35886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_232_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34837_ _36181_/CLK _34837_/D VGND VGND VPWR VPWR _34837_/Q sky130_fd_sc_hd__dfxtp_1
X_22851_ _20618_/X _22849_/X _22850_/X _20627_/X VGND VGND VPWR VPWR _22851_/X sky130_fd_sc_hd__a22o_1
XFILLER_42_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21802_ _33654_/Q _33590_/Q _33526_/Q _33462_/Q _21800_/X _21801_/X VGND VGND VPWR
+ VPWR _21802_/X sky130_fd_sc_hd__mux4_1
X_25570_ _25570_/A VGND VGND VPWR VPWR _33250_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34768_ _34897_/CLK _34768_/D VGND VGND VPWR VPWR _34768_/Q sky130_fd_sc_hd__dfxtp_1
X_22782_ _20648_/X _22780_/X _22781_/X _20658_/X VGND VGND VPWR VPWR _22782_/X sky130_fd_sc_hd__a22o_1
XFILLER_231_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24521_ _24521_/A VGND VGND VPWR VPWR _32787_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21733_ _21726_/X _21731_/X _21732_/X VGND VGND VPWR VPWR _21767_/A sky130_fd_sc_hd__o21ba_1
X_33719_ _35768_/CLK _33719_/D VGND VGND VPWR VPWR _33719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34699_ _36167_/CLK _34699_/D VGND VGND VPWR VPWR _34699_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27240_ _34008_/Q _27041_/X _27254_/S VGND VGND VPWR VPWR _27241_/A sky130_fd_sc_hd__mux2_1
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24452_ _24452_/A VGND VGND VPWR VPWR _32754_/D sky130_fd_sc_hd__clkbuf_1
X_21664_ _33138_/Q _36018_/Q _33010_/Q _32946_/Q _21662_/X _21663_/X VGND VGND VPWR
+ VPWR _21664_/X sky130_fd_sc_hd__mux4_1
XFILLER_24_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23403_ _32213_/Q _23402_/X _23418_/S VGND VGND VPWR VPWR _23404_/A sky130_fd_sc_hd__mux2_1
X_27171_ input39/X VGND VGND VPWR VPWR _27171_/X sky130_fd_sc_hd__clkbuf_4
X_20615_ _22438_/A VGND VGND VPWR VPWR _20615_/X sky130_fd_sc_hd__buf_4
XFILLER_131_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24383_ _23073_/X _32722_/Q _24389_/S VGND VGND VPWR VPWR _24384_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_894 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21595_ _32880_/Q _32816_/Q _32752_/Q _32688_/Q _21593_/X _21594_/X VGND VGND VPWR
+ VPWR _21595_/X sky130_fd_sc_hd__mux4_1
XFILLER_201_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26122_ _26122_/A VGND VGND VPWR VPWR _33512_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23334_ _23334_/A VGND VGND VPWR VPWR _32184_/D sky130_fd_sc_hd__clkbuf_1
X_20546_ _20542_/X _20545_/X _20171_/A VGND VGND VPWR VPWR _20547_/D sky130_fd_sc_hd__o21ba_1
XFILLER_193_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26053_ _26080_/S VGND VGND VPWR VPWR _26072_/S sky130_fd_sc_hd__buf_4
XFILLER_193_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23265_ input3/X VGND VGND VPWR VPWR _23265_/X sky130_fd_sc_hd__buf_4
X_20477_ _33106_/Q _32082_/Q _35858_/Q _35794_/Q _18379_/X _18380_/X VGND VGND VPWR
+ VPWR _20477_/X sky130_fd_sc_hd__mux4_1
XFILLER_193_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_52_CLK clkbuf_leaf_57_CLK/A VGND VGND VPWR VPWR _35945_/CLK sky130_fd_sc_hd__clkbuf_16
X_25004_ _25004_/A VGND VGND VPWR VPWR _32984_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22216_ _34433_/Q _36161_/Q _34305_/Q _34241_/Q _22182_/X _22183_/X VGND VGND VPWR
+ VPWR _22216_/X sky130_fd_sc_hd__mux4_1
XFILLER_193_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_558 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23196_ _23223_/S VGND VGND VPWR VPWR _23215_/S sky130_fd_sc_hd__buf_4
XTAP_6702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29812_ _29812_/A VGND VGND VPWR VPWR _35164_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22147_ _34943_/Q _34879_/Q _34815_/Q _34751_/Q _22113_/X _22114_/X VGND VGND VPWR
+ VPWR _22147_/X sky130_fd_sc_hd__mux4_1
XFILLER_121_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29743_ _35132_/Q _29447_/X _29745_/S VGND VGND VPWR VPWR _29744_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22078_ _34174_/Q _34110_/Q _34046_/Q _33982_/Q _22046_/X _22047_/X VGND VGND VPWR
+ VPWR _22078_/X sky130_fd_sc_hd__mux4_1
X_26955_ _26955_/A VGND VGND VPWR VPWR _33904_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25906_ _24936_/X _33410_/Q _25916_/S VGND VGND VPWR VPWR _25907_/A sky130_fd_sc_hd__mux2_1
X_21029_ _33120_/Q _36000_/Q _32992_/Q _32928_/Q _20956_/X _20957_/X VGND VGND VPWR
+ VPWR _21029_/X sky130_fd_sc_hd__mux4_1
X_29674_ _35099_/Q _29345_/X _29682_/S VGND VGND VPWR VPWR _29675_/A sky130_fd_sc_hd__mux2_1
X_26886_ _33872_/Q _23481_/X _26888_/S VGND VGND VPWR VPWR _26887_/A sky130_fd_sc_hd__mux2_1
XFILLER_208_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28625_ _28625_/A VGND VGND VPWR VPWR _34633_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25837_ _24834_/X _33377_/Q _25853_/S VGND VGND VPWR VPWR _25838_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28556_ _27701_/X _34601_/Q _28556_/S VGND VGND VPWR VPWR _28557_/A sky130_fd_sc_hd__mux2_1
X_16570_ _17982_/A VGND VGND VPWR VPWR _16570_/X sky130_fd_sc_hd__buf_6
X_25768_ _25768_/A VGND VGND VPWR VPWR _33344_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_216_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27507_ _27507_/A VGND VGND VPWR VPWR _34134_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24719_ _22971_/X _32881_/Q _24723_/S VGND VGND VPWR VPWR _24720_/A sky130_fd_sc_hd__mux2_1
X_28487_ _27797_/X _34568_/Q _28505_/S VGND VGND VPWR VPWR _28488_/A sky130_fd_sc_hd__mux2_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25699_ _25810_/S VGND VGND VPWR VPWR _25718_/S sky130_fd_sc_hd__buf_4
XFILLER_187_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18240_ _34708_/Q _34644_/Q _34580_/Q _34516_/Q _17998_/X _17999_/X VGND VGND VPWR
+ VPWR _18240_/X sky130_fd_sc_hd__mux4_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27438_ _34102_/Q _27134_/X _27452_/S VGND VGND VPWR VPWR _27439_/A sky130_fd_sc_hd__mux2_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18171_ _17158_/A _18169_/X _18170_/X _17163_/A VGND VGND VPWR VPWR _18171_/X sky130_fd_sc_hd__a22o_1
X_27369_ _29662_/B _31688_/B VGND VGND VPWR VPWR _27502_/S sky130_fd_sc_hd__nor2_8
XFILLER_156_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1066 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29108_ _34861_/Q _27106_/X _29120_/S VGND VGND VPWR VPWR _29109_/A sky130_fd_sc_hd__mux2_1
X_17122_ _17122_/A _17122_/B _17122_/C _17122_/D VGND VGND VPWR VPWR _17123_/A sky130_fd_sc_hd__or4_4
XFILLER_7_532 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30380_ _30470_/S VGND VGND VPWR VPWR _30399_/S sky130_fd_sc_hd__buf_6
XFILLER_89_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17053_ _34162_/Q _34098_/Q _34034_/Q _33970_/Q _16740_/X _16741_/X VGND VGND VPWR
+ VPWR _17053_/X sky130_fd_sc_hd__mux4_1
XFILLER_13_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29039_ _29039_/A VGND VGND VPWR VPWR _34828_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_221_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1020 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_43_CLK clkbuf_6_6__f_CLK/X VGND VGND VPWR VPWR _35812_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_183_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16004_ _33366_/Q _33302_/Q _33238_/Q _33174_/Q _16002_/X _16003_/X VGND VGND VPWR
+ VPWR _16004_/X sky130_fd_sc_hd__mux4_1
XFILLER_137_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32050_ _35187_/CLK _32050_/D VGND VGND VPWR VPWR _32050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31001_ _31001_/A VGND VGND VPWR VPWR _35728_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_912 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17955_ _17773_/X _17953_/X _17954_/X _17777_/X VGND VGND VPWR VPWR _17955_/X sky130_fd_sc_hd__a22o_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1015 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35740_ _35804_/CLK _35740_/D VGND VGND VPWR VPWR _35740_/Q sky130_fd_sc_hd__dfxtp_1
X_16906_ _16900_/X _16905_/X _16798_/X VGND VGND VPWR VPWR _16914_/C sky130_fd_sc_hd__o21ba_1
X_32952_ _36024_/CLK _32952_/D VGND VGND VPWR VPWR _32952_/Q sky130_fd_sc_hd__dfxtp_1
X_17886_ _32905_/Q _32841_/Q _32777_/Q _32713_/Q _17699_/X _17700_/X VGND VGND VPWR
+ VPWR _17886_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19625_ _19621_/X _19624_/X _19451_/X VGND VGND VPWR VPWR _19633_/C sky130_fd_sc_hd__o21ba_1
X_31903_ _31903_/A VGND VGND VPWR VPWR _36155_/D sky130_fd_sc_hd__clkbuf_1
X_35671_ _35735_/CLK _35671_/D VGND VGND VPWR VPWR _35671_/Q sky130_fd_sc_hd__dfxtp_1
X_16837_ _34667_/Q _34603_/Q _34539_/Q _34475_/Q _16586_/X _16587_/X VGND VGND VPWR
+ VPWR _16837_/X sky130_fd_sc_hd__mux4_1
XFILLER_19_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32883_ _32904_/CLK _32883_/D VGND VGND VPWR VPWR _32883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34622_ _36103_/CLK _34622_/D VGND VGND VPWR VPWR _34622_/Q sky130_fd_sc_hd__dfxtp_1
X_31834_ _31834_/A VGND VGND VPWR VPWR _36122_/D sky130_fd_sc_hd__clkbuf_1
X_19556_ _35447_/Q _35383_/Q _35319_/Q _35255_/Q _19554_/X _19555_/X VGND VGND VPWR
+ VPWR _19556_/X sky130_fd_sc_hd__mux4_1
XFILLER_47_992 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_22_0_CLK clkbuf_2_2_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_22_0_CLK/X sky130_fd_sc_hd__clkbuf_8
X_16768_ _16764_/X _16767_/X _16459_/X VGND VGND VPWR VPWR _16769_/D sky130_fd_sc_hd__o21ba_1
XFILLER_207_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18507_ _18503_/X _18506_/X _18404_/X VGND VGND VPWR VPWR _18508_/D sky130_fd_sc_hd__o21ba_1
XFILLER_34_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34553_ _36152_/CLK _34553_/D VGND VGND VPWR VPWR _34553_/Q sky130_fd_sc_hd__dfxtp_1
X_31765_ _36090_/Q input30/X _31771_/S VGND VGND VPWR VPWR _31766_/A sky130_fd_sc_hd__mux2_1
X_19487_ _33077_/Q _32053_/Q _35829_/Q _35765_/Q _19378_/X _19379_/X VGND VGND VPWR
+ VPWR _19487_/X sky130_fd_sc_hd__mux4_1
X_16699_ _33640_/Q _33576_/Q _33512_/Q _33448_/Q _16494_/X _16495_/X VGND VGND VPWR
+ VPWR _16699_/X sky130_fd_sc_hd__mux4_1
XFILLER_59_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33504_ _36202_/CLK _33504_/D VGND VGND VPWR VPWR _33504_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18438_ _18438_/A _18438_/B _18438_/C _18438_/D VGND VGND VPWR VPWR _18439_/A sky130_fd_sc_hd__or4_2
X_30716_ _35593_/Q _29488_/X _30732_/S VGND VGND VPWR VPWR _30717_/A sky130_fd_sc_hd__mux2_1
X_34484_ _34612_/CLK _34484_/D VGND VGND VPWR VPWR _34484_/Q sky130_fd_sc_hd__dfxtp_1
X_31696_ _36057_/Q input34/X _31708_/S VGND VGND VPWR VPWR _31697_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36223_ _36223_/CLK _36223_/D VGND VGND VPWR VPWR _36223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33435_ _33753_/CLK _33435_/D VGND VGND VPWR VPWR _33435_/Q sky130_fd_sc_hd__dfxtp_1
X_18369_ _20236_/A VGND VGND VPWR VPWR _18369_/X sky130_fd_sc_hd__buf_4
X_30647_ _30647_/A VGND VGND VPWR VPWR _35560_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20400_ _34192_/Q _34128_/Q _34064_/Q _34000_/Q _20099_/X _20100_/X VGND VGND VPWR
+ VPWR _20400_/X sky130_fd_sc_hd__mux4_1
XFILLER_159_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36154_ _36154_/CLK _36154_/D VGND VGND VPWR VPWR _36154_/Q sky130_fd_sc_hd__dfxtp_1
X_33366_ _35804_/CLK _33366_/D VGND VGND VPWR VPWR _33366_/Q sky130_fd_sc_hd__dfxtp_1
X_21380_ _21373_/X _21378_/X _21379_/X VGND VGND VPWR VPWR _21414_/A sky130_fd_sc_hd__o21ba_1
X_30578_ _30605_/S VGND VGND VPWR VPWR _30597_/S sky130_fd_sc_hd__buf_4
XFILLER_120_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35105_ _35168_/CLK _35105_/D VGND VGND VPWR VPWR _35105_/Q sky130_fd_sc_hd__dfxtp_1
X_20331_ _35213_/Q _35149_/Q _35085_/Q _32269_/Q _20016_/X _20017_/X VGND VGND VPWR
+ VPWR _20331_/X sky130_fd_sc_hd__mux4_1
XFILLER_175_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32317_ _32575_/CLK _32317_/D VGND VGND VPWR VPWR _32317_/Q sky130_fd_sc_hd__dfxtp_1
X_36085_ _36085_/CLK _36085_/D VGND VGND VPWR VPWR _36085_/Q sky130_fd_sc_hd__dfxtp_1
X_33297_ _36106_/CLK _33297_/D VGND VGND VPWR VPWR _33297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_34_CLK clkbuf_6_7__f_CLK/X VGND VGND VPWR VPWR _36005_/CLK sky130_fd_sc_hd__clkbuf_16
X_35036_ _36219_/CLK _35036_/D VGND VGND VPWR VPWR _35036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23050_ _23049_/X _32074_/Q _23071_/S VGND VGND VPWR VPWR _23051_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20262_ _35467_/Q _35403_/Q _35339_/Q _35275_/Q _20260_/X _20261_/X VGND VGND VPWR
+ VPWR _20262_/X sky130_fd_sc_hd__mux4_1
XFILLER_150_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32248_ _36150_/CLK _32248_/D VGND VGND VPWR VPWR _32248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22001_ _21758_/X _21999_/X _22000_/X _21763_/X VGND VGND VPWR VPWR _22001_/X sky130_fd_sc_hd__a22o_1
XTAP_6009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20193_ _33097_/Q _32073_/Q _35849_/Q _35785_/Q _20084_/X _20085_/X VGND VGND VPWR
+ VPWR _20193_/X sky130_fd_sc_hd__mux4_1
XFILLER_143_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32179_ _35482_/CLK _32179_/D VGND VGND VPWR VPWR _32179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26740_ _26740_/A VGND VGND VPWR VPWR _33802_/D sky130_fd_sc_hd__clkbuf_1
X_23952_ _23952_/A VGND VGND VPWR VPWR _32520_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_233_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35938_ _35938_/CLK _35938_/D VGND VGND VPWR VPWR _35938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_244_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22903_ input56/X VGND VGND VPWR VPWR _22903_/X sky130_fd_sc_hd__buf_2
XTAP_3917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26671_ _26761_/S VGND VGND VPWR VPWR _26690_/S sky130_fd_sc_hd__buf_4
XFILLER_84_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35869_ _35997_/CLK _35869_/D VGND VGND VPWR VPWR _35869_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23883_ _22943_/X _32488_/Q _23885_/S VGND VGND VPWR VPWR _23884_/A sky130_fd_sc_hd__mux2_1
XFILLER_217_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28410_ _28410_/A VGND VGND VPWR VPWR _34531_/D sky130_fd_sc_hd__clkbuf_1
X_22834_ _35668_/Q _35028_/Q _34388_/Q _33748_/Q _20712_/X _20713_/X VGND VGND VPWR
+ VPWR _22834_/X sky130_fd_sc_hd__mux4_1
X_25622_ _25622_/A VGND VGND VPWR VPWR _33275_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29390_ _29390_/A VGND VGND VPWR VPWR _34985_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28341_ _27782_/X _34499_/Q _28349_/S VGND VGND VPWR VPWR _28342_/A sky130_fd_sc_hd__mux2_1
X_25553_ _25553_/A VGND VGND VPWR VPWR _33242_/D sky130_fd_sc_hd__clkbuf_1
X_22765_ _22761_/X _22764_/X _22438_/A VGND VGND VPWR VPWR _22787_/A sky130_fd_sc_hd__o21ba_1
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24504_ _23052_/X _32779_/Q _24516_/S VGND VGND VPWR VPWR _24505_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_826 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21716_ _35187_/Q _35123_/Q _35059_/Q _32220_/Q _21610_/X _21611_/X VGND VGND VPWR
+ VPWR _21716_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28272_ _27680_/X _34466_/Q _28286_/S VGND VGND VPWR VPWR _28273_/A sky130_fd_sc_hd__mux2_1
XFILLER_212_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25484_ _24911_/X _33210_/Q _25490_/S VGND VGND VPWR VPWR _25485_/A sky130_fd_sc_hd__mux2_1
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22696_ _22692_/X _22695_/X _22471_/X VGND VGND VPWR VPWR _22697_/D sky130_fd_sc_hd__o21ba_1
XFILLER_169_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1099 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27223_ input58/X VGND VGND VPWR VPWR _27223_/X sky130_fd_sc_hd__clkbuf_4
X_24435_ _22949_/X _32746_/Q _24453_/S VGND VGND VPWR VPWR _24436_/A sky130_fd_sc_hd__mux2_1
X_21647_ _34929_/Q _34865_/Q _34801_/Q _34737_/Q _21407_/X _21408_/X VGND VGND VPWR
+ VPWR _21647_/X sky130_fd_sc_hd__mux4_1
XFILLER_197_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27154_ _27154_/A VGND VGND VPWR VPWR _33980_/D sky130_fd_sc_hd__clkbuf_1
X_24366_ _24366_/A VGND VGND VPWR VPWR _32713_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21578_ _21405_/X _21576_/X _21577_/X _21410_/X VGND VGND VPWR VPWR _21578_/X sky130_fd_sc_hd__a22o_1
XFILLER_240_1299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26105_ _24830_/X _33504_/Q _26123_/S VGND VGND VPWR VPWR _26106_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23317_ _32176_/Q _23316_/X _23424_/S VGND VGND VPWR VPWR _23318_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20529_ _32148_/Q _32340_/Q _32404_/Q _35924_/Q _20286_/X _19311_/A VGND VGND VPWR
+ VPWR _20529_/X sky130_fd_sc_hd__mux4_1
X_27085_ _33958_/Q _27084_/X _27094_/S VGND VGND VPWR VPWR _27086_/A sky130_fd_sc_hd__mux2_1
X_24297_ _22946_/X _32681_/Q _24297_/S VGND VGND VPWR VPWR _24298_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_25_CLK clkbuf_6_4__f_CLK/X VGND VGND VPWR VPWR _35168_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_193_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26036_ _26036_/A VGND VGND VPWR VPWR _33471_/D sky130_fd_sc_hd__clkbuf_1
X_23248_ _23248_/A VGND VGND VPWR VPWR _32155_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23179_ _23179_/A VGND VGND VPWR VPWR _32127_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27987_ _34331_/Q _27050_/X _27995_/S VGND VGND VPWR VPWR _27988_/A sky130_fd_sc_hd__mux2_1
XTAP_6576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17740_ _17420_/X _17738_/X _17739_/X _17424_/X VGND VGND VPWR VPWR _17740_/X sky130_fd_sc_hd__a22o_1
X_29726_ _29795_/S VGND VGND VPWR VPWR _29745_/S sky130_fd_sc_hd__buf_6
XTAP_6598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26938_ _26938_/A VGND VGND VPWR VPWR _33896_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_12__f_CLK clkbuf_5_6_0_CLK/X VGND VGND VPWR VPWR clkbuf_leaf_49_CLK/A sky130_fd_sc_hd__clkbuf_16
XFILLER_248_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29657_ _29657_/A VGND VGND VPWR VPWR _35091_/D sky130_fd_sc_hd__clkbuf_1
X_17671_ _17800_/A VGND VGND VPWR VPWR _17671_/X sky130_fd_sc_hd__clkbuf_4
X_26869_ _26896_/S VGND VGND VPWR VPWR _26888_/S sky130_fd_sc_hd__buf_4
XFILLER_235_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19410_ _19298_/X _19408_/X _19409_/X _19301_/X VGND VGND VPWR VPWR _19410_/X sky130_fd_sc_hd__a22o_1
XFILLER_78_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28608_ _28608_/A VGND VGND VPWR VPWR _34625_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16622_ _16447_/X _16620_/X _16621_/X _16450_/X VGND VGND VPWR VPWR _16622_/X sky130_fd_sc_hd__a22o_1
XFILLER_112_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29588_ _29588_/A VGND VGND VPWR VPWR _35058_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19341_ _19303_/X _19339_/X _19340_/X _19306_/X VGND VGND VPWR VPWR _19341_/X sky130_fd_sc_hd__a22o_1
XFILLER_56_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16553_ _16547_/X _16552_/X _16445_/X VGND VGND VPWR VPWR _16561_/C sky130_fd_sc_hd__o21ba_1
X_28539_ _28539_/A VGND VGND VPWR VPWR _34592_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_245_1144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31550_ _31550_/A VGND VGND VPWR VPWR _35988_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19272_ _19268_/X _19271_/X _19098_/X VGND VGND VPWR VPWR _19280_/C sky130_fd_sc_hd__o21ba_1
XFILLER_245_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16484_ _34657_/Q _34593_/Q _34529_/Q _34465_/Q _16233_/X _16234_/X VGND VGND VPWR
+ VPWR _16484_/X sky130_fd_sc_hd__mux4_1
XFILLER_231_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18223_ _33940_/Q _33876_/Q _33812_/Q _36116_/Q _16062_/X _16064_/X VGND VGND VPWR
+ VPWR _18223_/X sky130_fd_sc_hd__mux4_1
XFILLER_62_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30501_ _35491_/Q _29370_/X _30513_/S VGND VGND VPWR VPWR _30502_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_223_1442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31481_ _31481_/A VGND VGND VPWR VPWR _35955_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_248_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33220_ _33415_/CLK _33220_/D VGND VGND VPWR VPWR _33220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18154_ _34961_/Q _34897_/Q _34833_/Q _34769_/Q _17866_/X _17867_/X VGND VGND VPWR
+ VPWR _18154_/X sky130_fd_sc_hd__mux4_1
X_30432_ _30432_/A VGND VGND VPWR VPWR _35458_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17105_ _32883_/Q _32819_/Q _32755_/Q _32691_/Q _16993_/X _16994_/X VGND VGND VPWR
+ VPWR _17105_/X sky130_fd_sc_hd__mux4_1
XFILLER_184_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33151_ _35903_/CLK _33151_/D VGND VGND VPWR VPWR _33151_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18085_ _15981_/X _18083_/X _18084_/X _15991_/X VGND VGND VPWR VPWR _18085_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30363_ _30363_/A VGND VGND VPWR VPWR _35425_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_16_CLK clkbuf_6_6__f_CLK/X VGND VGND VPWR VPWR _36135_/CLK sky130_fd_sc_hd__clkbuf_16
X_32102_ _32552_/CLK _32102_/D VGND VGND VPWR VPWR _32102_/Q sky130_fd_sc_hd__dfxtp_1
X_17036_ _35697_/Q _32205_/Q _35569_/Q _35505_/Q _16964_/X _16965_/X VGND VGND VPWR
+ VPWR _17036_/X sky130_fd_sc_hd__mux4_1
X_30294_ _35393_/Q _29463_/X _30306_/S VGND VGND VPWR VPWR _30295_/A sky130_fd_sc_hd__mux2_1
X_33082_ _36026_/CLK _33082_/D VGND VGND VPWR VPWR _33082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32033_ _35943_/CLK _32033_/D VGND VGND VPWR VPWR _32033_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18987_ _33063_/Q _32039_/Q _35815_/Q _35751_/Q _18672_/X _18673_/X VGND VGND VPWR
+ VPWR _18987_/X sky130_fd_sc_hd__mux4_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17938_ _34954_/Q _34890_/Q _34826_/Q _34762_/Q _17866_/X _17867_/X VGND VGND VPWR
+ VPWR _17938_/X sky130_fd_sc_hd__mux4_1
XFILLER_230_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33984_ _33984_/CLK _33984_/D VGND VGND VPWR VPWR _33984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35723_ _35723_/CLK _35723_/D VGND VGND VPWR VPWR _35723_/Q sky130_fd_sc_hd__dfxtp_1
X_32935_ _36007_/CLK _32935_/D VGND VGND VPWR VPWR _32935_/Q sky130_fd_sc_hd__dfxtp_1
X_17869_ _17869_/A VGND VGND VPWR VPWR _17869_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_22_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19608_ _19506_/X _19606_/X _19607_/X _19509_/X VGND VGND VPWR VPWR _19608_/X sky130_fd_sc_hd__a22o_1
X_35654_ _35655_/CLK _35654_/D VGND VGND VPWR VPWR _35654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20880_ _33884_/Q _33820_/Q _33756_/Q _36060_/Q _20712_/X _20713_/X VGND VGND VPWR
+ VPWR _20880_/X sky130_fd_sc_hd__mux4_1
X_32866_ _32869_/CLK _32866_/D VGND VGND VPWR VPWR _32866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34605_ _35181_/CLK _34605_/D VGND VGND VPWR VPWR _34605_/Q sky130_fd_sc_hd__dfxtp_1
X_31817_ _36115_/Q input58/X _31821_/S VGND VGND VPWR VPWR _31818_/A sky130_fd_sc_hd__mux2_1
X_19539_ _19499_/X _19537_/X _19538_/X _19504_/X VGND VGND VPWR VPWR _19539_/X sky130_fd_sc_hd__a22o_1
XFILLER_241_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35585_ _35646_/CLK _35585_/D VGND VGND VPWR VPWR _35585_/Q sky130_fd_sc_hd__dfxtp_1
X_32797_ _32797_/CLK _32797_/D VGND VGND VPWR VPWR _32797_/Q sky130_fd_sc_hd__dfxtp_1
X_22550_ _32651_/Q _32587_/Q _32523_/Q _35979_/Q _22229_/X _22366_/X VGND VGND VPWR
+ VPWR _22550_/X sky130_fd_sc_hd__mux4_1
X_34536_ _35684_/CLK _34536_/D VGND VGND VPWR VPWR _34536_/Q sky130_fd_sc_hd__dfxtp_1
X_31748_ _36082_/Q input21/X _31750_/S VGND VGND VPWR VPWR _31749_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21501_ _22560_/A VGND VGND VPWR VPWR _21501_/X sky130_fd_sc_hd__buf_4
XFILLER_50_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22481_ _22477_/X _22480_/X _22438_/X VGND VGND VPWR VPWR _22503_/A sky130_fd_sc_hd__o21ba_1
XFILLER_179_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34467_ _36209_/CLK _34467_/D VGND VGND VPWR VPWR _34467_/Q sky130_fd_sc_hd__dfxtp_1
X_31679_ _31679_/A VGND VGND VPWR VPWR _36049_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_829 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36206_ _36211_/CLK _36206_/D VGND VGND VPWR VPWR _36206_/Q sky130_fd_sc_hd__dfxtp_1
X_24220_ _32646_/Q _23447_/X _24222_/S VGND VGND VPWR VPWR _24221_/A sky130_fd_sc_hd__mux2_1
X_33418_ _33673_/CLK _33418_/D VGND VGND VPWR VPWR _33418_/Q sky130_fd_sc_hd__dfxtp_1
X_21432_ _21245_/X _21430_/X _21431_/X _21248_/X VGND VGND VPWR VPWR _21432_/X sky130_fd_sc_hd__a22o_1
XFILLER_194_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34398_ _36235_/CLK _34398_/D VGND VGND VPWR VPWR _34398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36137_ _36137_/CLK _36137_/D VGND VGND VPWR VPWR _36137_/Q sky130_fd_sc_hd__dfxtp_1
X_24151_ _32613_/Q _23277_/X _24159_/S VGND VGND VPWR VPWR _24152_/A sky130_fd_sc_hd__mux2_1
X_33349_ _34177_/CLK _33349_/D VGND VGND VPWR VPWR _33349_/Q sky130_fd_sc_hd__dfxtp_1
X_21363_ _35177_/Q _35113_/Q _35049_/Q _32169_/Q _21257_/X _21258_/X VGND VGND VPWR
+ VPWR _21363_/X sky130_fd_sc_hd__mux4_1
XFILLER_238_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23102_ _22903_/X _32091_/Q _23110_/S VGND VGND VPWR VPWR _23103_/A sky130_fd_sc_hd__mux2_1
X_20314_ _20212_/X _20312_/X _20313_/X _20215_/X VGND VGND VPWR VPWR _20314_/X sky130_fd_sc_hd__a22o_1
X_24082_ _23036_/X _32582_/Q _24084_/S VGND VGND VPWR VPWR _24083_/A sky130_fd_sc_hd__mux2_1
X_36068_ _36068_/CLK _36068_/D VGND VGND VPWR VPWR _36068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21294_ _34919_/Q _34855_/Q _34791_/Q _34727_/Q _21054_/X _21055_/X VGND VGND VPWR
+ VPWR _21294_/X sky130_fd_sc_hd__mux4_1
XFILLER_163_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35019_ _35724_/CLK _35019_/D VGND VGND VPWR VPWR _35019_/Q sky130_fd_sc_hd__dfxtp_1
X_23033_ input42/X VGND VGND VPWR VPWR _23033_/X sky130_fd_sc_hd__buf_2
X_27910_ _27910_/A VGND VGND VPWR VPWR _34294_/D sky130_fd_sc_hd__clkbuf_1
X_20245_ _20205_/X _20243_/X _20244_/X _20210_/X VGND VGND VPWR VPWR _20245_/X sky130_fd_sc_hd__a22o_1
XFILLER_235_1324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28890_ _34758_/Q _27183_/X _28892_/S VGND VGND VPWR VPWR _28891_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27841_ _27973_/S VGND VGND VPWR VPWR _27860_/S sky130_fd_sc_hd__buf_4
XTAP_5105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20176_ _34185_/Q _34121_/Q _34057_/Q _33993_/Q _20099_/X _20100_/X VGND VGND VPWR
+ VPWR _20176_/X sky130_fd_sc_hd__mux4_1
XTAP_5116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27772_ _27772_/A VGND VGND VPWR VPWR _34239_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_1109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24984_ _24984_/A VGND VGND VPWR VPWR _32977_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29511_ _29511_/A VGND VGND VPWR VPWR _35024_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26723_ _26723_/A VGND VGND VPWR VPWR _33794_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23935_ _23935_/A VGND VGND VPWR VPWR _32512_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29442_ _35002_/Q _29441_/X _29451_/S VGND VGND VPWR VPWR _29443_/A sky130_fd_sc_hd__mux2_1
XFILLER_244_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26654_ _26654_/A VGND VGND VPWR VPWR _33761_/D sky130_fd_sc_hd__clkbuf_1
X_23866_ _23977_/S VGND VGND VPWR VPWR _23885_/S sky130_fd_sc_hd__buf_4
XTAP_3769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22817_ _22817_/A _22817_/B _22817_/C _22817_/D VGND VGND VPWR VPWR _22818_/A sky130_fd_sc_hd__or4_4
X_25605_ _25605_/A VGND VGND VPWR VPWR _33267_/D sky130_fd_sc_hd__clkbuf_1
X_29373_ input6/X VGND VGND VPWR VPWR _29373_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_72_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26585_ _24939_/X _33731_/Q _26593_/S VGND VGND VPWR VPWR _26586_/A sky130_fd_sc_hd__mux2_1
X_23797_ _23018_/X _32384_/Q _23811_/S VGND VGND VPWR VPWR _23798_/A sky130_fd_sc_hd__mux2_1
XFILLER_246_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28324_ _27757_/X _34491_/Q _28328_/S VGND VGND VPWR VPWR _28325_/A sky130_fd_sc_hd__mux2_1
X_25536_ _24988_/X _33235_/Q _25540_/S VGND VGND VPWR VPWR _25537_/A sky130_fd_sc_hd__mux2_1
X_22748_ _20601_/X _22746_/X _22747_/X _20607_/X VGND VGND VPWR VPWR _22748_/X sky130_fd_sc_hd__a22o_1
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28255_ _27655_/X _34458_/Q _28265_/S VGND VGND VPWR VPWR _28256_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25467_ _24886_/X _33202_/Q _25469_/S VGND VGND VPWR VPWR _25468_/A sky130_fd_sc_hd__mux2_1
X_22679_ _32143_/Q _32335_/Q _32399_/Q _35919_/Q _22586_/X _22374_/X VGND VGND VPWR
+ VPWR _22679_/X sky130_fd_sc_hd__mux4_1
XFILLER_197_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27206_ _33997_/Q _27205_/X _27218_/S VGND VGND VPWR VPWR _27207_/A sky130_fd_sc_hd__mux2_1
X_24418_ _22925_/X _32738_/Q _24432_/S VGND VGND VPWR VPWR _24419_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25398_ _25398_/A VGND VGND VPWR VPWR _33170_/D sky130_fd_sc_hd__clkbuf_1
X_28186_ _28186_/A VGND VGND VPWR VPWR _34425_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24349_ _24349_/A VGND VGND VPWR VPWR _32705_/D sky130_fd_sc_hd__clkbuf_1
X_27137_ input27/X VGND VGND VPWR VPWR _27137_/X sky130_fd_sc_hd__buf_2
XFILLER_103_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27068_ _27068_/A VGND VGND VPWR VPWR _33952_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26019_ _26019_/A VGND VGND VPWR VPWR _33463_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18910_ _18906_/X _18909_/X _18734_/X _18735_/X VGND VGND VPWR VPWR _18927_/B sky130_fd_sc_hd__o211a_1
XTAP_7030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19890_ _33665_/Q _33601_/Q _33537_/Q _33473_/Q _19853_/X _19854_/X VGND VGND VPWR
+ VPWR _19890_/X sky130_fd_sc_hd__mux4_1
XFILLER_175_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18841_ _32099_/Q _32291_/Q _32355_/Q _35875_/Q _18521_/X _18662_/X VGND VGND VPWR
+ VPWR _18841_/X sky130_fd_sc_hd__mux4_1
XTAP_7085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18772_ _18653_/X _18770_/X _18771_/X _18659_/X VGND VGND VPWR VPWR _18772_/X sky130_fd_sc_hd__a22o_1
XTAP_6395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15984_ _17906_/A VGND VGND VPWR VPWR _15984_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_48_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17723_ _17719_/X _17722_/X _17518_/X VGND VGND VPWR VPWR _17724_/D sky130_fd_sc_hd__o21ba_1
X_29709_ _29709_/A VGND VGND VPWR VPWR _35115_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30981_ _35719_/Q input44/X _30981_/S VGND VGND VPWR VPWR _30982_/A sky130_fd_sc_hd__mux2_1
XTAP_4960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32720_ _32914_/CLK _32720_/D VGND VGND VPWR VPWR _32720_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17654_ _17654_/A _17654_/B _17654_/C _17654_/D VGND VGND VPWR VPWR _17655_/A sky130_fd_sc_hd__or4_2
XFILLER_75_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_5_CLK clkbuf_leaf_9_CLK/A VGND VGND VPWR VPWR _34918_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_91_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16605_ _33125_/Q _36005_/Q _32997_/Q _32933_/Q _16356_/X _16357_/X VGND VGND VPWR
+ VPWR _16605_/X sky130_fd_sc_hd__mux4_1
XFILLER_223_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32651_ _36044_/CLK _32651_/D VGND VGND VPWR VPWR _32651_/Q sky130_fd_sc_hd__dfxtp_1
X_17585_ _34944_/Q _34880_/Q _34816_/Q _34752_/Q _17513_/X _17514_/X VGND VGND VPWR
+ VPWR _17585_/X sky130_fd_sc_hd__mux4_1
XFILLER_189_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19324_ _20150_/A VGND VGND VPWR VPWR _19324_/X sky130_fd_sc_hd__buf_4
X_31602_ _31602_/A VGND VGND VPWR VPWR _36012_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16536_ _16500_/X _16534_/X _16535_/X _16503_/X VGND VGND VPWR VPWR _16536_/X sky130_fd_sc_hd__a22o_1
X_35370_ _35685_/CLK _35370_/D VGND VGND VPWR VPWR _35370_/Q sky130_fd_sc_hd__dfxtp_1
X_32582_ _35974_/CLK _32582_/D VGND VGND VPWR VPWR _32582_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_232_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34321_ _36177_/CLK _34321_/D VGND VGND VPWR VPWR _34321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31533_ _27810_/X _35980_/Q _31543_/S VGND VGND VPWR VPWR _31534_/A sky130_fd_sc_hd__mux2_1
X_19255_ _19153_/X _19253_/X _19254_/X _19156_/X VGND VGND VPWR VPWR _19255_/X sky130_fd_sc_hd__a22o_1
XFILLER_31_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16467_ _33889_/Q _33825_/Q _33761_/Q _36065_/Q _16318_/X _16319_/X VGND VGND VPWR
+ VPWR _16467_/X sky130_fd_sc_hd__mux4_1
XFILLER_176_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18206_ _35475_/Q _35411_/Q _35347_/Q _35283_/Q _17960_/X _17961_/X VGND VGND VPWR
+ VPWR _18206_/X sky130_fd_sc_hd__mux4_1
X_34252_ _36173_/CLK _34252_/D VGND VGND VPWR VPWR _34252_/Q sky130_fd_sc_hd__dfxtp_1
X_19186_ _19146_/X _19184_/X _19185_/X _19151_/X VGND VGND VPWR VPWR _19186_/X sky130_fd_sc_hd__a22o_1
X_31464_ _27708_/X _35947_/Q _31480_/S VGND VGND VPWR VPWR _31465_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16398_ _32095_/Q _32287_/Q _32351_/Q _35871_/Q _16221_/X _16362_/X VGND VGND VPWR
+ VPWR _16398_/X sky130_fd_sc_hd__mux4_1
XFILLER_106_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_970 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33203_ _33393_/CLK _33203_/D VGND VGND VPWR VPWR _33203_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18137_ _33169_/Q _36049_/Q _33041_/Q _32977_/Q _16032_/X _17161_/A VGND VGND VPWR
+ VPWR _18137_/X sky130_fd_sc_hd__mux4_1
XFILLER_129_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30415_ _30415_/A VGND VGND VPWR VPWR _35450_/D sky130_fd_sc_hd__clkbuf_1
X_34183_ _34183_/CLK _34183_/D VGND VGND VPWR VPWR _34183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31395_ _31395_/A VGND VGND VPWR VPWR _35914_/D sky130_fd_sc_hd__clkbuf_1
X_33134_ _36015_/CLK _33134_/D VGND VGND VPWR VPWR _33134_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30346_ _30346_/A VGND VGND VPWR VPWR _35417_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_176_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18068_ _18068_/A VGND VGND VPWR VPWR _32014_/D sky130_fd_sc_hd__buf_2
X_17019_ _17019_/A VGND VGND VPWR VPWR _31984_/D sky130_fd_sc_hd__clkbuf_1
X_33065_ _35755_/CLK _33065_/D VGND VGND VPWR VPWR _33065_/Q sky130_fd_sc_hd__dfxtp_1
X_30277_ _35385_/Q _29438_/X _30285_/S VGND VGND VPWR VPWR _30278_/A sky130_fd_sc_hd__mux2_1
X_20030_ _20150_/A VGND VGND VPWR VPWR _20030_/X sky130_fd_sc_hd__buf_4
X_32016_ _36202_/CLK _32016_/D VGND VGND VPWR VPWR _32016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_246_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33967_ _34991_/CLK _33967_/D VGND VGND VPWR VPWR _33967_/Q sky130_fd_sc_hd__dfxtp_1
X_21981_ _21975_/X _21980_/X _21732_/X VGND VGND VPWR VPWR _22003_/A sky130_fd_sc_hd__o21ba_1
XFILLER_67_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23720_ _23720_/A VGND VGND VPWR VPWR _32347_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32918_ _35863_/CLK _32918_/D VGND VGND VPWR VPWR _32918_/Q sky130_fd_sc_hd__dfxtp_1
X_20932_ _20892_/X _20930_/X _20931_/X _20895_/X VGND VGND VPWR VPWR _20932_/X sky130_fd_sc_hd__a22o_1
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35706_ _35709_/CLK _35706_/D VGND VGND VPWR VPWR _35706_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33898_ _34091_/CLK _33898_/D VGND VGND VPWR VPWR _33898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23651_ _23651_/A VGND VGND VPWR VPWR _32316_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_226_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20863_ _35419_/Q _35355_/Q _35291_/Q _35227_/Q _20795_/X _20796_/X VGND VGND VPWR
+ VPWR _20863_/X sky130_fd_sc_hd__mux4_1
X_32849_ _32913_/CLK _32849_/D VGND VGND VPWR VPWR _32849_/Q sky130_fd_sc_hd__dfxtp_1
X_35637_ _35701_/CLK _35637_/D VGND VGND VPWR VPWR _35637_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22602_ _22459_/X _22600_/X _22601_/X _22462_/X VGND VGND VPWR VPWR _22602_/X sky130_fd_sc_hd__a22o_1
XFILLER_228_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26370_ _26370_/A VGND VGND VPWR VPWR _33629_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23582_ _23582_/A VGND VGND VPWR VPWR _32283_/D sky130_fd_sc_hd__clkbuf_1
X_35568_ _35635_/CLK _35568_/D VGND VGND VPWR VPWR _35568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20794_ _20648_/X _20792_/X _20793_/X _20658_/X VGND VGND VPWR VPWR _20794_/X sky130_fd_sc_hd__a22o_1
XFILLER_165_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25321_ _25321_/A VGND VGND VPWR VPWR _33133_/D sky130_fd_sc_hd__clkbuf_1
X_34519_ _34903_/CLK _34519_/D VGND VGND VPWR VPWR _34519_/Q sky130_fd_sc_hd__dfxtp_1
X_22533_ _35210_/Q _35146_/Q _35082_/Q _32266_/Q _22316_/X _22317_/X VGND VGND VPWR
+ VPWR _22533_/X sky130_fd_sc_hd__mux4_1
X_35499_ _35691_/CLK _35499_/D VGND VGND VPWR VPWR _35499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25252_ _25252_/A VGND VGND VPWR VPWR _33101_/D sky130_fd_sc_hd__clkbuf_1
X_28040_ _34356_/Q _27127_/X _28058_/S VGND VGND VPWR VPWR _28041_/A sky130_fd_sc_hd__mux2_1
X_22464_ _22464_/A VGND VGND VPWR VPWR _22464_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_155_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24203_ _24251_/S VGND VGND VPWR VPWR _24222_/S sky130_fd_sc_hd__buf_4
XFILLER_185_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21415_ _21415_/A VGND VGND VPWR VPWR _36202_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25183_ _25183_/A VGND VGND VPWR VPWR _33068_/D sky130_fd_sc_hd__clkbuf_1
X_22395_ _22391_/X _22394_/X _22118_/X VGND VGND VPWR VPWR _22396_/D sky130_fd_sc_hd__o21ba_1
XFILLER_175_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_1389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_1282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24134_ _32605_/Q _23252_/X _24138_/S VGND VGND VPWR VPWR _24135_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21346_ _21100_/X _21344_/X _21345_/X _21103_/X VGND VGND VPWR VPWR _21346_/X sky130_fd_sc_hd__a22o_1
XFILLER_163_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29991_ _29991_/A VGND VGND VPWR VPWR _35249_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28942_ _28942_/A VGND VGND VPWR VPWR _34782_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24065_ _24113_/S VGND VGND VPWR VPWR _24084_/S sky130_fd_sc_hd__buf_4
XFILLER_11_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21277_ _33127_/Q _36007_/Q _32999_/Q _32935_/Q _20956_/X _20957_/X VGND VGND VPWR
+ VPWR _21277_/X sky130_fd_sc_hd__mux4_1
X_23016_ _23015_/X _32063_/Q _23040_/S VGND VGND VPWR VPWR _23017_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20228_ _35466_/Q _35402_/Q _35338_/Q _35274_/Q _19907_/X _19908_/X VGND VGND VPWR
+ VPWR _20228_/X sky130_fd_sc_hd__mux4_1
X_28873_ _28921_/S VGND VGND VPWR VPWR _28892_/S sky130_fd_sc_hd__buf_4
XFILLER_131_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_231_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27824_ _27824_/A VGND VGND VPWR VPWR _34256_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_1439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20159_ _20159_/A VGND VGND VPWR VPWR _20159_/X sky130_fd_sc_hd__clkbuf_4
XTAP_4201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27755_ _27754_/X _34234_/Q _27764_/S VGND VGND VPWR VPWR _27756_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24967_ input50/X VGND VGND VPWR VPWR _24967_/X sky130_fd_sc_hd__buf_4
XTAP_4256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26706_ _26706_/A VGND VGND VPWR VPWR _33786_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_246_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23918_ _23918_/A VGND VGND VPWR VPWR _32504_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27686_ input6/X VGND VGND VPWR VPWR _27686_/X sky130_fd_sc_hd__buf_4
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24898_ _24898_/A VGND VGND VPWR VPWR _32949_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29425_ _29425_/A VGND VGND VPWR VPWR _34996_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26637_ _26637_/A VGND VGND VPWR VPWR _33753_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23849_ _23849_/A VGND VGND VPWR VPWR _32471_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29356_ _29356_/A VGND VGND VPWR VPWR _34974_/D sky130_fd_sc_hd__clkbuf_1
X_17370_ _17366_/X _17369_/X _17165_/X VGND VGND VPWR VPWR _17371_/D sky130_fd_sc_hd__o21ba_1
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26568_ _24914_/X _33723_/Q _26572_/S VGND VGND VPWR VPWR _26569_/A sky130_fd_sc_hd__mux2_1
XFILLER_232_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16321_ _16147_/X _16317_/X _16320_/X _16150_/X VGND VGND VPWR VPWR _16321_/X sky130_fd_sc_hd__a22o_1
X_28307_ _27732_/X _34483_/Q _28307_/S VGND VGND VPWR VPWR _28308_/A sky130_fd_sc_hd__mux2_1
XFILLER_242_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25519_ _25519_/A VGND VGND VPWR VPWR _33226_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29287_ _34946_/Q _27171_/X _29297_/S VGND VGND VPWR VPWR _29288_/A sky130_fd_sc_hd__mux2_1
XFILLER_203_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26499_ _24812_/X _33690_/Q _26509_/S VGND VGND VPWR VPWR _26500_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19040_ _20260_/A VGND VGND VPWR VPWR _19040_/X sky130_fd_sc_hd__buf_4
X_28238_ _28238_/A VGND VGND VPWR VPWR _34450_/D sky130_fd_sc_hd__clkbuf_1
X_16252_ _33115_/Q _35995_/Q _32987_/Q _32923_/Q _16024_/X _16025_/X VGND VGND VPWR
+ VPWR _16252_/X sky130_fd_sc_hd__mux4_1
XFILLER_51_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16183_ _16147_/X _16181_/X _16182_/X _16150_/X VGND VGND VPWR VPWR _16183_/X sky130_fd_sc_hd__a22o_1
XFILLER_154_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28169_ _28169_/A VGND VGND VPWR VPWR _34417_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30200_ _35349_/Q _29524_/X _30200_/S VGND VGND VPWR VPWR _30201_/A sky130_fd_sc_hd__mux2_1
Xoutput209 _36187_/Q VGND VGND VPWR VPWR D2[5] sky130_fd_sc_hd__buf_2
X_31180_ _31180_/A VGND VGND VPWR VPWR _35812_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_1328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19942_ _33090_/Q _32066_/Q _35842_/Q _35778_/Q _19731_/X _19732_/X VGND VGND VPWR
+ VPWR _19942_/X sky130_fd_sc_hd__mux4_1
XFILLER_154_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30131_ _30200_/S VGND VGND VPWR VPWR _30150_/S sky130_fd_sc_hd__buf_6
XFILLER_4_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30062_ _30062_/A VGND VGND VPWR VPWR _35283_/D sky130_fd_sc_hd__clkbuf_1
X_19873_ _35648_/Q _35008_/Q _34368_/Q _33728_/Q _19797_/X _19798_/X VGND VGND VPWR
+ VPWR _19873_/X sky130_fd_sc_hd__mux4_1
XFILLER_110_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18824_ _19177_/A VGND VGND VPWR VPWR _18824_/X sky130_fd_sc_hd__buf_4
XFILLER_95_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34870_ _35830_/CLK _34870_/D VGND VGND VPWR VPWR _34870_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33821_ _33821_/CLK _33821_/D VGND VGND VPWR VPWR _33821_/Q sky130_fd_sc_hd__dfxtp_1
X_18755_ _19461_/A VGND VGND VPWR VPWR _18755_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_209_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17706_ _35652_/Q _35012_/Q _34372_/Q _33732_/Q _17497_/X _17498_/X VGND VGND VPWR
+ VPWR _17706_/X sky130_fd_sc_hd__mux4_1
X_33752_ _36057_/CLK _33752_/D VGND VGND VPWR VPWR _33752_/Q sky130_fd_sc_hd__dfxtp_1
X_30964_ _30964_/A VGND VGND VPWR VPWR _35710_/D sky130_fd_sc_hd__clkbuf_1
X_18686_ _33631_/Q _33567_/Q _33503_/Q _33439_/Q _18441_/X _18442_/X VGND VGND VPWR
+ VPWR _18686_/X sky130_fd_sc_hd__mux4_1
XFILLER_97_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32703_ _32894_/CLK _32703_/D VGND VGND VPWR VPWR _32703_/Q sky130_fd_sc_hd__dfxtp_1
X_17637_ _17632_/X _17636_/X _17493_/X _17494_/X VGND VGND VPWR VPWR _17654_/B sky130_fd_sc_hd__o211a_1
XFILLER_247_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33683_ _33875_/CLK _33683_/D VGND VGND VPWR VPWR _33683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30895_ _35678_/Q input63/X _30897_/S VGND VGND VPWR VPWR _30896_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35422_ _35677_/CLK _35422_/D VGND VGND VPWR VPWR _35422_/Q sky130_fd_sc_hd__dfxtp_1
X_32634_ _35451_/CLK _32634_/D VGND VGND VPWR VPWR _32634_/Q sky130_fd_sc_hd__dfxtp_1
X_17568_ _32128_/Q _32320_/Q _32384_/Q _35904_/Q _17280_/X _17421_/X VGND VGND VPWR
+ VPWR _17568_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19307_ _19303_/X _19304_/X _19305_/X _19306_/X VGND VGND VPWR VPWR _19307_/X sky130_fd_sc_hd__a22o_1
XFILLER_232_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35353_ _35674_/CLK _35353_/D VGND VGND VPWR VPWR _35353_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_1072 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1075 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16519_ _16515_/X _16518_/X _16445_/X VGND VGND VPWR VPWR _16529_/C sky130_fd_sc_hd__o21ba_1
X_32565_ _36021_/CLK _32565_/D VGND VGND VPWR VPWR _32565_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_1209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17499_ _35646_/Q _35006_/Q _34366_/Q _33726_/Q _17497_/X _17498_/X VGND VGND VPWR
+ VPWR _17499_/X sky130_fd_sc_hd__mux4_1
XFILLER_220_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34304_ _34815_/CLK _34304_/D VGND VGND VPWR VPWR _34304_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31516_ _27785_/X _35972_/Q _31522_/S VGND VGND VPWR VPWR _31517_/A sky130_fd_sc_hd__mux2_1
X_19238_ _19234_/X _19237_/X _19098_/X VGND VGND VPWR VPWR _19248_/C sky130_fd_sc_hd__o21ba_1
X_35284_ _35668_/CLK _35284_/D VGND VGND VPWR VPWR _35284_/Q sky130_fd_sc_hd__dfxtp_1
X_32496_ _35952_/CLK _32496_/D VGND VGND VPWR VPWR _32496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34235_ _36157_/CLK _34235_/D VGND VGND VPWR VPWR _34235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19169_ _35436_/Q _35372_/Q _35308_/Q _35244_/Q _18848_/X _18849_/X VGND VGND VPWR
+ VPWR _19169_/X sky130_fd_sc_hd__mux4_1
X_31447_ _27683_/X _35939_/Q _31459_/S VGND VGND VPWR VPWR _31448_/A sky130_fd_sc_hd__mux2_1
X_21200_ _33381_/Q _33317_/Q _33253_/Q _33189_/Q _21021_/X _21022_/X VGND VGND VPWR
+ VPWR _21200_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22180_ _35200_/Q _35136_/Q _35072_/Q _32256_/Q _21963_/X _21964_/X VGND VGND VPWR
+ VPWR _22180_/X sky130_fd_sc_hd__mux4_1
X_34166_ _34166_/CLK _34166_/D VGND VGND VPWR VPWR _34166_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31378_ _31378_/A VGND VGND VPWR VPWR _35906_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_1138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33117_ _36054_/CLK _33117_/D VGND VGND VPWR VPWR _33117_/Q sky130_fd_sc_hd__dfxtp_1
X_21131_ _33635_/Q _33571_/Q _33507_/Q _33443_/Q _21094_/X _21095_/X VGND VGND VPWR
+ VPWR _21131_/X sky130_fd_sc_hd__mux4_1
XFILLER_191_1319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30329_ _35410_/Q _29515_/X _30335_/S VGND VGND VPWR VPWR _30330_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34097_ _35632_/CLK _34097_/D VGND VGND VPWR VPWR _34097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_236_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33048_ _35799_/CLK _33048_/D VGND VGND VPWR VPWR _33048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21062_ _21062_/A VGND VGND VPWR VPWR _36192_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20013_ _20009_/X _20010_/X _20011_/X _20012_/X VGND VGND VPWR VPWR _20013_/X sky130_fd_sc_hd__a22o_1
XFILLER_140_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25870_ _24883_/X _33393_/Q _25874_/S VGND VGND VPWR VPWR _25871_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_247_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24821_ input62/X VGND VGND VPWR VPWR _24821_/X sky130_fd_sc_hd__buf_2
XFILLER_58_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34999_ _35768_/CLK _34999_/D VGND VGND VPWR VPWR _34999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27540_ _27540_/A VGND VGND VPWR VPWR _34150_/D sky130_fd_sc_hd__clkbuf_1
X_21964_ _22317_/A VGND VGND VPWR VPWR _21964_/X sky130_fd_sc_hd__buf_6
X_24752_ _24752_/A VGND VGND VPWR VPWR _32896_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20915_ _34141_/Q _34077_/Q _34013_/Q _33949_/Q _20609_/X _20611_/X VGND VGND VPWR
+ VPWR _20915_/X sky130_fd_sc_hd__mux4_1
X_23703_ _23703_/A VGND VGND VPWR VPWR _32341_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27471_ _34118_/Q _27183_/X _27473_/S VGND VGND VPWR VPWR _27472_/A sky130_fd_sc_hd__mux2_1
XFILLER_214_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24683_ _24794_/S VGND VGND VPWR VPWR _24702_/S sky130_fd_sc_hd__buf_4
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21895_ _35192_/Q _35128_/Q _35064_/Q _32248_/Q _21610_/X _21611_/X VGND VGND VPWR
+ VPWR _21895_/X sky130_fd_sc_hd__mux4_1
XFILLER_81_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29210_ _29210_/A VGND VGND VPWR VPWR _34909_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26422_ _33654_/Q _23396_/X _26436_/S VGND VGND VPWR VPWR _26423_/A sky130_fd_sc_hd__mux2_1
X_23634_ _22980_/X _32308_/Q _23652_/S VGND VGND VPWR VPWR _23635_/A sky130_fd_sc_hd__mux2_1
X_20846_ _20740_/X _20844_/X _20845_/X _20745_/X VGND VGND VPWR VPWR _20846_/X sky130_fd_sc_hd__a22o_1
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29141_ _34877_/Q _27155_/X _29141_/S VGND VGND VPWR VPWR _29142_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23565_ _32277_/Q _23498_/X _23565_/S VGND VGND VPWR VPWR _23566_/A sky130_fd_sc_hd__mux2_1
X_26353_ _26353_/A VGND VGND VPWR VPWR _26486_/S sky130_fd_sc_hd__buf_12
X_20777_ _20777_/A VGND VGND VPWR VPWR _36184_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_35_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22516_ _22512_/X _22513_/X _22514_/X _22515_/X VGND VGND VPWR VPWR _22516_/X sky130_fd_sc_hd__a22o_1
X_25304_ _25304_/A VGND VGND VPWR VPWR _33125_/D sky130_fd_sc_hd__clkbuf_1
X_29072_ _34844_/Q _27053_/X _29078_/S VGND VGND VPWR VPWR _29073_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26284_ _24896_/X _33589_/Q _26300_/S VGND VGND VPWR VPWR _26285_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23496_ _32244_/Q _23495_/X _23499_/S VGND VGND VPWR VPWR _23497_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28023_ _34348_/Q _27103_/X _28037_/S VGND VGND VPWR VPWR _28024_/A sky130_fd_sc_hd__mux2_1
X_25235_ _25235_/A VGND VGND VPWR VPWR _33093_/D sky130_fd_sc_hd__clkbuf_1
X_22447_ _22447_/A VGND VGND VPWR VPWR _22447_/X sky130_fd_sc_hd__buf_2
XFILLER_6_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25166_ _25166_/A VGND VGND VPWR VPWR _33060_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22378_ _22373_/X _22375_/X _22376_/X _22377_/X VGND VGND VPWR VPWR _22378_/X sky130_fd_sc_hd__a22o_1
XFILLER_191_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24117_ _24117_/A VGND VGND VPWR VPWR _30877_/B sky130_fd_sc_hd__buf_8
XFILLER_124_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21329_ _21323_/X _21328_/X _21045_/X VGND VGND VPWR VPWR _21337_/C sky130_fd_sc_hd__o21ba_1
X_25097_ _24945_/X _33029_/Q _25101_/S VGND VGND VPWR VPWR _25098_/A sky130_fd_sc_hd__mux2_1
X_29974_ _29974_/A VGND VGND VPWR VPWR _35241_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28925_ _34774_/Q _27033_/X _28943_/S VGND VGND VPWR VPWR _28926_/A sky130_fd_sc_hd__mux2_1
X_24048_ _24048_/A VGND VGND VPWR VPWR _32565_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28856_ _28856_/A VGND VGND VPWR VPWR _34741_/D sky130_fd_sc_hd__clkbuf_1
X_16870_ _33068_/Q _32044_/Q _35820_/Q _35756_/Q _16725_/X _16726_/X VGND VGND VPWR
+ VPWR _16870_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27807_ input49/X VGND VGND VPWR VPWR _27807_/X sky130_fd_sc_hd__clkbuf_4
XTAP_4020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28787_ _28787_/A VGND VGND VPWR VPWR _31688_/A sky130_fd_sc_hd__buf_6
XFILLER_38_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25999_ _24874_/X _33454_/Q _26009_/S VGND VGND VPWR VPWR _26000_/A sky130_fd_sc_hd__mux2_1
XTAP_4053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18540_ _18391_/X _18538_/X _18539_/X _18401_/X VGND VGND VPWR VPWR _18540_/X sky130_fd_sc_hd__a22o_1
XTAP_4064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27738_ _27738_/A VGND VGND VPWR VPWR _34228_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_1042 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_218_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18471_ _19177_/A VGND VGND VPWR VPWR _18471_/X sky130_fd_sc_hd__buf_6
XTAP_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27669_ _27669_/A VGND VGND VPWR VPWR _34206_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_206_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29408_ _34991_/Q _29407_/X _29420_/S VGND VGND VPWR VPWR _29409_/A sky130_fd_sc_hd__mux2_1
X_17422_ _32124_/Q _32316_/Q _32380_/Q _35900_/Q _17280_/X _17421_/X VGND VGND VPWR
+ VPWR _17422_/X sky130_fd_sc_hd__mux4_1
XFILLER_205_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30680_ _35576_/Q _29435_/X _30690_/S VGND VGND VPWR VPWR _30681_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29339_ input34/X VGND VGND VPWR VPWR _29339_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17353_ _35642_/Q _35002_/Q _34362_/Q _33722_/Q _17144_/X _17145_/X VGND VGND VPWR
+ VPWR _17353_/X sky130_fd_sc_hd__mux4_1
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16304_ _17716_/A VGND VGND VPWR VPWR _16304_/X sky130_fd_sc_hd__buf_6
XFILLER_9_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32350_ _32802_/CLK _32350_/D VGND VGND VPWR VPWR _32350_/Q sky130_fd_sc_hd__dfxtp_1
X_17284_ _17279_/X _17283_/X _17140_/X _17141_/X VGND VGND VPWR VPWR _17301_/B sky130_fd_sc_hd__o211a_1
XFILLER_144_1398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31301_ _27667_/X _35870_/Q _31303_/S VGND VGND VPWR VPWR _31302_/A sky130_fd_sc_hd__mux2_1
X_19023_ _18945_/X _19021_/X _19022_/X _18948_/X VGND VGND VPWR VPWR _19023_/X sky130_fd_sc_hd__a22o_1
X_16235_ _34650_/Q _34586_/Q _34522_/Q _34458_/Q _16233_/X _16234_/X VGND VGND VPWR
+ VPWR _16235_/X sky130_fd_sc_hd__mux4_1
X_32281_ _35733_/CLK _32281_/D VGND VGND VPWR VPWR _32281_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34020_ _34148_/CLK _34020_/D VGND VGND VPWR VPWR _34020_/Q sky130_fd_sc_hd__dfxtp_1
X_31232_ _31232_/A VGND VGND VPWR VPWR _35837_/D sky130_fd_sc_hd__clkbuf_1
X_16166_ _16162_/X _16165_/X _16075_/X VGND VGND VPWR VPWR _16176_/C sky130_fd_sc_hd__o21ba_1
XFILLER_86_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31163_ _31163_/A VGND VGND VPWR VPWR _35804_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16097_ _17774_/A VGND VGND VPWR VPWR _17161_/A sky130_fd_sc_hd__buf_12
XFILLER_47_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30114_ _30114_/A VGND VGND VPWR VPWR _35307_/D sky130_fd_sc_hd__clkbuf_1
X_19925_ _33410_/Q _33346_/Q _33282_/Q _33218_/Q _19780_/X _19781_/X VGND VGND VPWR
+ VPWR _19925_/X sky130_fd_sc_hd__mux4_1
X_35971_ _36037_/CLK _35971_/D VGND VGND VPWR VPWR _35971_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31094_ _31094_/A VGND VGND VPWR VPWR _35772_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_296_CLK clkbuf_6_56__f_CLK/X VGND VGND VPWR VPWR _35779_/CLK sky130_fd_sc_hd__clkbuf_16
X_19856_ _34176_/Q _34112_/Q _34048_/Q _33984_/Q _19746_/X _19747_/X VGND VGND VPWR
+ VPWR _19856_/X sky130_fd_sc_hd__mux4_1
X_30045_ _35275_/Q _29494_/X _30057_/S VGND VGND VPWR VPWR _30046_/A sky130_fd_sc_hd__mux2_1
X_34922_ _35692_/CLK _34922_/D VGND VGND VPWR VPWR _34922_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18807_ _33122_/Q _36002_/Q _32994_/Q _32930_/Q _18656_/X _18657_/X VGND VGND VPWR
+ VPWR _18807_/X sky130_fd_sc_hd__mux4_1
X_19787_ _32638_/Q _32574_/Q _32510_/Q _35966_/Q _19576_/X _19713_/X VGND VGND VPWR
+ VPWR _19787_/X sky130_fd_sc_hd__mux4_1
X_34853_ _34920_/CLK _34853_/D VGND VGND VPWR VPWR _34853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16999_ _35696_/Q _32204_/Q _35568_/Q _35504_/Q _16964_/X _16965_/X VGND VGND VPWR
+ VPWR _16999_/X sky130_fd_sc_hd__mux4_1
XFILLER_62_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33804_ _36109_/CLK _33804_/D VGND VGND VPWR VPWR _33804_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18738_ _20298_/A VGND VGND VPWR VPWR _18738_/X sky130_fd_sc_hd__buf_6
X_34784_ _34915_/CLK _34784_/D VGND VGND VPWR VPWR _34784_/Q sky130_fd_sc_hd__dfxtp_1
X_31996_ _34405_/CLK _31996_/D VGND VGND VPWR VPWR _31996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33735_ _35715_/CLK _33735_/D VGND VGND VPWR VPWR _33735_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18669_ _35614_/Q _34974_/Q _34334_/Q _33694_/Q _18353_/X _18355_/X VGND VGND VPWR
+ VPWR _18669_/X sky130_fd_sc_hd__mux4_1
X_30947_ _30947_/A VGND VGND VPWR VPWR _35702_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20700_ _22377_/A VGND VGND VPWR VPWR _21763_/A sky130_fd_sc_hd__buf_12
XFILLER_34_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33666_ _36161_/CLK _33666_/D VGND VGND VPWR VPWR _33666_/Q sky130_fd_sc_hd__dfxtp_1
X_21680_ _33074_/Q _32050_/Q _35826_/Q _35762_/Q _21678_/X _21679_/X VGND VGND VPWR
+ VPWR _21680_/X sky130_fd_sc_hd__mux4_1
XFILLER_149_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30878_ _31010_/S VGND VGND VPWR VPWR _30897_/S sky130_fd_sc_hd__buf_6
X_35405_ _35853_/CLK _35405_/D VGND VGND VPWR VPWR _35405_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20631_ _20661_/A VGND VGND VPWR VPWR _22586_/A sky130_fd_sc_hd__buf_8
X_32617_ _35944_/CLK _32617_/D VGND VGND VPWR VPWR _32617_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33597_ _33661_/CLK _33597_/D VGND VGND VPWR VPWR _33597_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_220_CLK clkbuf_6_53__f_CLK/X VGND VGND VPWR VPWR _36173_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_162_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35336_ _35785_/CLK _35336_/D VGND VGND VPWR VPWR _35336_/Q sky130_fd_sc_hd__dfxtp_1
X_23350_ _23350_/A VGND VGND VPWR VPWR _32191_/D sky130_fd_sc_hd__clkbuf_1
X_20562_ _20558_/X _20561_/X _20146_/A _20147_/A VGND VGND VPWR VPWR _20577_/B sky130_fd_sc_hd__o211a_1
X_32548_ _35941_/CLK _32548_/D VGND VGND VPWR VPWR _32548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22301_ _32900_/Q _32836_/Q _32772_/Q _32708_/Q _22299_/X _22300_/X VGND VGND VPWR
+ VPWR _22301_/X sky130_fd_sc_hd__mux4_1
XFILLER_177_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35267_ _35716_/CLK _35267_/D VGND VGND VPWR VPWR _35267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23281_ _32166_/Q _23280_/X _23290_/S VGND VGND VPWR VPWR _23282_/A sky130_fd_sc_hd__mux2_1
X_20493_ _33939_/Q _33875_/Q _33811_/Q _36115_/Q _18362_/X _18364_/X VGND VGND VPWR
+ VPWR _20493_/X sky130_fd_sc_hd__mux4_1
XFILLER_164_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32479_ _35999_/CLK _32479_/D VGND VGND VPWR VPWR _32479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25020_ _24830_/X _32992_/Q _25038_/S VGND VGND VPWR VPWR _25021_/A sky130_fd_sc_hd__mux2_1
X_22232_ _22012_/X _22230_/X _22231_/X _22018_/X VGND VGND VPWR VPWR _22232_/X sky130_fd_sc_hd__a22o_1
XFILLER_117_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34218_ _36140_/CLK _34218_/D VGND VGND VPWR VPWR _34218_/Q sky130_fd_sc_hd__dfxtp_1
X_35198_ _36100_/CLK _35198_/D VGND VGND VPWR VPWR _35198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22163_ _22159_/X _22160_/X _22161_/X _22162_/X VGND VGND VPWR VPWR _22163_/X sky130_fd_sc_hd__a22o_1
X_34149_ _34149_/CLK _34149_/D VGND VGND VPWR VPWR _34149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21114_ _35618_/Q _34978_/Q _34338_/Q _33698_/Q _21038_/X _21039_/X VGND VGND VPWR
+ VPWR _21114_/X sky130_fd_sc_hd__mux4_1
XTAP_6917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22094_ _22447_/A VGND VGND VPWR VPWR _22094_/X sky130_fd_sc_hd__clkbuf_4
X_26971_ _33912_/Q _23402_/X _26981_/S VGND VGND VPWR VPWR _26972_/A sky130_fd_sc_hd__mux2_1
XTAP_6939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_287_CLK clkbuf_6_58__f_CLK/X VGND VGND VPWR VPWR _35839_/CLK sky130_fd_sc_hd__clkbuf_16
X_28710_ _28710_/A VGND VGND VPWR VPWR _34673_/D sky130_fd_sc_hd__clkbuf_1
X_25922_ _25922_/A VGND VGND VPWR VPWR _33417_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21045_ _22457_/A VGND VGND VPWR VPWR _21045_/X sky130_fd_sc_hd__buf_2
XFILLER_43_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29690_ _29690_/A VGND VGND VPWR VPWR _35106_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_247_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28641_ _28641_/A VGND VGND VPWR VPWR _34641_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25853_ _24858_/X _33385_/Q _25853_/S VGND VGND VPWR VPWR _25854_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24804_ _24803_/X _32919_/Q _24828_/S VGND VGND VPWR VPWR _24805_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_832 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28572_ _28572_/A VGND VGND VPWR VPWR _34608_/D sky130_fd_sc_hd__clkbuf_1
X_25784_ _24954_/X _33352_/Q _25802_/S VGND VGND VPWR VPWR _25785_/A sky130_fd_sc_hd__mux2_1
XFILLER_228_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22996_ input29/X VGND VGND VPWR VPWR _22996_/X sky130_fd_sc_hd__buf_2
XFILLER_227_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27523_ _27523_/A VGND VGND VPWR VPWR _34142_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24735_ _24735_/A VGND VGND VPWR VPWR _32888_/D sky130_fd_sc_hd__clkbuf_1
X_21947_ _22434_/A VGND VGND VPWR VPWR _21947_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27454_ _27502_/S VGND VGND VPWR VPWR _27473_/S sky130_fd_sc_hd__buf_6
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24666_ _24666_/A VGND VGND VPWR VPWR _32855_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_199_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_1338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21878_ _33144_/Q _36024_/Q _33016_/Q _32952_/Q _21662_/X _21663_/X VGND VGND VPWR
+ VPWR _21878_/X sky130_fd_sc_hd__mux4_1
XFILLER_203_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26405_ _33646_/Q _23305_/X _26415_/S VGND VGND VPWR VPWR _26406_/A sky130_fd_sc_hd__mux2_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20829_ _35418_/Q _35354_/Q _35290_/Q _35226_/Q _20795_/X _20796_/X VGND VGND VPWR
+ VPWR _20829_/X sky130_fd_sc_hd__mux4_1
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23617_ _22956_/X _32300_/Q _23631_/S VGND VGND VPWR VPWR _23618_/A sky130_fd_sc_hd__mux2_1
X_27385_ _34077_/Q _27056_/X _27389_/S VGND VGND VPWR VPWR _27386_/A sky130_fd_sc_hd__mux2_1
XFILLER_202_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24597_ _22990_/X _32823_/Q _24609_/S VGND VGND VPWR VPWR _24598_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_211_CLK clkbuf_6_52__f_CLK/X VGND VGND VPWR VPWR _35210_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_11_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29124_ _29124_/A VGND VGND VPWR VPWR _34868_/D sky130_fd_sc_hd__clkbuf_1
X_26336_ _24973_/X _33614_/Q _26342_/S VGND VGND VPWR VPWR _26337_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23548_ _23548_/A VGND VGND VPWR VPWR _32268_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29055_ _29055_/A VGND VGND VPWR VPWR _34836_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23479_ _32238_/Q _23478_/X _23485_/S VGND VGND VPWR VPWR _23480_/A sky130_fd_sc_hd__mux2_1
X_26267_ _24871_/X _33581_/Q _26279_/S VGND VGND VPWR VPWR _26268_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16020_ _17982_/A VGND VGND VPWR VPWR _17866_/A sky130_fd_sc_hd__buf_12
X_28006_ _34340_/Q _27078_/X _28016_/S VGND VGND VPWR VPWR _28007_/A sky130_fd_sc_hd__mux2_1
X_25218_ _25218_/A VGND VGND VPWR VPWR _33085_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26198_ _26198_/A VGND VGND VPWR VPWR _33548_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_1366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25149_ _25149_/A VGND VGND VPWR VPWR _33052_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17971_ _17864_/X _17969_/X _17970_/X _17869_/X VGND VGND VPWR VPWR _17971_/X sky130_fd_sc_hd__a22o_1
X_29957_ _35233_/Q _29364_/X _29973_/S VGND VGND VPWR VPWR _29958_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_1322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_278_CLK clkbuf_6_59__f_CLK/X VGND VGND VPWR VPWR _33924_/CLK sky130_fd_sc_hd__clkbuf_16
X_19710_ _19506_/X _19708_/X _19709_/X _19509_/X VGND VGND VPWR VPWR _19710_/X sky130_fd_sc_hd__a22o_1
X_28908_ _28908_/A VGND VGND VPWR VPWR _34766_/D sky130_fd_sc_hd__clkbuf_1
X_16922_ _16918_/X _16921_/X _16779_/X VGND VGND VPWR VPWR _16948_/A sky130_fd_sc_hd__o21ba_1
X_29888_ _29888_/A VGND VGND VPWR VPWR _35200_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19641_ _19637_/X _19640_/X _19432_/X VGND VGND VPWR VPWR _19671_/A sky130_fd_sc_hd__o21ba_1
XFILLER_38_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16853_ _17912_/A VGND VGND VPWR VPWR _16853_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_4_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28839_ _28839_/A VGND VGND VPWR VPWR _34733_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19572_ _33400_/Q _33336_/Q _33272_/Q _33208_/Q _19427_/X _19428_/X VGND VGND VPWR
+ VPWR _19572_/X sky130_fd_sc_hd__mux4_1
X_31850_ _23268_/X _36130_/Q _31864_/S VGND VGND VPWR VPWR _31851_/A sky130_fd_sc_hd__mux2_1
X_16784_ _32106_/Q _32298_/Q _32362_/Q _35882_/Q _16574_/X _16715_/X VGND VGND VPWR
+ VPWR _16784_/X sky130_fd_sc_hd__mux4_1
XFILLER_219_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_1394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18523_ _32858_/Q _32794_/Q _32730_/Q _32666_/Q _18337_/X _18339_/X VGND VGND VPWR
+ VPWR _18523_/X sky130_fd_sc_hd__mux4_1
X_30801_ _30801_/A VGND VGND VPWR VPWR _35633_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31781_ _31781_/A VGND VGND VPWR VPWR _36097_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33520_ _36080_/CLK _33520_/D VGND VGND VPWR VPWR _33520_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_450_CLK clkbuf_6_14__f_CLK/X VGND VGND VPWR VPWR _36015_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18454_ _33112_/Q _35992_/Q _32984_/Q _32920_/Q _18324_/X _18325_/X VGND VGND VPWR
+ VPWR _18454_/X sky130_fd_sc_hd__mux4_1
X_30732_ _35601_/Q _29512_/X _30732_/S VGND VGND VPWR VPWR _30733_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17405_ _33660_/Q _33596_/Q _33532_/Q _33468_/Q _17200_/X _17201_/X VGND VGND VPWR
+ VPWR _17405_/X sky130_fd_sc_hd__mux4_1
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33451_ _34153_/CLK _33451_/D VGND VGND VPWR VPWR _33451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18385_ _19311_/A VGND VGND VPWR VPWR _18385_/X sky130_fd_sc_hd__buf_4
X_30663_ _35568_/Q _29410_/X _30669_/S VGND VGND VPWR VPWR _30664_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_202_CLK clkbuf_6_51__f_CLK/X VGND VGND VPWR VPWR _35466_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32402_ _35922_/CLK _32402_/D VGND VGND VPWR VPWR _32402_/Q sky130_fd_sc_hd__dfxtp_1
X_36170_ _36171_/CLK _36170_/D VGND VGND VPWR VPWR _36170_/Q sky130_fd_sc_hd__dfxtp_1
X_17336_ _34170_/Q _34106_/Q _34042_/Q _33978_/Q _17093_/X _17094_/X VGND VGND VPWR
+ VPWR _17336_/X sky130_fd_sc_hd__mux4_1
XFILLER_60_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33382_ _33697_/CLK _33382_/D VGND VGND VPWR VPWR _33382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30594_ _30594_/A VGND VGND VPWR VPWR _35535_/D sky130_fd_sc_hd__clkbuf_1
X_35121_ _35377_/CLK _35121_/D VGND VGND VPWR VPWR _35121_/Q sky130_fd_sc_hd__dfxtp_1
X_32333_ _35916_/CLK _32333_/D VGND VGND VPWR VPWR _32333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17267_ _17267_/A _17267_/B _17267_/C _17267_/D VGND VGND VPWR VPWR _17268_/A sky130_fd_sc_hd__or4_4
XFILLER_88_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1050 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19006_ _20205_/A VGND VGND VPWR VPWR _19006_/X sky130_fd_sc_hd__clkbuf_4
X_16218_ _32602_/Q _32538_/Q _32474_/Q _35930_/Q _16217_/X _17717_/A VGND VGND VPWR
+ VPWR _16218_/X sky130_fd_sc_hd__mux4_1
X_35052_ _35564_/CLK _35052_/D VGND VGND VPWR VPWR _35052_/Q sky130_fd_sc_hd__dfxtp_1
X_32264_ _35212_/CLK _32264_/D VGND VGND VPWR VPWR _32264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17198_ _17198_/A VGND VGND VPWR VPWR _31989_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34003_ _34897_/CLK _34003_/D VGND VGND VPWR VPWR _34003_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31215_ _27739_/X _35829_/Q _31231_/S VGND VGND VPWR VPWR _31216_/A sky130_fd_sc_hd__mux2_1
X_16149_ _33880_/Q _33816_/Q _33752_/Q _36056_/Q _16112_/X _16113_/X VGND VGND VPWR
+ VPWR _16149_/X sky130_fd_sc_hd__mux4_1
XFILLER_127_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32195_ _35687_/CLK _32195_/D VGND VGND VPWR VPWR _32195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_216_1108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31146_ _31146_/A VGND VGND VPWR VPWR _35797_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_269_CLK clkbuf_6_60__f_CLK/X VGND VGND VPWR VPWR _34691_/CLK sky130_fd_sc_hd__clkbuf_16
X_19908_ _20261_/A VGND VGND VPWR VPWR _19908_/X sky130_fd_sc_hd__buf_4
X_31077_ _35764_/Q input24/X _31095_/S VGND VGND VPWR VPWR _31078_/A sky130_fd_sc_hd__mux2_1
X_35954_ _35955_/CLK _35954_/D VGND VGND VPWR VPWR _35954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_233_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34905_ _34907_/CLK _34905_/D VGND VGND VPWR VPWR _34905_/Q sky130_fd_sc_hd__dfxtp_1
X_30028_ _35267_/Q _29469_/X _30036_/S VGND VGND VPWR VPWR _30029_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19839_ _35455_/Q _35391_/Q _35327_/Q _35263_/Q _19554_/X _19555_/X VGND VGND VPWR
+ VPWR _19839_/X sky130_fd_sc_hd__mux4_1
XFILLER_232_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35885_ _35951_/CLK _35885_/D VGND VGND VPWR VPWR _35885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34836_ _34964_/CLK _34836_/D VGND VGND VPWR VPWR _34836_/Q sky130_fd_sc_hd__dfxtp_1
X_22850_ _34197_/Q _34133_/Q _34069_/Q _34005_/Q _20649_/X _20650_/X VGND VGND VPWR
+ VPWR _22850_/X sky130_fd_sc_hd__mux4_1
XFILLER_232_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21801_ _22507_/A VGND VGND VPWR VPWR _21801_/X sky130_fd_sc_hd__buf_4
XFILLER_232_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22781_ _35218_/Q _35154_/Q _35090_/Q _32274_/Q _20692_/X _20694_/X VGND VGND VPWR
+ VPWR _22781_/X sky130_fd_sc_hd__mux4_1
XFILLER_37_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34767_ _34961_/CLK _34767_/D VGND VGND VPWR VPWR _34767_/Q sky130_fd_sc_hd__dfxtp_1
X_31979_ _34790_/CLK _31979_/D VGND VGND VPWR VPWR _31979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_441_CLK clkbuf_6_37__f_CLK/X VGND VGND VPWR VPWR _35953_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_225_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24520_ _23076_/X _32787_/Q _24524_/S VGND VGND VPWR VPWR _24521_/A sky130_fd_sc_hd__mux2_1
X_21732_ _22438_/A VGND VGND VPWR VPWR _21732_/X sky130_fd_sc_hd__clkbuf_4
X_33718_ _35703_/CLK _33718_/D VGND VGND VPWR VPWR _33718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34698_ _34698_/CLK _34698_/D VGND VGND VPWR VPWR _34698_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21663_ _22374_/A VGND VGND VPWR VPWR _21663_/X sky130_fd_sc_hd__clkbuf_4
X_24451_ _22974_/X _32754_/Q _24453_/S VGND VGND VPWR VPWR _24452_/A sky130_fd_sc_hd__mux2_1
X_33649_ _34098_/CLK _33649_/D VGND VGND VPWR VPWR _33649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20614_ input75/X input76/X VGND VGND VPWR VPWR _22438_/A sky130_fd_sc_hd__or2b_4
X_23402_ input28/X VGND VGND VPWR VPWR _23402_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_71_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27170_ _27170_/A VGND VGND VPWR VPWR _33985_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24382_ _24382_/A VGND VGND VPWR VPWR _32721_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21594_ _22434_/A VGND VGND VPWR VPWR _21594_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_71_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23333_ _32184_/Q _23255_/X _23335_/S VGND VGND VPWR VPWR _23334_/A sky130_fd_sc_hd__mux2_1
X_26121_ _24855_/X _33512_/Q _26123_/S VGND VGND VPWR VPWR _26122_/A sky130_fd_sc_hd__mux2_1
X_20545_ _18360_/X _20543_/X _20544_/X _18372_/X VGND VGND VPWR VPWR _20545_/X sky130_fd_sc_hd__a22o_1
XFILLER_137_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35319_ _35769_/CLK _35319_/D VGND VGND VPWR VPWR _35319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26052_ _26052_/A VGND VGND VPWR VPWR _33479_/D sky130_fd_sc_hd__clkbuf_1
X_23264_ _23264_/A VGND VGND VPWR VPWR _32160_/D sky130_fd_sc_hd__clkbuf_1
X_20476_ _35474_/Q _35410_/Q _35346_/Q _35282_/Q _20260_/X _20261_/X VGND VGND VPWR
+ VPWR _20476_/X sky130_fd_sc_hd__mux4_1
XFILLER_106_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25003_ _24806_/X _32984_/Q _25017_/S VGND VGND VPWR VPWR _25004_/A sky130_fd_sc_hd__mux2_1
X_22215_ _22106_/X _22213_/X _22214_/X _22109_/X VGND VGND VPWR VPWR _22215_/X sky130_fd_sc_hd__a22o_1
XFILLER_152_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23195_ _23195_/A VGND VGND VPWR VPWR _32135_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29811_ _35164_/Q _29348_/X _29817_/S VGND VGND VPWR VPWR _29812_/A sky130_fd_sc_hd__mux2_1
XTAP_6703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22146_ _34431_/Q _36159_/Q _34303_/Q _34239_/Q _21829_/X _21830_/X VGND VGND VPWR
+ VPWR _22146_/X sky130_fd_sc_hd__mux4_1
XFILLER_105_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29742_ _29742_/A VGND VGND VPWR VPWR _35131_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_248_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26954_ _33904_/Q _23340_/X _26960_/S VGND VGND VPWR VPWR _26955_/A sky130_fd_sc_hd__mux2_1
X_22077_ _33662_/Q _33598_/Q _33534_/Q _33470_/Q _21800_/X _21801_/X VGND VGND VPWR
+ VPWR _22077_/X sky130_fd_sc_hd__mux4_1
XTAP_6769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25905_ _25905_/A VGND VGND VPWR VPWR _33409_/D sky130_fd_sc_hd__clkbuf_1
X_21028_ _32608_/Q _32544_/Q _32480_/Q _35936_/Q _20817_/X _20954_/X VGND VGND VPWR
+ VPWR _21028_/X sky130_fd_sc_hd__mux4_1
X_29673_ _29673_/A VGND VGND VPWR VPWR _35098_/D sky130_fd_sc_hd__clkbuf_1
X_26885_ _26885_/A VGND VGND VPWR VPWR _33871_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28624_ _27801_/X _34633_/Q _28640_/S VGND VGND VPWR VPWR _28625_/A sky130_fd_sc_hd__mux2_1
X_25836_ _25836_/A VGND VGND VPWR VPWR _33376_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_216_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28555_ _28555_/A VGND VGND VPWR VPWR _34600_/D sky130_fd_sc_hd__clkbuf_1
X_25767_ _24930_/X _33344_/Q _25781_/S VGND VGND VPWR VPWR _25768_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22979_ _22979_/A VGND VGND VPWR VPWR _32051_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_432_CLK clkbuf_6_36__f_CLK/X VGND VGND VPWR VPWR _36019_/CLK sky130_fd_sc_hd__clkbuf_16
X_27506_ _34134_/Q _27033_/X _27524_/S VGND VGND VPWR VPWR _27507_/A sky130_fd_sc_hd__mux2_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_231_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24718_ _24718_/A VGND VGND VPWR VPWR _32880_/D sky130_fd_sc_hd__clkbuf_1
X_28486_ _28513_/S VGND VGND VPWR VPWR _28505_/S sky130_fd_sc_hd__buf_4
XFILLER_203_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25698_ _25698_/A VGND VGND VPWR VPWR _33311_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27437_ _27437_/A VGND VGND VPWR VPWR _34101_/D sky130_fd_sc_hd__clkbuf_1
X_24649_ _23067_/X _32848_/Q _24651_/S VGND VGND VPWR VPWR _24650_/A sky130_fd_sc_hd__mux2_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18170_ _32914_/Q _32850_/Q _32786_/Q _32722_/Q _15984_/X _15987_/X VGND VGND VPWR
+ VPWR _18170_/X sky130_fd_sc_hd__mux4_1
X_27368_ _27368_/A VGND VGND VPWR VPWR _34069_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_230_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29107_ _29107_/A VGND VGND VPWR VPWR _34860_/D sky130_fd_sc_hd__clkbuf_1
X_17121_ _17117_/X _17120_/X _16812_/X VGND VGND VPWR VPWR _17122_/D sky130_fd_sc_hd__o21ba_1
X_26319_ _24948_/X _33606_/Q _26321_/S VGND VGND VPWR VPWR _26320_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_1078 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27299_ _34036_/Q _27127_/X _27317_/S VGND VGND VPWR VPWR _27300_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_6_35__f_CLK clkbuf_5_17_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_35__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_7_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29038_ _34828_/Q _27202_/X _29048_/S VGND VGND VPWR VPWR _29039_/A sky130_fd_sc_hd__mux2_1
X_17052_ _33650_/Q _33586_/Q _33522_/Q _33458_/Q _16847_/X _16848_/X VGND VGND VPWR
+ VPWR _17052_/X sky130_fd_sc_hd__mux4_1
XFILLER_156_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16003_ _17800_/A VGND VGND VPWR VPWR _16003_/X sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_499_CLK clkbuf_6_2__f_CLK/X VGND VGND VPWR VPWR _36073_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_100_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31000_ _35728_/Q input54/X _31002_/S VGND VGND VPWR VPWR _31001_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17954_ _32907_/Q _32843_/Q _32779_/Q _32715_/Q _17699_/X _17700_/X VGND VGND VPWR
+ VPWR _17954_/X sky130_fd_sc_hd__mux4_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16905_ _16650_/X _16903_/X _16904_/X _16653_/X VGND VGND VPWR VPWR _16905_/X sky130_fd_sc_hd__a22o_1
XFILLER_111_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32951_ _36024_/CLK _32951_/D VGND VGND VPWR VPWR _32951_/Q sky130_fd_sc_hd__dfxtp_1
X_17885_ _32137_/Q _32329_/Q _32393_/Q _35913_/Q _17633_/X _17774_/X VGND VGND VPWR
+ VPWR _17885_/X sky130_fd_sc_hd__mux4_1
XFILLER_120_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31902_ _23411_/X _36155_/Q _31906_/S VGND VGND VPWR VPWR _31903_/A sky130_fd_sc_hd__mux2_1
X_19624_ _19303_/X _19622_/X _19623_/X _19306_/X VGND VGND VPWR VPWR _19624_/X sky130_fd_sc_hd__a22o_1
X_16836_ _16832_/X _16835_/X _16798_/X VGND VGND VPWR VPWR _16844_/C sky130_fd_sc_hd__o21ba_1
XFILLER_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35670_ _35735_/CLK _35670_/D VGND VGND VPWR VPWR _35670_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32882_ _32882_/CLK _32882_/D VGND VGND VPWR VPWR _32882_/Q sky130_fd_sc_hd__dfxtp_1
X_31833_ _23243_/X _36122_/Q _31843_/S VGND VGND VPWR VPWR _31834_/A sky130_fd_sc_hd__mux2_1
XFILLER_207_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34621_ _36153_/CLK _34621_/D VGND VGND VPWR VPWR _34621_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19555_ _20261_/A VGND VGND VPWR VPWR _19555_/X sky130_fd_sc_hd__buf_4
XFILLER_202_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16767_ _16452_/X _16765_/X _16766_/X _16457_/X VGND VGND VPWR VPWR _16767_/X sky130_fd_sc_hd__a22o_1
XFILLER_81_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18506_ _18391_/X _18504_/X _18505_/X _18401_/X VGND VGND VPWR VPWR _18506_/X sky130_fd_sc_hd__a22o_1
XFILLER_206_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_423_CLK clkbuf_6_33__f_CLK/X VGND VGND VPWR VPWR _35634_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_59_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34552_ _35193_/CLK _34552_/D VGND VGND VPWR VPWR _34552_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_1134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31764_ _31764_/A VGND VGND VPWR VPWR _36089_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19486_ _35445_/Q _35381_/Q _35317_/Q _35253_/Q _19201_/X _19202_/X VGND VGND VPWR
+ VPWR _19486_/X sky130_fd_sc_hd__mux4_1
X_16698_ _16698_/A VGND VGND VPWR VPWR _31975_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_1107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18437_ _18433_/X _18436_/X _18404_/X VGND VGND VPWR VPWR _18438_/D sky130_fd_sc_hd__o21ba_1
X_30715_ _30715_/A VGND VGND VPWR VPWR _35592_/D sky130_fd_sc_hd__clkbuf_1
X_33503_ _36191_/CLK _33503_/D VGND VGND VPWR VPWR _33503_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34483_ _34611_/CLK _34483_/D VGND VGND VPWR VPWR _34483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31695_ _31695_/A VGND VGND VPWR VPWR _36056_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36222_ _36229_/CLK _36222_/D VGND VGND VPWR VPWR _36222_/Q sky130_fd_sc_hd__dfxtp_1
X_33434_ _36212_/CLK _33434_/D VGND VGND VPWR VPWR _33434_/Q sky130_fd_sc_hd__dfxtp_1
X_30646_ _35560_/Q _29385_/X _30648_/S VGND VGND VPWR VPWR _30647_/A sky130_fd_sc_hd__mux2_1
X_18368_ _20066_/A VGND VGND VPWR VPWR _20236_/A sky130_fd_sc_hd__buf_12
XFILLER_33_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36153_ _36153_/CLK _36153_/D VGND VGND VPWR VPWR _36153_/Q sky130_fd_sc_hd__dfxtp_1
X_17319_ _35705_/Q _32214_/Q _35577_/Q _35513_/Q _17317_/X _17318_/X VGND VGND VPWR
+ VPWR _17319_/X sky130_fd_sc_hd__mux4_2
X_33365_ _33685_/CLK _33365_/D VGND VGND VPWR VPWR _33365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30577_ _30577_/A VGND VGND VPWR VPWR _35527_/D sky130_fd_sc_hd__clkbuf_1
X_18299_ _18299_/A VGND VGND VPWR VPWR _20073_/A sky130_fd_sc_hd__buf_2
XFILLER_30_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20330_ _34701_/Q _34637_/Q _34573_/Q _34509_/Q _20298_/X _20299_/X VGND VGND VPWR
+ VPWR _20330_/X sky130_fd_sc_hd__mux4_1
X_35104_ _35168_/CLK _35104_/D VGND VGND VPWR VPWR _35104_/Q sky130_fd_sc_hd__dfxtp_1
X_32316_ _35964_/CLK _32316_/D VGND VGND VPWR VPWR _32316_/Q sky130_fd_sc_hd__dfxtp_1
X_36084_ _36085_/CLK _36084_/D VGND VGND VPWR VPWR _36084_/Q sky130_fd_sc_hd__dfxtp_1
X_33296_ _34186_/CLK _33296_/D VGND VGND VPWR VPWR _33296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35035_ _35482_/CLK _35035_/D VGND VGND VPWR VPWR _35035_/Q sky130_fd_sc_hd__dfxtp_1
X_20261_ _20261_/A VGND VGND VPWR VPWR _20261_/X sky130_fd_sc_hd__clkbuf_4
X_32247_ _36024_/CLK _32247_/D VGND VGND VPWR VPWR _32247_/Q sky130_fd_sc_hd__dfxtp_1
X_22000_ _34939_/Q _34875_/Q _34811_/Q _34747_/Q _21760_/X _21761_/X VGND VGND VPWR
+ VPWR _22000_/X sky130_fd_sc_hd__mux4_1
XFILLER_192_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32178_ _35482_/CLK _32178_/D VGND VGND VPWR VPWR _32178_/Q sky130_fd_sc_hd__dfxtp_1
X_20192_ _35465_/Q _35401_/Q _35337_/Q _35273_/Q _19907_/X _19908_/X VGND VGND VPWR
+ VPWR _20192_/X sky130_fd_sc_hd__mux4_1
XFILLER_153_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_935 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31129_ _35789_/Q input51/X _31137_/S VGND VGND VPWR VPWR _31130_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23951_ _23042_/X _32520_/Q _23969_/S VGND VGND VPWR VPWR _23952_/A sky130_fd_sc_hd__mux2_1
X_35937_ _35938_/CLK _35937_/D VGND VGND VPWR VPWR _35937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22902_ _22902_/A VGND VGND VPWR VPWR _32026_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26670_ _26670_/A VGND VGND VPWR VPWR _33769_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35868_ _35997_/CLK _35868_/D VGND VGND VPWR VPWR _35868_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23882_ _23882_/A VGND VGND VPWR VPWR _32487_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25621_ _24914_/X _33275_/Q _25625_/S VGND VGND VPWR VPWR _25622_/A sky130_fd_sc_hd__mux2_1
X_34819_ _34949_/CLK _34819_/D VGND VGND VPWR VPWR _34819_/Q sky130_fd_sc_hd__dfxtp_1
X_22833_ _35732_/Q _32244_/Q _35604_/Q _35540_/Q _20593_/X _20595_/X VGND VGND VPWR
+ VPWR _22833_/X sky130_fd_sc_hd__mux4_1
XFILLER_186_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_1048 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35799_ _35799_/CLK _35799_/D VGND VGND VPWR VPWR _35799_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_414_CLK clkbuf_6_32__f_CLK/X VGND VGND VPWR VPWR _34035_/CLK sky130_fd_sc_hd__clkbuf_16
X_28340_ _28340_/A VGND VGND VPWR VPWR _34498_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25552_ _24812_/X _33242_/Q _25562_/S VGND VGND VPWR VPWR _25553_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22764_ _22512_/X _22762_/X _22763_/X _22515_/X VGND VGND VPWR VPWR _22764_/X sky130_fd_sc_hd__a22o_1
XFILLER_168_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24503_ _24503_/A VGND VGND VPWR VPWR _32778_/D sky130_fd_sc_hd__clkbuf_1
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21715_ _34675_/Q _34611_/Q _34547_/Q _34483_/Q _21539_/X _21540_/X VGND VGND VPWR
+ VPWR _21715_/X sky130_fd_sc_hd__mux4_1
X_28271_ _28271_/A VGND VGND VPWR VPWR _34465_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_241_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22695_ _22464_/X _22693_/X _22694_/X _22469_/X VGND VGND VPWR VPWR _22695_/X sky130_fd_sc_hd__a22o_1
XFILLER_13_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25483_ _25483_/A VGND VGND VPWR VPWR _33209_/D sky130_fd_sc_hd__clkbuf_1
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27222_ _27222_/A VGND VGND VPWR VPWR _34002_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24434_ _24524_/S VGND VGND VPWR VPWR _24453_/S sky130_fd_sc_hd__buf_4
XFILLER_40_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21646_ _34417_/Q _36145_/Q _34289_/Q _34225_/Q _21476_/X _21477_/X VGND VGND VPWR
+ VPWR _21646_/X sky130_fd_sc_hd__mux4_1
XFILLER_12_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1062 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27153_ _33980_/Q _27152_/X _27156_/S VGND VGND VPWR VPWR _27154_/A sky130_fd_sc_hd__mux2_1
X_24365_ _23046_/X _32713_/Q _24381_/S VGND VGND VPWR VPWR _24366_/A sky130_fd_sc_hd__mux2_1
X_21577_ _34927_/Q _34863_/Q _34799_/Q _34735_/Q _21407_/X _21408_/X VGND VGND VPWR
+ VPWR _21577_/X sky130_fd_sc_hd__mux4_1
XFILLER_193_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26104_ _26215_/S VGND VGND VPWR VPWR _26123_/S sky130_fd_sc_hd__buf_6
XFILLER_193_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20528_ _19453_/A _20526_/X _20527_/X _19456_/A VGND VGND VPWR VPWR _20528_/X sky130_fd_sc_hd__a22o_1
X_23316_ input18/X VGND VGND VPWR VPWR _23316_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_138_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24296_ _24296_/A VGND VGND VPWR VPWR _32680_/D sky130_fd_sc_hd__clkbuf_1
X_27084_ input8/X VGND VGND VPWR VPWR _27084_/X sky130_fd_sc_hd__buf_2
XFILLER_153_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26035_ _24927_/X _33471_/Q _26051_/S VGND VGND VPWR VPWR _26036_/A sky130_fd_sc_hd__mux2_1
X_20459_ _33682_/Q _33618_/Q _33554_/Q _33490_/Q _20206_/X _20207_/X VGND VGND VPWR
+ VPWR _20459_/X sky130_fd_sc_hd__mux4_1
X_23247_ _32155_/Q _23246_/X _23259_/S VGND VGND VPWR VPWR _23248_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23178_ _23015_/X _32127_/Q _23194_/S VGND VGND VPWR VPWR _23179_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22129_ _32639_/Q _32575_/Q _32511_/Q _35967_/Q _21876_/X _22013_/X VGND VGND VPWR
+ VPWR _22129_/X sky130_fd_sc_hd__mux4_1
XTAP_6544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27986_ _27986_/A VGND VGND VPWR VPWR _34330_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29725_ _29725_/A VGND VGND VPWR VPWR _35123_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26937_ _33896_/Q _23286_/X _26939_/S VGND VGND VPWR VPWR _26938_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_248_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29656_ _35091_/Q _29518_/X _29660_/S VGND VGND VPWR VPWR _29657_/A sky130_fd_sc_hd__mux2_1
X_17670_ _17799_/A VGND VGND VPWR VPWR _17670_/X sky130_fd_sc_hd__buf_4
XFILLER_43_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26868_ _26868_/A VGND VGND VPWR VPWR _33863_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28607_ _27776_/X _34625_/Q _28619_/S VGND VGND VPWR VPWR _28608_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16621_ _35173_/Q _35109_/Q _35045_/Q _32165_/Q _16304_/X _16305_/X VGND VGND VPWR
+ VPWR _16621_/X sky130_fd_sc_hd__mux4_1
X_25819_ _25819_/A VGND VGND VPWR VPWR _33368_/D sky130_fd_sc_hd__clkbuf_1
X_29587_ _35058_/Q _29416_/X _29589_/S VGND VGND VPWR VPWR _29588_/A sky130_fd_sc_hd__mux2_1
X_26799_ _26799_/A VGND VGND VPWR VPWR _33830_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_405_CLK clkbuf_6_34__f_CLK/X VGND VGND VPWR VPWR _34100_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_210_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_902 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_941 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19340_ _33073_/Q _32049_/Q _35825_/Q _35761_/Q _19025_/X _19026_/X VGND VGND VPWR
+ VPWR _19340_/X sky130_fd_sc_hd__mux4_1
XFILLER_16_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16552_ _16297_/X _16550_/X _16551_/X _16300_/X VGND VGND VPWR VPWR _16552_/X sky130_fd_sc_hd__a22o_1
XFILLER_95_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28538_ _27673_/X _34592_/Q _28556_/S VGND VGND VPWR VPWR _28539_/A sky130_fd_sc_hd__mux2_1
XFILLER_244_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_245_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19271_ _18950_/X _19269_/X _19270_/X _18953_/X VGND VGND VPWR VPWR _19271_/X sky130_fd_sc_hd__a22o_1
XFILLER_91_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28469_ _28469_/A VGND VGND VPWR VPWR _34559_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16483_ _16479_/X _16482_/X _16445_/X VGND VGND VPWR VPWR _16491_/C sky130_fd_sc_hd__o21ba_1
X_18222_ _33428_/Q _33364_/Q _33300_/Q _33236_/Q _16037_/X _16039_/X VGND VGND VPWR
+ VPWR _18222_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30500_ _30500_/A VGND VGND VPWR VPWR _35490_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31480_ _27732_/X _35955_/Q _31480_/S VGND VGND VPWR VPWR _31481_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18153_ _34449_/Q _36177_/Q _34321_/Q _34257_/Q _17935_/X _17936_/X VGND VGND VPWR
+ VPWR _18153_/X sky130_fd_sc_hd__mux4_1
X_30431_ _35458_/Q _29466_/X _30441_/S VGND VGND VPWR VPWR _30432_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17104_ _32115_/Q _32307_/Q _32371_/Q _35891_/Q _16927_/X _17068_/X VGND VGND VPWR
+ VPWR _17104_/X sky130_fd_sc_hd__mux4_1
XFILLER_106_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33150_ _36031_/CLK _33150_/D VGND VGND VPWR VPWR _33150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18084_ _35663_/Q _35023_/Q _34383_/Q _33743_/Q _17850_/X _17851_/X VGND VGND VPWR
+ VPWR _18084_/X sky130_fd_sc_hd__mux4_1
X_30362_ _35425_/Q _29364_/X _30378_/S VGND VGND VPWR VPWR _30363_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32101_ _35945_/CLK _32101_/D VGND VGND VPWR VPWR _32101_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17035_ _17031_/X _17034_/X _16787_/X _16788_/X VGND VGND VPWR VPWR _17050_/B sky130_fd_sc_hd__o211a_1
X_33081_ _35833_/CLK _33081_/D VGND VGND VPWR VPWR _33081_/Q sky130_fd_sc_hd__dfxtp_1
X_30293_ _30293_/A VGND VGND VPWR VPWR _35392_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32032_ _35941_/CLK _32032_/D VGND VGND VPWR VPWR _32032_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18986_ _35431_/Q _35367_/Q _35303_/Q _35239_/Q _18848_/X _18849_/X VGND VGND VPWR
+ VPWR _18986_/X sky130_fd_sc_hd__mux4_1
XFILLER_140_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17937_ _34442_/Q _36170_/Q _34314_/Q _34250_/Q _17935_/X _17936_/X VGND VGND VPWR
+ VPWR _17937_/X sky130_fd_sc_hd__mux4_1
XFILLER_140_798 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33983_ _35454_/CLK _33983_/D VGND VGND VPWR VPWR _33983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35722_ _35722_/CLK _35722_/D VGND VGND VPWR VPWR _35722_/Q sky130_fd_sc_hd__dfxtp_1
X_17868_ _34952_/Q _34888_/Q _34824_/Q _34760_/Q _17866_/X _17867_/X VGND VGND VPWR
+ VPWR _17868_/X sky130_fd_sc_hd__mux4_1
XFILLER_27_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32934_ _36003_/CLK _32934_/D VGND VGND VPWR VPWR _32934_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19607_ _33913_/Q _33849_/Q _33785_/Q _36089_/Q _19324_/X _19325_/X VGND VGND VPWR
+ VPWR _19607_/X sky130_fd_sc_hd__mux4_1
X_35653_ _35655_/CLK _35653_/D VGND VGND VPWR VPWR _35653_/Q sky130_fd_sc_hd__dfxtp_1
X_16819_ _33387_/Q _33323_/Q _33259_/Q _33195_/Q _16774_/X _16775_/X VGND VGND VPWR
+ VPWR _16819_/X sky130_fd_sc_hd__mux4_1
X_17799_ _17799_/A VGND VGND VPWR VPWR _17799_/X sky130_fd_sc_hd__clkbuf_8
X_32865_ _35871_/CLK _32865_/D VGND VGND VPWR VPWR _32865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34604_ _36140_/CLK _34604_/D VGND VGND VPWR VPWR _34604_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31816_ _31816_/A VGND VGND VPWR VPWR _36114_/D sky130_fd_sc_hd__clkbuf_1
X_19538_ _34167_/Q _34103_/Q _34039_/Q _33975_/Q _19393_/X _19394_/X VGND VGND VPWR
+ VPWR _19538_/X sky130_fd_sc_hd__mux4_1
XFILLER_81_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35584_ _35713_/CLK _35584_/D VGND VGND VPWR VPWR _35584_/Q sky130_fd_sc_hd__dfxtp_1
X_32796_ _36053_/CLK _32796_/D VGND VGND VPWR VPWR _32796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19469_ _33653_/Q _33589_/Q _33525_/Q _33461_/Q _19147_/X _19148_/X VGND VGND VPWR
+ VPWR _19469_/X sky130_fd_sc_hd__mux4_1
X_31747_ _31747_/A VGND VGND VPWR VPWR _36081_/D sky130_fd_sc_hd__clkbuf_1
X_34535_ _35365_/CLK _34535_/D VGND VGND VPWR VPWR _34535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21500_ _21245_/X _21498_/X _21499_/X _21248_/X VGND VGND VPWR VPWR _21500_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22480_ _22159_/X _22478_/X _22479_/X _22162_/X VGND VGND VPWR VPWR _22480_/X sky130_fd_sc_hd__a22o_1
X_31678_ _27825_/X _36049_/Q _31678_/S VGND VGND VPWR VPWR _31679_/A sky130_fd_sc_hd__mux2_1
X_34466_ _36209_/CLK _34466_/D VGND VGND VPWR VPWR _34466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36205_ _36205_/CLK _36205_/D VGND VGND VPWR VPWR _36205_/Q sky130_fd_sc_hd__dfxtp_1
X_21431_ _35627_/Q _34987_/Q _34347_/Q _33707_/Q _21391_/X _21392_/X VGND VGND VPWR
+ VPWR _21431_/X sky130_fd_sc_hd__mux4_1
X_33417_ _34121_/CLK _33417_/D VGND VGND VPWR VPWR _33417_/Q sky130_fd_sc_hd__dfxtp_1
X_30629_ _30740_/S VGND VGND VPWR VPWR _30648_/S sky130_fd_sc_hd__buf_4
XFILLER_72_1284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34397_ _36235_/CLK _34397_/D VGND VGND VPWR VPWR _34397_/Q sky130_fd_sc_hd__dfxtp_1
X_24150_ _24150_/A VGND VGND VPWR VPWR _32612_/D sky130_fd_sc_hd__clkbuf_1
X_33348_ _34177_/CLK _33348_/D VGND VGND VPWR VPWR _33348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21362_ _34665_/Q _34601_/Q _34537_/Q _34473_/Q _21186_/X _21187_/X VGND VGND VPWR
+ VPWR _21362_/X sky130_fd_sc_hd__mux4_1
X_36136_ _36136_/CLK _36136_/D VGND VGND VPWR VPWR _36136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20313_ _33933_/Q _33869_/Q _33805_/Q _36109_/Q _20030_/X _20031_/X VGND VGND VPWR
+ VPWR _20313_/X sky130_fd_sc_hd__mux4_1
X_23101_ _23101_/A VGND VGND VPWR VPWR _32090_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24081_ _24081_/A VGND VGND VPWR VPWR _32581_/D sky130_fd_sc_hd__clkbuf_1
Xinput80 R3[3] VGND VGND VPWR VPWR input80/X sky130_fd_sc_hd__buf_4
X_33279_ _35648_/CLK _33279_/D VGND VGND VPWR VPWR _33279_/Q sky130_fd_sc_hd__dfxtp_1
X_36067_ _36070_/CLK _36067_/D VGND VGND VPWR VPWR _36067_/Q sky130_fd_sc_hd__dfxtp_1
X_21293_ _34407_/Q _36135_/Q _34279_/Q _34215_/Q _21123_/X _21124_/X VGND VGND VPWR
+ VPWR _21293_/X sky130_fd_sc_hd__mux4_1
XFILLER_200_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23032_ _23032_/A VGND VGND VPWR VPWR _32068_/D sky130_fd_sc_hd__clkbuf_1
X_20244_ _34187_/Q _34123_/Q _34059_/Q _33995_/Q _20099_/X _20100_/X VGND VGND VPWR
+ VPWR _20244_/X sky130_fd_sc_hd__mux4_1
X_35018_ _35724_/CLK _35018_/D VGND VGND VPWR VPWR _35018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_946 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_646 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27840_ _27840_/A _31823_/B VGND VGND VPWR VPWR _27973_/S sky130_fd_sc_hd__nand2_8
X_20175_ _33673_/Q _33609_/Q _33545_/Q _33481_/Q _19853_/X _19854_/X VGND VGND VPWR
+ VPWR _20175_/X sky130_fd_sc_hd__mux4_1
XFILLER_192_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27771_ _27770_/X _34239_/Q _27795_/S VGND VGND VPWR VPWR _27772_/A sky130_fd_sc_hd__mux2_1
XTAP_4405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24983_ _24982_/X _32977_/Q _24983_/S VGND VGND VPWR VPWR _24984_/A sky130_fd_sc_hd__mux2_1
XTAP_4416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29510_ _35024_/Q _29509_/X _29513_/S VGND VGND VPWR VPWR _29511_/A sky130_fd_sc_hd__mux2_1
XTAP_4427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26722_ _33794_/Q _23435_/X _26732_/S VGND VGND VPWR VPWR _26723_/A sky130_fd_sc_hd__mux2_1
XTAP_4438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23934_ _23018_/X _32512_/Q _23948_/S VGND VGND VPWR VPWR _23935_/A sky130_fd_sc_hd__mux2_1
XTAP_3704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29441_ input30/X VGND VGND VPWR VPWR _29441_/X sky130_fd_sc_hd__buf_2
XTAP_3748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26653_ _33761_/Q _23265_/X _26669_/S VGND VGND VPWR VPWR _26654_/A sky130_fd_sc_hd__mux2_1
XFILLER_217_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23865_ _23865_/A VGND VGND VPWR VPWR _32479_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25604_ _24889_/X _33267_/Q _25604_/S VGND VGND VPWR VPWR _25605_/A sky130_fd_sc_hd__mux2_1
XFILLER_246_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22816_ _22812_/X _22815_/X _22471_/A VGND VGND VPWR VPWR _22817_/D sky130_fd_sc_hd__o21ba_1
X_29372_ _29372_/A VGND VGND VPWR VPWR _34979_/D sky130_fd_sc_hd__clkbuf_1
X_26584_ _26584_/A VGND VGND VPWR VPWR _33730_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23796_ _23796_/A VGND VGND VPWR VPWR _32383_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28323_ _28323_/A VGND VGND VPWR VPWR _34490_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_246_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25535_ _25535_/A VGND VGND VPWR VPWR _33234_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22747_ _33105_/Q _32081_/Q _35857_/Q _35793_/Q _20679_/X _20680_/X VGND VGND VPWR
+ VPWR _22747_/X sky130_fd_sc_hd__mux4_1
XFILLER_13_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28254_ _28254_/A VGND VGND VPWR VPWR _34457_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25466_ _25466_/A VGND VGND VPWR VPWR _33201_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22678_ _22365_/X _22676_/X _22677_/X _22371_/X VGND VGND VPWR VPWR _22678_/X sky130_fd_sc_hd__a22o_1
XFILLER_51_1302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27205_ input51/X VGND VGND VPWR VPWR _27205_/X sky130_fd_sc_hd__buf_4
X_24417_ _24417_/A VGND VGND VPWR VPWR _32737_/D sky130_fd_sc_hd__clkbuf_1
X_28185_ _27751_/X _34425_/Q _28193_/S VGND VGND VPWR VPWR _28186_/A sky130_fd_sc_hd__mux2_1
X_21629_ _32625_/Q _32561_/Q _32497_/Q _35953_/Q _21523_/X _21307_/X VGND VGND VPWR
+ VPWR _21629_/X sky130_fd_sc_hd__mux4_1
X_25397_ _33170_/Q _23487_/X _25403_/S VGND VGND VPWR VPWR _25398_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27136_ _27136_/A VGND VGND VPWR VPWR _33974_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24348_ _23021_/X _32705_/Q _24360_/S VGND VGND VPWR VPWR _24349_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27067_ _33952_/Q _27065_/X _27094_/S VGND VGND VPWR VPWR _27068_/A sky130_fd_sc_hd__mux2_1
X_24279_ _22918_/X _32672_/Q _24297_/S VGND VGND VPWR VPWR _24280_/A sky130_fd_sc_hd__mux2_1
XFILLER_181_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_5_21_0_CLK clkbuf_2_2_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_21_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_49_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26018_ _24902_/X _33463_/Q _26030_/S VGND VGND VPWR VPWR _26019_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18840_ _18653_/X _18838_/X _18839_/X _18659_/X VGND VGND VPWR VPWR _18840_/X sky130_fd_sc_hd__a22o_1
XTAP_7075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18771_ _33121_/Q _36001_/Q _32993_/Q _32929_/Q _18656_/X _18657_/X VGND VGND VPWR
+ VPWR _18771_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27969_ _27831_/X _34323_/Q _27973_/S VGND VGND VPWR VPWR _27970_/A sky130_fd_sc_hd__mux2_1
XTAP_5640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15983_ _16061_/A VGND VGND VPWR VPWR _17906_/A sky130_fd_sc_hd__buf_12
XTAP_6385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17722_ _17511_/X _17720_/X _17721_/X _17516_/X VGND VGND VPWR VPWR _17722_/X sky130_fd_sc_hd__a22o_1
XTAP_5662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29708_ _35115_/Q _29395_/X _29724_/S VGND VGND VPWR VPWR _29709_/A sky130_fd_sc_hd__mux2_1
XTAP_5684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30980_ _30980_/A VGND VGND VPWR VPWR _35718_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17653_ _17649_/X _17652_/X _17518_/X VGND VGND VPWR VPWR _17654_/D sky130_fd_sc_hd__o21ba_1
XTAP_4972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29639_ _29639_/A VGND VGND VPWR VPWR _35082_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16604_ _32613_/Q _32549_/Q _32485_/Q _35941_/Q _16570_/X _16354_/X VGND VGND VPWR
+ VPWR _16604_/X sky130_fd_sc_hd__mux4_1
X_32650_ _36040_/CLK _32650_/D VGND VGND VPWR VPWR _32650_/Q sky130_fd_sc_hd__dfxtp_1
X_17584_ _34432_/Q _36160_/Q _34304_/Q _34240_/Q _17582_/X _17583_/X VGND VGND VPWR
+ VPWR _17584_/X sky130_fd_sc_hd__mux4_1
XFILLER_51_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19323_ _33393_/Q _33329_/Q _33265_/Q _33201_/Q _19074_/X _19075_/X VGND VGND VPWR
+ VPWR _19323_/X sky130_fd_sc_hd__mux4_1
X_31601_ _27711_/X _36012_/Q _31615_/S VGND VGND VPWR VPWR _31602_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_1390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16535_ _33891_/Q _33827_/Q _33763_/Q _36067_/Q _16318_/X _16319_/X VGND VGND VPWR
+ VPWR _16535_/X sky130_fd_sc_hd__mux4_1
X_32581_ _35907_/CLK _32581_/D VGND VGND VPWR VPWR _32581_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34320_ _36176_/CLK _34320_/D VGND VGND VPWR VPWR _34320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31532_ _31532_/A VGND VGND VPWR VPWR _35979_/D sky130_fd_sc_hd__clkbuf_1
X_19254_ _33903_/Q _33839_/Q _33775_/Q _36079_/Q _18971_/X _18972_/X VGND VGND VPWR
+ VPWR _19254_/X sky130_fd_sc_hd__mux4_1
XFILLER_204_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16466_ _33377_/Q _33313_/Q _33249_/Q _33185_/Q _16421_/X _16422_/X VGND VGND VPWR
+ VPWR _16466_/X sky130_fd_sc_hd__mux4_1
XFILLER_32_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18205_ _15981_/X _18203_/X _18204_/X _15991_/X VGND VGND VPWR VPWR _18205_/X sky130_fd_sc_hd__a22o_1
X_34251_ _36173_/CLK _34251_/D VGND VGND VPWR VPWR _34251_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19185_ _34157_/Q _34093_/Q _34029_/Q _33965_/Q _19040_/X _19041_/X VGND VGND VPWR
+ VPWR _19185_/X sky130_fd_sc_hd__mux4_1
X_31463_ _31463_/A VGND VGND VPWR VPWR _35946_/D sky130_fd_sc_hd__clkbuf_1
X_16397_ _16353_/X _16395_/X _16396_/X _16359_/X VGND VGND VPWR VPWR _16397_/X sky130_fd_sc_hd__a22o_1
X_33202_ _33393_/CLK _33202_/D VGND VGND VPWR VPWR _33202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_982 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18136_ _32657_/Q _32593_/Q _32529_/Q _35985_/Q _17982_/X _16877_/A VGND VGND VPWR
+ VPWR _18136_/X sky130_fd_sc_hd__mux4_1
X_30414_ _35450_/Q _29441_/X _30420_/S VGND VGND VPWR VPWR _30415_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_1022 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34182_ _34182_/CLK _34182_/D VGND VGND VPWR VPWR _34182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31394_ _27804_/X _35914_/Q _31408_/S VGND VGND VPWR VPWR _31395_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33133_ _36013_/CLK _33133_/D VGND VGND VPWR VPWR _33133_/Q sky130_fd_sc_hd__dfxtp_1
X_30345_ _35417_/Q _29339_/X _30357_/S VGND VGND VPWR VPWR _30346_/A sky130_fd_sc_hd__mux2_1
X_18067_ _18067_/A _18067_/B _18067_/C _18067_/D VGND VGND VPWR VPWR _18068_/A sky130_fd_sc_hd__or4_2
XFILLER_160_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17018_ _17018_/A _17018_/B _17018_/C _17018_/D VGND VGND VPWR VPWR _17019_/A sky130_fd_sc_hd__or4_4
XFILLER_67_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33064_ _35755_/CLK _33064_/D VGND VGND VPWR VPWR _33064_/Q sky130_fd_sc_hd__dfxtp_1
X_30276_ _30276_/A VGND VGND VPWR VPWR _35384_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32015_ _36202_/CLK _32015_/D VGND VGND VPWR VPWR _32015_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18969_ _18793_/X _18967_/X _18968_/X _18798_/X VGND VGND VPWR VPWR _18969_/X sky130_fd_sc_hd__a22o_1
XFILLER_246_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_1391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33966_ _35630_/CLK _33966_/D VGND VGND VPWR VPWR _33966_/Q sky130_fd_sc_hd__dfxtp_1
X_21980_ _21806_/X _21976_/X _21979_/X _21809_/X VGND VGND VPWR VPWR _21980_/X sky130_fd_sc_hd__a22o_1
XFILLER_187_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35705_ _35835_/CLK _35705_/D VGND VGND VPWR VPWR _35705_/Q sky130_fd_sc_hd__dfxtp_1
X_20931_ _35613_/Q _34973_/Q _34333_/Q _33693_/Q _20653_/X _20655_/X VGND VGND VPWR
+ VPWR _20931_/X sky130_fd_sc_hd__mux4_1
X_32917_ _35989_/CLK _32917_/D VGND VGND VPWR VPWR _32917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_214_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33897_ _33897_/CLK _33897_/D VGND VGND VPWR VPWR _33897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20862_ _20648_/X _20860_/X _20861_/X _20658_/X VGND VGND VPWR VPWR _20862_/X sky130_fd_sc_hd__a22o_1
X_35636_ _35701_/CLK _35636_/D VGND VGND VPWR VPWR _35636_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23650_ _23005_/X _32316_/Q _23652_/S VGND VGND VPWR VPWR _23651_/A sky130_fd_sc_hd__mux2_1
X_32848_ _32914_/CLK _32848_/D VGND VGND VPWR VPWR _32848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22601_ _35212_/Q _35148_/Q _35084_/Q _32268_/Q _22316_/X _22317_/X VGND VGND VPWR
+ VPWR _22601_/X sky130_fd_sc_hd__mux4_1
XFILLER_240_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20793_ _35609_/Q _34969_/Q _34329_/Q _33689_/Q _20653_/X _20655_/X VGND VGND VPWR
+ VPWR _20793_/X sky130_fd_sc_hd__mux4_1
X_23581_ _22903_/X _32283_/Q _23589_/S VGND VGND VPWR VPWR _23582_/A sky130_fd_sc_hd__mux2_1
X_35567_ _35567_/CLK _35567_/D VGND VGND VPWR VPWR _35567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32779_ _32907_/CLK _32779_/D VGND VGND VPWR VPWR _32779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25320_ _33133_/Q _23302_/X _25332_/S VGND VGND VPWR VPWR _25321_/A sky130_fd_sc_hd__mux2_1
X_34518_ _34647_/CLK _34518_/D VGND VGND VPWR VPWR _34518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22532_ _34698_/Q _34634_/Q _34570_/Q _34506_/Q _22245_/X _22246_/X VGND VGND VPWR
+ VPWR _22532_/X sky130_fd_sc_hd__mux4_1
XFILLER_210_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35498_ _35690_/CLK _35498_/D VGND VGND VPWR VPWR _35498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25251_ _33101_/Q _23472_/X _25259_/S VGND VGND VPWR VPWR _25252_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34449_ _36175_/CLK _34449_/D VGND VGND VPWR VPWR _34449_/Q sky130_fd_sc_hd__dfxtp_1
X_22463_ _22459_/X _22460_/X _22461_/X _22462_/X VGND VGND VPWR VPWR _22463_/X sky130_fd_sc_hd__a22o_1
XFILLER_33_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24202_ _24202_/A VGND VGND VPWR VPWR _32637_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21414_ _21414_/A _21414_/B _21414_/C _21414_/D VGND VGND VPWR VPWR _21415_/A sky130_fd_sc_hd__or4_4
X_22394_ _22111_/X _22392_/X _22393_/X _22116_/X VGND VGND VPWR VPWR _22394_/X sky130_fd_sc_hd__a22o_1
X_25182_ _33068_/Q _23299_/X _25196_/S VGND VGND VPWR VPWR _25183_/A sky130_fd_sc_hd__mux2_1
XFILLER_136_835 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36119_ _36119_/CLK _36119_/D VGND VGND VPWR VPWR _36119_/Q sky130_fd_sc_hd__dfxtp_1
X_24133_ _24133_/A VGND VGND VPWR VPWR _32604_/D sky130_fd_sc_hd__clkbuf_1
X_21345_ _33897_/Q _33833_/Q _33769_/Q _36073_/Q _21271_/X _21272_/X VGND VGND VPWR
+ VPWR _21345_/X sky130_fd_sc_hd__mux4_1
XFILLER_198_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29990_ _35249_/Q _29413_/X _29994_/S VGND VGND VPWR VPWR _29991_/A sky130_fd_sc_hd__mux2_1
XFILLER_191_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28941_ _34782_/Q _27059_/X _28943_/S VGND VGND VPWR VPWR _28942_/A sky130_fd_sc_hd__mux2_1
X_21276_ _32615_/Q _32551_/Q _32487_/Q _35943_/Q _21170_/X _20954_/X VGND VGND VPWR
+ VPWR _21276_/X sky130_fd_sc_hd__mux4_1
X_24064_ _24064_/A VGND VGND VPWR VPWR _32573_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20227_ _20004_/X _20225_/X _20226_/X _20007_/X VGND VGND VPWR VPWR _20227_/X sky130_fd_sc_hd__a22o_1
X_23015_ input36/X VGND VGND VPWR VPWR _23015_/X sky130_fd_sc_hd__clkbuf_2
X_28872_ _28872_/A VGND VGND VPWR VPWR _34749_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27823_ _27822_/X _34256_/Q _27826_/S VGND VGND VPWR VPWR _27824_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20158_ _20153_/X _20156_/X _20157_/X VGND VGND VPWR VPWR _20173_/C sky130_fd_sc_hd__o21ba_1
XFILLER_77_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27754_ input30/X VGND VGND VPWR VPWR _27754_/X sky130_fd_sc_hd__buf_2
X_20089_ _34694_/Q _34630_/Q _34566_/Q _34502_/Q _19945_/X _19946_/X VGND VGND VPWR
+ VPWR _20089_/X sky130_fd_sc_hd__mux4_1
X_24966_ _24966_/A VGND VGND VPWR VPWR _32971_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26705_ _33786_/Q _23408_/X _26711_/S VGND VGND VPWR VPWR _26706_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23917_ _22993_/X _32504_/Q _23927_/S VGND VGND VPWR VPWR _23918_/A sky130_fd_sc_hd__mux2_1
XFILLER_206_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27685_ _27685_/A VGND VGND VPWR VPWR _34211_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24897_ _24896_/X _32949_/Q _24921_/S VGND VGND VPWR VPWR _24898_/A sky130_fd_sc_hd__mux2_1
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29424_ _34996_/Q _29422_/X _29451_/S VGND VGND VPWR VPWR _29425_/A sky130_fd_sc_hd__mux2_1
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26636_ _33753_/Q _23240_/X _26648_/S VGND VGND VPWR VPWR _26637_/A sky130_fd_sc_hd__mux2_1
XTAP_3578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23848_ _22891_/X _32471_/Q _23864_/S VGND VGND VPWR VPWR _23849_/A sky130_fd_sc_hd__mux2_1
XTAP_3589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29355_ _34974_/Q _29354_/X _29358_/S VGND VGND VPWR VPWR _29356_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_782 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26567_ _26567_/A VGND VGND VPWR VPWR _33722_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23779_ _23779_/A VGND VGND VPWR VPWR _32375_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16320_ _33885_/Q _33821_/Q _33757_/Q _36061_/Q _16318_/X _16319_/X VGND VGND VPWR
+ VPWR _16320_/X sky130_fd_sc_hd__mux4_1
X_28306_ _28306_/A VGND VGND VPWR VPWR _34482_/D sky130_fd_sc_hd__clkbuf_1
X_25518_ _24961_/X _33226_/Q _25532_/S VGND VGND VPWR VPWR _25519_/A sky130_fd_sc_hd__mux2_1
X_29286_ _29286_/A VGND VGND VPWR VPWR _34945_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26498_ _26498_/A VGND VGND VPWR VPWR _33689_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28237_ _27828_/X _34450_/Q _28243_/S VGND VGND VPWR VPWR _28238_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16251_ _32603_/Q _32539_/Q _32475_/Q _35931_/Q _16217_/X _17717_/A VGND VGND VPWR
+ VPWR _16251_/X sky130_fd_sc_hd__mux4_1
X_25449_ _25449_/A VGND VGND VPWR VPWR _33193_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16182_ _33881_/Q _33817_/Q _33753_/Q _36057_/Q _16112_/X _16113_/X VGND VGND VPWR
+ VPWR _16182_/X sky130_fd_sc_hd__mux4_1
X_28168_ _27726_/X _34417_/Q _28172_/S VGND VGND VPWR VPWR _28169_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27119_ _33969_/Q _27118_/X _27125_/S VGND VGND VPWR VPWR _27120_/A sky130_fd_sc_hd__mux2_1
X_28099_ _28099_/A VGND VGND VPWR VPWR _34384_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30130_ _30130_/A VGND VGND VPWR VPWR _35315_/D sky130_fd_sc_hd__clkbuf_1
X_19941_ _35458_/Q _35394_/Q _35330_/Q _35266_/Q _19907_/X _19908_/X VGND VGND VPWR
+ VPWR _19941_/X sky130_fd_sc_hd__mux4_1
XFILLER_141_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_218_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30061_ _35283_/Q _29518_/X _30065_/S VGND VGND VPWR VPWR _30062_/A sky130_fd_sc_hd__mux2_1
X_19872_ _35712_/Q _32222_/Q _35584_/Q _35520_/Q _19617_/X _19618_/X VGND VGND VPWR
+ VPWR _19872_/X sky130_fd_sc_hd__mux4_1
XFILLER_4_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18823_ _20016_/A VGND VGND VPWR VPWR _18823_/X sky130_fd_sc_hd__buf_6
XFILLER_228_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33820_ _36058_/CLK _33820_/D VGND VGND VPWR VPWR _33820_/Q sky130_fd_sc_hd__dfxtp_1
X_18754_ _20166_/A VGND VGND VPWR VPWR _18754_/X sky130_fd_sc_hd__buf_4
XTAP_5470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17705_ _35716_/Q _32226_/Q _35588_/Q _35524_/Q _17670_/X _17671_/X VGND VGND VPWR
+ VPWR _17705_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33751_ _36059_/CLK _33751_/D VGND VGND VPWR VPWR _33751_/Q sky130_fd_sc_hd__dfxtp_1
X_30963_ _35710_/Q input35/X _30981_/S VGND VGND VPWR VPWR _30964_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18685_ _18685_/A VGND VGND VPWR VPWR _32414_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32702_ _32894_/CLK _32702_/D VGND VGND VPWR VPWR _32702_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17636_ _17420_/X _17634_/X _17635_/X _17424_/X VGND VGND VPWR VPWR _17636_/X sky130_fd_sc_hd__a22o_1
X_33682_ _33875_/CLK _33682_/D VGND VGND VPWR VPWR _33682_/Q sky130_fd_sc_hd__dfxtp_1
X_30894_ _30894_/A VGND VGND VPWR VPWR _35677_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_224_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35421_ _35805_/CLK _35421_/D VGND VGND VPWR VPWR _35421_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17567_ _17412_/X _17565_/X _17566_/X _17418_/X VGND VGND VPWR VPWR _17567_/X sky130_fd_sc_hd__a22o_1
X_32633_ _36025_/CLK _32633_/D VGND VGND VPWR VPWR _32633_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19306_ _20169_/A VGND VGND VPWR VPWR _19306_/X sky130_fd_sc_hd__clkbuf_4
X_16518_ _16297_/X _16516_/X _16517_/X _16300_/X VGND VGND VPWR VPWR _16518_/X sky130_fd_sc_hd__a22o_1
X_35352_ _35799_/CLK _35352_/D VGND VGND VPWR VPWR _35352_/Q sky130_fd_sc_hd__dfxtp_1
X_32564_ _35956_/CLK _32564_/D VGND VGND VPWR VPWR _32564_/Q sky130_fd_sc_hd__dfxtp_1
X_17498_ _17851_/A VGND VGND VPWR VPWR _17498_/X sky130_fd_sc_hd__buf_4
XFILLER_182_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34303_ _36103_/CLK _34303_/D VGND VGND VPWR VPWR _34303_/Q sky130_fd_sc_hd__dfxtp_1
X_31515_ _31515_/A VGND VGND VPWR VPWR _35971_/D sky130_fd_sc_hd__clkbuf_1
X_19237_ _18950_/X _19235_/X _19236_/X _18953_/X VGND VGND VPWR VPWR _19237_/X sky130_fd_sc_hd__a22o_1
X_16449_ _35168_/Q _35104_/Q _35040_/Q _32160_/Q _16304_/X _16305_/X VGND VGND VPWR
+ VPWR _16449_/X sky130_fd_sc_hd__mux4_1
X_35283_ _35666_/CLK _35283_/D VGND VGND VPWR VPWR _35283_/Q sky130_fd_sc_hd__dfxtp_1
X_32495_ _35951_/CLK _32495_/D VGND VGND VPWR VPWR _32495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31446_ _31446_/A VGND VGND VPWR VPWR _35938_/D sky130_fd_sc_hd__clkbuf_1
X_19168_ _18945_/X _19166_/X _19167_/X _18948_/X VGND VGND VPWR VPWR _19168_/X sky130_fd_sc_hd__a22o_1
X_34234_ _36153_/CLK _34234_/D VGND VGND VPWR VPWR _34234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18119_ _18115_/X _18118_/X _17857_/X VGND VGND VPWR VPWR _18127_/C sky130_fd_sc_hd__o21ba_1
XFILLER_118_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34165_ _35703_/CLK _34165_/D VGND VGND VPWR VPWR _34165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31377_ _27779_/X _35906_/Q _31387_/S VGND VGND VPWR VPWR _31378_/A sky130_fd_sc_hd__mux2_1
X_19099_ _19094_/X _19097_/X _19098_/X VGND VGND VPWR VPWR _19114_/C sky130_fd_sc_hd__o21ba_1
XFILLER_133_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21130_ _21130_/A VGND VGND VPWR VPWR _36194_/D sky130_fd_sc_hd__clkbuf_1
X_30328_ _30328_/A VGND VGND VPWR VPWR _35409_/D sky130_fd_sc_hd__clkbuf_1
X_33116_ _36054_/CLK _33116_/D VGND VGND VPWR VPWR _33116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34096_ _35632_/CLK _34096_/D VGND VGND VPWR VPWR _34096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_890 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33047_ _36118_/CLK _33047_/D VGND VGND VPWR VPWR _33047_/Q sky130_fd_sc_hd__dfxtp_1
X_21061_ _21061_/A _21061_/B _21061_/C _21061_/D VGND VGND VPWR VPWR _21062_/A sky130_fd_sc_hd__or4_1
X_30259_ _30259_/A VGND VGND VPWR VPWR _35376_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20012_ _20169_/A VGND VGND VPWR VPWR _20012_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_113_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24820_ _24820_/A VGND VGND VPWR VPWR _32924_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_230_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34998_ _35768_/CLK _34998_/D VGND VGND VPWR VPWR _34998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24751_ _23018_/X _32896_/Q _24765_/S VGND VGND VPWR VPWR _24752_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33949_ _36188_/CLK _33949_/D VGND VGND VPWR VPWR _33949_/Q sky130_fd_sc_hd__dfxtp_1
X_21963_ _22316_/A VGND VGND VPWR VPWR _21963_/X sky130_fd_sc_hd__buf_6
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23702_ _23082_/X _32341_/Q _23702_/S VGND VGND VPWR VPWR _23703_/A sky130_fd_sc_hd__mux2_1
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27470_ _27470_/A VGND VGND VPWR VPWR _34117_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_199_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20914_ _33629_/Q _33565_/Q _33501_/Q _33437_/Q _20741_/X _20742_/X VGND VGND VPWR
+ VPWR _20914_/X sky130_fd_sc_hd__mux4_1
X_24682_ _24682_/A VGND VGND VPWR VPWR _32863_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21894_ _34680_/Q _34616_/Q _34552_/Q _34488_/Q _21892_/X _21893_/X VGND VGND VPWR
+ VPWR _21894_/X sky130_fd_sc_hd__mux4_1
XFILLER_82_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_243_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26421_ _26421_/A VGND VGND VPWR VPWR _33653_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23633_ _23702_/S VGND VGND VPWR VPWR _23652_/S sky130_fd_sc_hd__buf_4
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35619_ _35620_/CLK _35619_/D VGND VGND VPWR VPWR _35619_/Q sky130_fd_sc_hd__dfxtp_1
X_20845_ _34139_/Q _34075_/Q _34011_/Q _33947_/Q _20609_/X _20611_/X VGND VGND VPWR
+ VPWR _20845_/X sky130_fd_sc_hd__mux4_1
X_29140_ _29140_/A VGND VGND VPWR VPWR _34876_/D sky130_fd_sc_hd__clkbuf_1
X_26352_ _30877_/B _26352_/B VGND VGND VPWR VPWR _26353_/A sky130_fd_sc_hd__and2b_1
X_23564_ _23564_/A VGND VGND VPWR VPWR _32276_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20776_ _20776_/A _20776_/B _20776_/C _20776_/D VGND VGND VPWR VPWR _20777_/A sky130_fd_sc_hd__or4_1
XFILLER_195_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25303_ _33125_/Q _23277_/X _25311_/S VGND VGND VPWR VPWR _25304_/A sky130_fd_sc_hd__mux2_1
X_29071_ _29071_/A VGND VGND VPWR VPWR _34843_/D sky130_fd_sc_hd__clkbuf_1
X_22515_ _22515_/A VGND VGND VPWR VPWR _22515_/X sky130_fd_sc_hd__clkbuf_4
X_26283_ _26283_/A VGND VGND VPWR VPWR _33588_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23495_ input59/X VGND VGND VPWR VPWR _23495_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_211_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28022_ _28022_/A VGND VGND VPWR VPWR _34347_/D sky130_fd_sc_hd__clkbuf_1
X_25234_ _33093_/Q _23444_/X _25238_/S VGND VGND VPWR VPWR _25235_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22446_ _22446_/A VGND VGND VPWR VPWR _22446_/X sky130_fd_sc_hd__buf_2
XFILLER_52_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25165_ _33060_/Q _23274_/X _25175_/S VGND VGND VPWR VPWR _25166_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22377_ _22377_/A VGND VGND VPWR VPWR _22377_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_129_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24116_ input85/X input84/X _27232_/A VGND VGND VPWR VPWR _24117_/A sky130_fd_sc_hd__or3_1
XFILLER_135_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21328_ _21250_/X _21324_/X _21327_/X _21253_/X VGND VGND VPWR VPWR _21328_/X sky130_fd_sc_hd__a22o_1
X_25096_ _25096_/A VGND VGND VPWR VPWR _33028_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29973_ _35241_/Q _29388_/X _29973_/S VGND VGND VPWR VPWR _29974_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28924_ _29056_/S VGND VGND VPWR VPWR _28943_/S sky130_fd_sc_hd__buf_4
X_21259_ _35174_/Q _35110_/Q _35046_/Q _32166_/Q _21257_/X _21258_/X VGND VGND VPWR
+ VPWR _21259_/X sky130_fd_sc_hd__mux4_1
X_24047_ _22984_/X _32565_/Q _24063_/S VGND VGND VPWR VPWR _24048_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28855_ _34741_/Q _27131_/X _28871_/S VGND VGND VPWR VPWR _28856_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27806_ _27806_/A VGND VGND VPWR VPWR _34250_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28786_ _28786_/A _28786_/B VGND VGND VPWR VPWR _28787_/A sky130_fd_sc_hd__or2_1
XTAP_4021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25998_ _25998_/A VGND VGND VPWR VPWR _33453_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27737_ _27735_/X _34228_/Q _27764_/S VGND VGND VPWR VPWR _27738_/A sky130_fd_sc_hd__mux2_1
XTAP_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24949_ _24948_/X _32966_/Q _24952_/S VGND VGND VPWR VPWR _24950_/A sky130_fd_sc_hd__mux2_1
XTAP_4065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18470_ _20016_/A VGND VGND VPWR VPWR _18470_/X sky130_fd_sc_hd__buf_6
XFILLER_79_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27668_ _27667_/X _34206_/Q _27671_/S VGND VGND VPWR VPWR _27669_/A sky130_fd_sc_hd__mux2_1
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17421_ _17774_/A VGND VGND VPWR VPWR _17421_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26619_ _26619_/A VGND VGND VPWR VPWR _33747_/D sky130_fd_sc_hd__clkbuf_1
X_29407_ input18/X VGND VGND VPWR VPWR _29407_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27599_ _27599_/A VGND VGND VPWR VPWR _34178_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17352_ _35706_/Q _32215_/Q _35578_/Q _35514_/Q _17317_/X _17318_/X VGND VGND VPWR
+ VPWR _17352_/X sky130_fd_sc_hd__mux4_1
X_29338_ _29338_/A VGND VGND VPWR VPWR _34968_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16303_ _34652_/Q _34588_/Q _34524_/Q _34460_/Q _16233_/X _16234_/X VGND VGND VPWR
+ VPWR _16303_/X sky130_fd_sc_hd__mux4_1
XFILLER_144_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29269_ _29269_/A VGND VGND VPWR VPWR _34937_/D sky130_fd_sc_hd__clkbuf_1
X_17283_ _17067_/X _17281_/X _17282_/X _17071_/X VGND VGND VPWR VPWR _17283_/X sky130_fd_sc_hd__a22o_1
XFILLER_220_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31300_ _31300_/A VGND VGND VPWR VPWR _35869_/D sky130_fd_sc_hd__clkbuf_1
X_19022_ _35624_/Q _34984_/Q _34344_/Q _33704_/Q _18738_/X _18739_/X VGND VGND VPWR
+ VPWR _19022_/X sky130_fd_sc_hd__mux4_1
X_16234_ _17999_/A VGND VGND VPWR VPWR _16234_/X sky130_fd_sc_hd__buf_6
XFILLER_16_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32280_ _32856_/CLK _32280_/D VGND VGND VPWR VPWR _32280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31231_ _27763_/X _35837_/Q _31231_/S VGND VGND VPWR VPWR _31232_/A sky130_fd_sc_hd__mux2_1
X_16165_ _16060_/X _16163_/X _16164_/X _16072_/X VGND VGND VPWR VPWR _16165_/X sky130_fd_sc_hd__a22o_1
XFILLER_86_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1074 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31162_ _27661_/X _35804_/Q _31168_/S VGND VGND VPWR VPWR _31163_/A sky130_fd_sc_hd__mux2_1
X_16096_ _17866_/A VGND VGND VPWR VPWR _16096_/X sky130_fd_sc_hd__buf_4
XFILLER_115_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30113_ _35307_/Q _29395_/X _30129_/S VGND VGND VPWR VPWR _30114_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19924_ _19852_/X _19922_/X _19923_/X _19857_/X VGND VGND VPWR VPWR _19924_/X sky130_fd_sc_hd__a22o_1
XFILLER_114_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35970_ _35970_/CLK _35970_/D VGND VGND VPWR VPWR _35970_/Q sky130_fd_sc_hd__dfxtp_1
X_31093_ _35772_/Q input32/X _31095_/S VGND VGND VPWR VPWR _31094_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30044_ _30044_/A VGND VGND VPWR VPWR _35274_/D sky130_fd_sc_hd__clkbuf_1
X_34921_ _34921_/CLK _34921_/D VGND VGND VPWR VPWR _34921_/Q sky130_fd_sc_hd__dfxtp_1
X_19855_ _33664_/Q _33600_/Q _33536_/Q _33472_/Q _19853_/X _19854_/X VGND VGND VPWR
+ VPWR _19855_/X sky130_fd_sc_hd__mux4_1
XFILLER_150_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18806_ _32610_/Q _32546_/Q _32482_/Q _35938_/Q _18517_/X _18654_/X VGND VGND VPWR
+ VPWR _18806_/X sky130_fd_sc_hd__mux4_1
XFILLER_116_1468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34852_ _34918_/CLK _34852_/D VGND VGND VPWR VPWR _34852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19786_ _19779_/X _19784_/X _19785_/X VGND VGND VPWR VPWR _19820_/A sky130_fd_sc_hd__o21ba_1
X_16998_ _17859_/A VGND VGND VPWR VPWR _16998_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1042 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33803_ _36109_/CLK _33803_/D VGND VGND VPWR VPWR _33803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18737_ _35680_/Q _32186_/Q _35552_/Q _35488_/Q _18558_/X _18559_/X VGND VGND VPWR
+ VPWR _18737_/X sky130_fd_sc_hd__mux4_1
X_34783_ _34911_/CLK _34783_/D VGND VGND VPWR VPWR _34783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31995_ _34405_/CLK _31995_/D VGND VGND VPWR VPWR _31995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33734_ _35525_/CLK _33734_/D VGND VGND VPWR VPWR _33734_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18668_ _35678_/Q _32184_/Q _35550_/Q _35486_/Q _18558_/X _18559_/X VGND VGND VPWR
+ VPWR _18668_/X sky130_fd_sc_hd__mux4_1
X_30946_ _35702_/Q input26/X _30960_/S VGND VGND VPWR VPWR _30947_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17619_ _17615_/X _17618_/X _17518_/X VGND VGND VPWR VPWR _17620_/D sky130_fd_sc_hd__o21ba_1
X_33665_ _34180_/CLK _33665_/D VGND VGND VPWR VPWR _33665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30877_ _30877_/A _30877_/B VGND VGND VPWR VPWR _31010_/S sky130_fd_sc_hd__nor2_8
X_18599_ _33052_/Q _32028_/Q _35804_/Q _35740_/Q _18367_/X _18369_/X VGND VGND VPWR
+ VPWR _18599_/X sky130_fd_sc_hd__mux4_1
XFILLER_52_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35404_ _35596_/CLK _35404_/D VGND VGND VPWR VPWR _35404_/Q sky130_fd_sc_hd__dfxtp_1
X_20630_ _22512_/A VGND VGND VPWR VPWR _20630_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_71_1305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32616_ _35944_/CLK _32616_/D VGND VGND VPWR VPWR _32616_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33596_ _33661_/CLK _33596_/D VGND VGND VPWR VPWR _33596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35335_ _35463_/CLK _35335_/D VGND VGND VPWR VPWR _35335_/Q sky130_fd_sc_hd__dfxtp_1
X_20561_ _19458_/A _20559_/X _20560_/X _19463_/A VGND VGND VPWR VPWR _20561_/X sky130_fd_sc_hd__a22o_1
X_32547_ _35939_/CLK _32547_/D VGND VGND VPWR VPWR _32547_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22300_ _22434_/A VGND VGND VPWR VPWR _22300_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_149_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20492_ _33427_/Q _33363_/Q _33299_/Q _33235_/Q _18337_/X _18339_/X VGND VGND VPWR
+ VPWR _20492_/X sky130_fd_sc_hd__mux4_1
X_35266_ _35458_/CLK _35266_/D VGND VGND VPWR VPWR _35266_/Q sky130_fd_sc_hd__dfxtp_1
X_23280_ input8/X VGND VGND VPWR VPWR _23280_/X sky130_fd_sc_hd__buf_6
X_32478_ _35999_/CLK _32478_/D VGND VGND VPWR VPWR _32478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22231_ _33154_/Q _36034_/Q _33026_/Q _32962_/Q _22015_/X _22016_/X VGND VGND VPWR
+ VPWR _22231_/X sky130_fd_sc_hd__mux4_1
X_34217_ _35554_/CLK _34217_/D VGND VGND VPWR VPWR _34217_/Q sky130_fd_sc_hd__dfxtp_1
X_31429_ _31429_/A VGND VGND VPWR VPWR _35930_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35197_ _35197_/CLK _35197_/D VGND VGND VPWR VPWR _35197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22162_ _22515_/A VGND VGND VPWR VPWR _22162_/X sky130_fd_sc_hd__buf_4
X_34148_ _34148_/CLK _34148_/D VGND VGND VPWR VPWR _34148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21113_ _35682_/Q _32189_/Q _35554_/Q _35490_/Q _20858_/X _20859_/X VGND VGND VPWR
+ VPWR _21113_/X sky130_fd_sc_hd__mux4_1
XFILLER_82_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22093_ _22446_/A VGND VGND VPWR VPWR _22093_/X sky130_fd_sc_hd__clkbuf_4
X_26970_ _26970_/A VGND VGND VPWR VPWR _33911_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34079_ _36207_/CLK _34079_/D VGND VGND VPWR VPWR _34079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25921_ _24958_/X _33417_/Q _25937_/S VGND VGND VPWR VPWR _25922_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21044_ _20897_/X _21042_/X _21043_/X _20900_/X VGND VGND VPWR VPWR _21044_/X sky130_fd_sc_hd__a22o_1
XFILLER_114_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_247_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_755 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28640_ _27825_/X _34641_/Q _28640_/S VGND VGND VPWR VPWR _28641_/A sky130_fd_sc_hd__mux2_1
X_25852_ _25852_/A VGND VGND VPWR VPWR _33384_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_917 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24803_ input12/X VGND VGND VPWR VPWR _24803_/X sky130_fd_sc_hd__buf_2
XFILLER_46_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28571_ _27723_/X _34608_/Q _28577_/S VGND VGND VPWR VPWR _28572_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25783_ _25810_/S VGND VGND VPWR VPWR _25802_/S sky130_fd_sc_hd__buf_4
XFILLER_28_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22995_ _22995_/A VGND VGND VPWR VPWR _32056_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_216_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27522_ _34142_/Q _27059_/X _27524_/S VGND VGND VPWR VPWR _27523_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24734_ _22993_/X _32888_/Q _24744_/S VGND VGND VPWR VPWR _24735_/A sky130_fd_sc_hd__mux2_1
X_21946_ _22433_/A VGND VGND VPWR VPWR _21946_/X sky130_fd_sc_hd__buf_4
XFILLER_227_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_1366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27453_ _27453_/A VGND VGND VPWR VPWR _34109_/D sky130_fd_sc_hd__clkbuf_1
X_24665_ _22891_/X _32855_/Q _24681_/S VGND VGND VPWR VPWR _24666_/A sky130_fd_sc_hd__mux2_1
XFILLER_231_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21877_ _32632_/Q _32568_/Q _32504_/Q _35960_/Q _21876_/X _21660_/X VGND VGND VPWR
+ VPWR _21877_/X sky130_fd_sc_hd__mux4_1
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26404_ _26404_/A VGND VGND VPWR VPWR _33645_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23616_ _23616_/A VGND VGND VPWR VPWR _32299_/D sky130_fd_sc_hd__clkbuf_1
X_20828_ _20648_/X _20826_/X _20827_/X _20658_/X VGND VGND VPWR VPWR _20828_/X sky130_fd_sc_hd__a22o_1
X_27384_ _27384_/A VGND VGND VPWR VPWR _34076_/D sky130_fd_sc_hd__clkbuf_1
X_24596_ _24596_/A VGND VGND VPWR VPWR _32822_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_204_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29123_ _34868_/Q _27127_/X _29141_/S VGND VGND VPWR VPWR _29124_/A sky130_fd_sc_hd__mux2_1
X_26335_ _26335_/A VGND VGND VPWR VPWR _33613_/D sky130_fd_sc_hd__clkbuf_1
X_23547_ _32268_/Q _23469_/X _23557_/S VGND VGND VPWR VPWR _23548_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20759_ _20755_/X _20758_/X _20644_/X _20646_/X VGND VGND VPWR VPWR _20776_/B sky130_fd_sc_hd__o211a_1
XFILLER_126_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29054_ _34836_/Q _27226_/X _29056_/S VGND VGND VPWR VPWR _29055_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26266_ _26266_/A VGND VGND VPWR VPWR _33580_/D sky130_fd_sc_hd__clkbuf_1
X_23478_ input53/X VGND VGND VPWR VPWR _23478_/X sky130_fd_sc_hd__buf_4
XFILLER_137_930 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28005_ _28005_/A VGND VGND VPWR VPWR _34339_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25217_ _33085_/Q _23417_/X _25217_/S VGND VGND VPWR VPWR _25218_/A sky130_fd_sc_hd__mux2_1
X_22429_ _22429_/A VGND VGND VPWR VPWR _36231_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26197_ _24967_/X _33548_/Q _26207_/S VGND VGND VPWR VPWR _26198_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25148_ _33052_/Q _23249_/X _25154_/S VGND VGND VPWR VPWR _25149_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17970_ _34955_/Q _34891_/Q _34827_/Q _34763_/Q _17866_/X _17867_/X VGND VGND VPWR
+ VPWR _17970_/X sky130_fd_sc_hd__mux4_1
X_25079_ _25079_/A VGND VGND VPWR VPWR _33020_/D sky130_fd_sc_hd__clkbuf_1
X_29956_ _29956_/A VGND VGND VPWR VPWR _35232_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_219_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28907_ _34766_/Q _27208_/X _28913_/S VGND VGND VPWR VPWR _28908_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16921_ _16853_/X _16919_/X _16920_/X _16856_/X VGND VGND VPWR VPWR _16921_/X sky130_fd_sc_hd__a22o_1
XFILLER_105_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29887_ _35200_/Q _29460_/X _29901_/S VGND VGND VPWR VPWR _29888_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19640_ _19506_/X _19638_/X _19639_/X _19509_/X VGND VGND VPWR VPWR _19640_/X sky130_fd_sc_hd__a22o_1
X_16852_ _16846_/X _16849_/X _16850_/X _16851_/X VGND VGND VPWR VPWR _16852_/X sky130_fd_sc_hd__a22o_1
X_28838_ _34733_/Q _27106_/X _28850_/S VGND VGND VPWR VPWR _28839_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19571_ _19499_/X _19569_/X _19570_/X _19504_/X VGND VGND VPWR VPWR _19571_/X sky130_fd_sc_hd__a22o_1
X_16783_ _16706_/X _16781_/X _16782_/X _16712_/X VGND VGND VPWR VPWR _16783_/X sky130_fd_sc_hd__a22o_1
XFILLER_93_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28769_ _28769_/A VGND VGND VPWR VPWR _34701_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_58__f_CLK clkbuf_5_29_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_58__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_93_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18522_ _32090_/Q _32282_/Q _32346_/Q _35866_/Q _18521_/X _20167_/A VGND VGND VPWR
+ VPWR _18522_/X sky130_fd_sc_hd__mux4_1
X_30800_ _35633_/Q input20/X _30804_/S VGND VGND VPWR VPWR _30801_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31780_ _36097_/Q input38/X _31792_/S VGND VGND VPWR VPWR _31781_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_1248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_786 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18453_ _32600_/Q _32536_/Q _32472_/Q _35928_/Q _20166_/A _20017_/A VGND VGND VPWR
+ VPWR _18453_/X sky130_fd_sc_hd__mux4_1
XFILLER_206_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30731_ _30731_/A VGND VGND VPWR VPWR _35600_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17404_ _17404_/A VGND VGND VPWR VPWR _31995_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18384_ _20066_/A VGND VGND VPWR VPWR _19311_/A sky130_fd_sc_hd__buf_12
X_33450_ _35690_/CLK _33450_/D VGND VGND VPWR VPWR _33450_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30662_ _30662_/A VGND VGND VPWR VPWR _35567_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32401_ _35921_/CLK _32401_/D VGND VGND VPWR VPWR _32401_/Q sky130_fd_sc_hd__dfxtp_1
X_17335_ _33658_/Q _33594_/Q _33530_/Q _33466_/Q _17200_/X _17201_/X VGND VGND VPWR
+ VPWR _17335_/X sky130_fd_sc_hd__mux4_1
XFILLER_14_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30593_ _35535_/Q _29506_/X _30597_/S VGND VGND VPWR VPWR _30594_/A sky130_fd_sc_hd__mux2_1
X_33381_ _36068_/CLK _33381_/D VGND VGND VPWR VPWR _33381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35120_ _35377_/CLK _35120_/D VGND VGND VPWR VPWR _35120_/Q sky130_fd_sc_hd__dfxtp_1
X_32332_ _32909_/CLK _32332_/D VGND VGND VPWR VPWR _32332_/Q sky130_fd_sc_hd__dfxtp_1
X_17266_ _17262_/X _17265_/X _17165_/X VGND VGND VPWR VPWR _17267_/D sky130_fd_sc_hd__o21ba_1
XFILLER_186_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16217_ _17982_/A VGND VGND VPWR VPWR _16217_/X sky130_fd_sc_hd__buf_6
X_19005_ _19001_/X _19004_/X _18726_/X VGND VGND VPWR VPWR _19037_/A sky130_fd_sc_hd__o21ba_1
XFILLER_220_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32263_ _35657_/CLK _32263_/D VGND VGND VPWR VPWR _32263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35051_ _35754_/CLK _35051_/D VGND VGND VPWR VPWR _35051_/Q sky130_fd_sc_hd__dfxtp_1
X_17197_ _17197_/A _17197_/B _17197_/C _17197_/D VGND VGND VPWR VPWR _17198_/A sky130_fd_sc_hd__or4_4
X_34002_ _34963_/CLK _34002_/D VGND VGND VPWR VPWR _34002_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31214_ _31214_/A VGND VGND VPWR VPWR _35828_/D sky130_fd_sc_hd__clkbuf_1
X_16148_ _33368_/Q _33304_/Q _33240_/Q _33176_/Q _16002_/X _16003_/X VGND VGND VPWR
+ VPWR _16148_/X sky130_fd_sc_hd__mux4_1
XFILLER_66_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32194_ _35687_/CLK _32194_/D VGND VGND VPWR VPWR _32194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31145_ _35797_/Q input60/X _31145_/S VGND VGND VPWR VPWR _31146_/A sky130_fd_sc_hd__mux2_1
X_16079_ _17935_/A VGND VGND VPWR VPWR _16079_/X sky130_fd_sc_hd__buf_6
XFILLER_233_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19907_ _20260_/A VGND VGND VPWR VPWR _19907_/X sky130_fd_sc_hd__buf_4
XFILLER_130_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35953_ _35953_/CLK _35953_/D VGND VGND VPWR VPWR _35953_/Q sky130_fd_sc_hd__dfxtp_1
X_31076_ _31145_/S VGND VGND VPWR VPWR _31095_/S sky130_fd_sc_hd__buf_8
XFILLER_229_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34904_ _34904_/CLK _34904_/D VGND VGND VPWR VPWR _34904_/Q sky130_fd_sc_hd__dfxtp_1
X_30027_ _30027_/A VGND VGND VPWR VPWR _35266_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19838_ _19651_/X _19836_/X _19837_/X _19654_/X VGND VGND VPWR VPWR _19838_/X sky130_fd_sc_hd__a22o_1
XFILLER_99_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35884_ _35949_/CLK _35884_/D VGND VGND VPWR VPWR _35884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34835_ _34963_/CLK _34835_/D VGND VGND VPWR VPWR _34835_/Q sky130_fd_sc_hd__dfxtp_1
Xinput1 DW[0] VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__buf_8
X_19769_ _35197_/Q _35133_/Q _35069_/Q _32253_/Q _19663_/X _19664_/X VGND VGND VPWR
+ VPWR _19769_/X sky130_fd_sc_hd__mux4_1
XFILLER_110_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21800_ _22506_/A VGND VGND VPWR VPWR _21800_/X sky130_fd_sc_hd__buf_6
XFILLER_65_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34766_ _34961_/CLK _34766_/D VGND VGND VPWR VPWR _34766_/Q sky130_fd_sc_hd__dfxtp_1
X_22780_ _34706_/Q _34642_/Q _34578_/Q _34514_/Q _22598_/X _22599_/X VGND VGND VPWR
+ VPWR _22780_/X sky130_fd_sc_hd__mux4_1
XFILLER_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31978_ _34790_/CLK _31978_/D VGND VGND VPWR VPWR _31978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21731_ _21453_/X _21729_/X _21730_/X _21456_/X VGND VGND VPWR VPWR _21731_/X sky130_fd_sc_hd__a22o_1
X_33717_ _35446_/CLK _33717_/D VGND VGND VPWR VPWR _33717_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30929_ _35694_/Q input17/X _30939_/S VGND VGND VPWR VPWR _30930_/A sky130_fd_sc_hd__mux2_1
X_34697_ _34698_/CLK _34697_/D VGND VGND VPWR VPWR _34697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24450_ _24450_/A VGND VGND VPWR VPWR _32753_/D sky130_fd_sc_hd__clkbuf_1
X_33648_ _34035_/CLK _33648_/D VGND VGND VPWR VPWR _33648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21662_ _22586_/A VGND VGND VPWR VPWR _21662_/X sky130_fd_sc_hd__buf_4
XFILLER_33_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23401_ _23401_/A VGND VGND VPWR VPWR _32212_/D sky130_fd_sc_hd__clkbuf_1
X_20613_ _20601_/X _20604_/X _20607_/X _20612_/X VGND VGND VPWR VPWR _20613_/X sky130_fd_sc_hd__a22o_1
XFILLER_162_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24381_ _23070_/X _32721_/Q _24381_/S VGND VGND VPWR VPWR _24382_/A sky130_fd_sc_hd__mux2_1
X_33579_ _33895_/CLK _33579_/D VGND VGND VPWR VPWR _33579_/Q sky130_fd_sc_hd__dfxtp_1
X_21593_ _22433_/A VGND VGND VPWR VPWR _21593_/X sky130_fd_sc_hd__buf_4
XFILLER_165_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26120_ _26120_/A VGND VGND VPWR VPWR _33511_/D sky130_fd_sc_hd__clkbuf_1
X_23332_ _23332_/A VGND VGND VPWR VPWR _32183_/D sky130_fd_sc_hd__clkbuf_1
X_35318_ _35446_/CLK _35318_/D VGND VGND VPWR VPWR _35318_/Q sky130_fd_sc_hd__dfxtp_1
X_20544_ _34964_/Q _34900_/Q _34836_/Q _34772_/Q _18383_/X _18385_/X VGND VGND VPWR
+ VPWR _20544_/X sky130_fd_sc_hd__mux4_1
XFILLER_177_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26051_ _24951_/X _33479_/Q _26051_/S VGND VGND VPWR VPWR _26052_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35249_ _35634_/CLK _35249_/D VGND VGND VPWR VPWR _35249_/Q sky130_fd_sc_hd__dfxtp_1
X_23263_ _32160_/Q _23261_/X _23290_/S VGND VGND VPWR VPWR _23264_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20475_ _18281_/X _20473_/X _20474_/X _18291_/X VGND VGND VPWR VPWR _20475_/X sky130_fd_sc_hd__a22o_1
XFILLER_117_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25002_ _25002_/A VGND VGND VPWR VPWR _32983_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22214_ _35201_/Q _35137_/Q _35073_/Q _32257_/Q _21963_/X _21964_/X VGND VGND VPWR
+ VPWR _22214_/X sky130_fd_sc_hd__mux4_1
XFILLER_195_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23194_ _23039_/X _32135_/Q _23194_/S VGND VGND VPWR VPWR _23195_/A sky130_fd_sc_hd__mux2_1
X_29810_ _29810_/A VGND VGND VPWR VPWR _35163_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22145_ _22106_/X _22143_/X _22144_/X _22109_/X VGND VGND VPWR VPWR _22145_/X sky130_fd_sc_hd__a22o_1
XFILLER_10_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29741_ _35131_/Q _29444_/X _29745_/S VGND VGND VPWR VPWR _29742_/A sky130_fd_sc_hd__mux2_1
X_22076_ _22076_/A VGND VGND VPWR VPWR _36221_/D sky130_fd_sc_hd__clkbuf_1
X_26953_ _26953_/A VGND VGND VPWR VPWR _33903_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25904_ _24933_/X _33409_/Q _25916_/S VGND VGND VPWR VPWR _25905_/A sky130_fd_sc_hd__mux2_1
X_21027_ _21020_/X _21025_/X _21026_/X VGND VGND VPWR VPWR _21061_/A sky130_fd_sc_hd__o21ba_1
X_29672_ _35098_/Q _29342_/X _29682_/S VGND VGND VPWR VPWR _29673_/A sky130_fd_sc_hd__mux2_1
X_26884_ _33871_/Q _23478_/X _26888_/S VGND VGND VPWR VPWR _26885_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28623_ _28623_/A VGND VGND VPWR VPWR _34632_/D sky130_fd_sc_hd__clkbuf_1
X_25835_ _24830_/X _33376_/Q _25853_/S VGND VGND VPWR VPWR _25836_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25766_ _25766_/A VGND VGND VPWR VPWR _33343_/D sky130_fd_sc_hd__clkbuf_1
X_28554_ _27698_/X _34600_/Q _28556_/S VGND VGND VPWR VPWR _28555_/A sky130_fd_sc_hd__mux2_1
X_22978_ _22977_/X _32051_/Q _22978_/S VGND VGND VPWR VPWR _22979_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27505_ _27637_/S VGND VGND VPWR VPWR _27524_/S sky130_fd_sc_hd__clkbuf_8
X_24717_ _22968_/X _32880_/Q _24723_/S VGND VGND VPWR VPWR _24718_/A sky130_fd_sc_hd__mux2_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28485_ _28485_/A VGND VGND VPWR VPWR _34567_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21929_ _34425_/Q _36153_/Q _34297_/Q _34233_/Q _21829_/X _21830_/X VGND VGND VPWR
+ VPWR _21929_/X sky130_fd_sc_hd__mux4_1
X_25697_ _24827_/X _33311_/Q _25697_/S VGND VGND VPWR VPWR _25698_/A sky130_fd_sc_hd__mux2_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27436_ _34101_/Q _27131_/X _27452_/S VGND VGND VPWR VPWR _27437_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24648_ _24648_/A VGND VGND VPWR VPWR _32847_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27367_ _34069_/Q _27229_/X _27367_/S VGND VGND VPWR VPWR _27368_/A sky130_fd_sc_hd__mux2_1
XFILLER_212_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_196_CLK clkbuf_6_49__f_CLK/X VGND VGND VPWR VPWR _35471_/CLK sky130_fd_sc_hd__clkbuf_16
X_24579_ _24579_/A VGND VGND VPWR VPWR _32814_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_212_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17120_ _16805_/X _17118_/X _17119_/X _16810_/X VGND VGND VPWR VPWR _17120_/X sky130_fd_sc_hd__a22o_1
XFILLER_106_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26318_ _26318_/A VGND VGND VPWR VPWR _33605_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29106_ _34860_/Q _27103_/X _29120_/S VGND VGND VPWR VPWR _29107_/A sky130_fd_sc_hd__mux2_1
X_27298_ _27367_/S VGND VGND VPWR VPWR _27317_/S sky130_fd_sc_hd__buf_4
XFILLER_156_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29037_ _29037_/A VGND VGND VPWR VPWR _34827_/D sky130_fd_sc_hd__clkbuf_1
X_17051_ _17051_/A VGND VGND VPWR VPWR _31985_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26249_ _26249_/A VGND VGND VPWR VPWR _33572_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16002_ _17799_/A VGND VGND VPWR VPWR _16002_/X sky130_fd_sc_hd__buf_6
XFILLER_109_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29939_ _29939_/A VGND VGND VPWR VPWR _35224_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17953_ _32139_/Q _32331_/Q _32395_/Q _35915_/Q _17633_/X _17774_/X VGND VGND VPWR
+ VPWR _17953_/X sky130_fd_sc_hd__mux4_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16904_ _33069_/Q _32045_/Q _35821_/Q _35757_/Q _16725_/X _16726_/X VGND VGND VPWR
+ VPWR _16904_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_120_CLK clkbuf_6_20__f_CLK/X VGND VGND VPWR VPWR _35544_/CLK sky130_fd_sc_hd__clkbuf_16
X_32950_ _34485_/CLK _32950_/D VGND VGND VPWR VPWR _32950_/Q sky130_fd_sc_hd__dfxtp_1
X_17884_ _17765_/X _17882_/X _17883_/X _17771_/X VGND VGND VPWR VPWR _17884_/X sky130_fd_sc_hd__a22o_1
XFILLER_65_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19623_ _33081_/Q _32057_/Q _35833_/Q _35769_/Q _19378_/X _19379_/X VGND VGND VPWR
+ VPWR _19623_/X sky130_fd_sc_hd__mux4_1
X_31901_ _31901_/A VGND VGND VPWR VPWR _36154_/D sky130_fd_sc_hd__clkbuf_1
X_16835_ _16650_/X _16833_/X _16834_/X _16653_/X VGND VGND VPWR VPWR _16835_/X sky130_fd_sc_hd__a22o_1
X_32881_ _35953_/CLK _32881_/D VGND VGND VPWR VPWR _32881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34620_ _35197_/CLK _34620_/D VGND VGND VPWR VPWR _34620_/Q sky130_fd_sc_hd__dfxtp_1
X_31832_ _31832_/A VGND VGND VPWR VPWR _36121_/D sky130_fd_sc_hd__clkbuf_1
X_19554_ _20260_/A VGND VGND VPWR VPWR _19554_/X sky130_fd_sc_hd__buf_6
XFILLER_0_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16766_ _34921_/Q _34857_/Q _34793_/Q _34729_/Q _16454_/X _16455_/X VGND VGND VPWR
+ VPWR _16766_/X sky130_fd_sc_hd__mux4_1
XFILLER_4_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18505_ _34905_/Q _34841_/Q _34777_/Q _34713_/Q _18396_/X _18398_/X VGND VGND VPWR
+ VPWR _18505_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34551_ _36024_/CLK _34551_/D VGND VGND VPWR VPWR _34551_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31763_ _36089_/Q input29/X _31771_/S VGND VGND VPWR VPWR _31764_/A sky130_fd_sc_hd__mux2_1
X_19485_ _19298_/X _19483_/X _19484_/X _19301_/X VGND VGND VPWR VPWR _19485_/X sky130_fd_sc_hd__a22o_1
X_16697_ _16697_/A _16697_/B _16697_/C _16697_/D VGND VGND VPWR VPWR _16698_/A sky130_fd_sc_hd__or4_2
XFILLER_94_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33502_ _36191_/CLK _33502_/D VGND VGND VPWR VPWR _33502_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18436_ _18391_/X _18434_/X _18435_/X _18401_/X VGND VGND VPWR VPWR _18436_/X sky130_fd_sc_hd__a22o_1
X_30714_ _35592_/Q _29484_/X _30732_/S VGND VGND VPWR VPWR _30715_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34482_ _34611_/CLK _34482_/D VGND VGND VPWR VPWR _34482_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31694_ _36056_/Q input23/X _31708_/S VGND VGND VPWR VPWR _31695_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36221_ _36223_/CLK _36221_/D VGND VGND VPWR VPWR _36221_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33433_ _34009_/CLK _33433_/D VGND VGND VPWR VPWR _33433_/Q sky130_fd_sc_hd__dfxtp_1
X_18367_ _20235_/A VGND VGND VPWR VPWR _18367_/X sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_187_CLK clkbuf_leaf_65_CLK/A VGND VGND VPWR VPWR _36047_/CLK sky130_fd_sc_hd__clkbuf_16
X_30645_ _30645_/A VGND VGND VPWR VPWR _35559_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17318_ _17800_/A VGND VGND VPWR VPWR _17318_/X sky130_fd_sc_hd__buf_4
X_36152_ _36152_/CLK _36152_/D VGND VGND VPWR VPWR _36152_/Q sky130_fd_sc_hd__dfxtp_1
X_33364_ _36180_/CLK _33364_/D VGND VGND VPWR VPWR _33364_/Q sky130_fd_sc_hd__dfxtp_1
X_30576_ _35527_/Q _29481_/X _30576_/S VGND VGND VPWR VPWR _30577_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18298_ input79/X input80/X VGND VGND VPWR VPWR _18299_/A sky130_fd_sc_hd__and2_1
X_35103_ _35610_/CLK _35103_/D VGND VGND VPWR VPWR _35103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32315_ _35962_/CLK _32315_/D VGND VGND VPWR VPWR _32315_/Q sky130_fd_sc_hd__dfxtp_1
X_36083_ _36085_/CLK _36083_/D VGND VGND VPWR VPWR _36083_/Q sky130_fd_sc_hd__dfxtp_1
X_17249_ _17067_/X _17247_/X _17248_/X _17071_/X VGND VGND VPWR VPWR _17249_/X sky130_fd_sc_hd__a22o_1
X_33295_ _33425_/CLK _33295_/D VGND VGND VPWR VPWR _33295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35034_ _35162_/CLK _35034_/D VGND VGND VPWR VPWR _35034_/Q sky130_fd_sc_hd__dfxtp_1
X_20260_ _20260_/A VGND VGND VPWR VPWR _20260_/X sky130_fd_sc_hd__buf_4
X_32246_ _36149_/CLK _32246_/D VGND VGND VPWR VPWR _32246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32177_ _35735_/CLK _32177_/D VGND VGND VPWR VPWR _32177_/Q sky130_fd_sc_hd__dfxtp_1
X_20191_ _20004_/X _20189_/X _20190_/X _20007_/X VGND VGND VPWR VPWR _20191_/X sky130_fd_sc_hd__a22o_1
XFILLER_88_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31128_ _31128_/A VGND VGND VPWR VPWR _35788_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_111_CLK clkbuf_6_22__f_CLK/X VGND VGND VPWR VPWR _35674_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23950_ _23977_/S VGND VGND VPWR VPWR _23969_/S sky130_fd_sc_hd__buf_4
X_35936_ _35938_/CLK _35936_/D VGND VGND VPWR VPWR _35936_/Q sky130_fd_sc_hd__dfxtp_1
X_31059_ _31059_/A VGND VGND VPWR VPWR _35755_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_229_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22901_ _22900_/X _32026_/Q _22916_/S VGND VGND VPWR VPWR _22902_/A sky130_fd_sc_hd__mux2_1
XTAP_3908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35867_ _35995_/CLK _35867_/D VGND VGND VPWR VPWR _35867_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23881_ _22940_/X _32487_/Q _23885_/S VGND VGND VPWR VPWR _23882_/A sky130_fd_sc_hd__mux2_1
XFILLER_245_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25620_ _25620_/A VGND VGND VPWR VPWR _33274_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34818_ _36163_/CLK _34818_/D VGND VGND VPWR VPWR _34818_/Q sky130_fd_sc_hd__dfxtp_1
X_22832_ _22828_/X _22831_/X _22446_/A _22447_/A VGND VGND VPWR VPWR _22847_/B sky130_fd_sc_hd__o211a_1
XFILLER_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35798_ _36118_/CLK _35798_/D VGND VGND VPWR VPWR _35798_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_6_41__f_CLK clkbuf_5_20_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_41__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_225_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25551_ _25551_/A VGND VGND VPWR VPWR _33241_/D sky130_fd_sc_hd__clkbuf_1
X_22763_ _33938_/Q _33874_/Q _33810_/Q _36114_/Q _20662_/X _20664_/X VGND VGND VPWR
+ VPWR _22763_/X sky130_fd_sc_hd__mux4_1
X_34749_ _34877_/CLK _34749_/D VGND VGND VPWR VPWR _34749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24502_ _23049_/X _32778_/Q _24516_/S VGND VGND VPWR VPWR _24503_/A sky130_fd_sc_hd__mux2_1
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_240_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21714_ _21710_/X _21713_/X _21398_/X VGND VGND VPWR VPWR _21722_/C sky130_fd_sc_hd__o21ba_1
X_28270_ _27677_/X _34465_/Q _28286_/S VGND VGND VPWR VPWR _28271_/A sky130_fd_sc_hd__mux2_1
X_25482_ _24908_/X _33209_/Q _25490_/S VGND VGND VPWR VPWR _25483_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22694_ _34959_/Q _34895_/Q _34831_/Q _34767_/Q _22466_/X _22467_/X VGND VGND VPWR
+ VPWR _22694_/X sky130_fd_sc_hd__mux4_1
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27221_ _34002_/Q _27220_/X _27230_/S VGND VGND VPWR VPWR _27222_/A sky130_fd_sc_hd__mux2_1
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24433_ _24433_/A VGND VGND VPWR VPWR _32745_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_178_CLK clkbuf_6_27__f_CLK/X VGND VGND VPWR VPWR _35666_/CLK sky130_fd_sc_hd__clkbuf_16
X_21645_ _21400_/X _21643_/X _21644_/X _21403_/X VGND VGND VPWR VPWR _21645_/X sky130_fd_sc_hd__a22o_1
XFILLER_234_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27152_ input32/X VGND VGND VPWR VPWR _27152_/X sky130_fd_sc_hd__clkbuf_4
X_24364_ _24364_/A VGND VGND VPWR VPWR _32712_/D sky130_fd_sc_hd__clkbuf_1
X_21576_ _34415_/Q _36143_/Q _34287_/Q _34223_/Q _21476_/X _21477_/X VGND VGND VPWR
+ VPWR _21576_/X sky130_fd_sc_hd__mux4_1
XFILLER_205_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26103_ _26103_/A VGND VGND VPWR VPWR _33503_/D sky130_fd_sc_hd__clkbuf_1
X_23315_ _23315_/A VGND VGND VPWR VPWR _32175_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20527_ _33172_/Q _36052_/Q _33044_/Q _32980_/Q _18332_/X _19461_/A VGND VGND VPWR
+ VPWR _20527_/X sky130_fd_sc_hd__mux4_1
X_27083_ _27083_/A VGND VGND VPWR VPWR _33957_/D sky130_fd_sc_hd__clkbuf_1
X_24295_ _22943_/X _32680_/Q _24297_/S VGND VGND VPWR VPWR _24296_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26034_ _26034_/A VGND VGND VPWR VPWR _33470_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23246_ input56/X VGND VGND VPWR VPWR _23246_/X sky130_fd_sc_hd__buf_4
XFILLER_4_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20458_ _20458_/A VGND VGND VPWR VPWR _32465_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_88_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23177_ _23177_/A VGND VGND VPWR VPWR _32126_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_350_CLK clkbuf_6_47__f_CLK/X VGND VGND VPWR VPWR _35453_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_6501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20389_ _20385_/X _20388_/X _20157_/X VGND VGND VPWR VPWR _20397_/C sky130_fd_sc_hd__o21ba_1
XFILLER_122_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22128_ _22124_/X _22127_/X _22085_/X VGND VGND VPWR VPWR _22150_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput190 _36224_/Q VGND VGND VPWR VPWR D2[42] sky130_fd_sc_hd__buf_2
XTAP_5800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27985_ _34330_/Q _27047_/X _27995_/S VGND VGND VPWR VPWR _27986_/A sky130_fd_sc_hd__mux2_1
XTAP_6556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29724_ _35123_/Q _29419_/X _29724_/S VGND VGND VPWR VPWR _29725_/A sky130_fd_sc_hd__mux2_1
XFILLER_212_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_102_CLK clkbuf_leaf_99_CLK/A VGND VGND VPWR VPWR _34009_/CLK sky130_fd_sc_hd__clkbuf_16
X_22059_ _22020_/X _22057_/X _22058_/X _22024_/X VGND VGND VPWR VPWR _22059_/X sky130_fd_sc_hd__a22o_1
X_26936_ _26936_/A VGND VGND VPWR VPWR _33895_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29655_ _29655_/A VGND VGND VPWR VPWR _35090_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26867_ _33863_/Q _23450_/X _26867_/S VGND VGND VPWR VPWR _26868_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28606_ _28606_/A VGND VGND VPWR VPWR _34624_/D sky130_fd_sc_hd__clkbuf_1
X_16620_ _34661_/Q _34597_/Q _34533_/Q _34469_/Q _16586_/X _16587_/X VGND VGND VPWR
+ VPWR _16620_/X sky130_fd_sc_hd__mux4_1
X_25818_ _24806_/X _33368_/Q _25832_/S VGND VGND VPWR VPWR _25819_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26798_ _33830_/Q _23280_/X _26804_/S VGND VGND VPWR VPWR _26799_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29586_ _29586_/A VGND VGND VPWR VPWR _35057_/D sky130_fd_sc_hd__clkbuf_1
X_16551_ _33059_/Q _32035_/Q _35811_/Q _35747_/Q _16372_/X _16373_/X VGND VGND VPWR
+ VPWR _16551_/X sky130_fd_sc_hd__mux4_1
X_25749_ _25749_/A VGND VGND VPWR VPWR _33335_/D sky130_fd_sc_hd__clkbuf_1
X_28537_ _28648_/S VGND VGND VPWR VPWR _28556_/S sky130_fd_sc_hd__buf_6
XFILLER_204_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19270_ _33071_/Q _32047_/Q _35823_/Q _35759_/Q _19025_/X _19026_/X VGND VGND VPWR
+ VPWR _19270_/X sky130_fd_sc_hd__mux4_1
X_16482_ _16297_/X _16480_/X _16481_/X _16300_/X VGND VGND VPWR VPWR _16482_/X sky130_fd_sc_hd__a22o_1
X_28468_ _27770_/X _34559_/Q _28484_/S VGND VGND VPWR VPWR _28469_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18221_ _16018_/X _18219_/X _18220_/X _16027_/X VGND VGND VPWR VPWR _18221_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_169_CLK clkbuf_6_30__f_CLK/X VGND VGND VPWR VPWR _34708_/CLK sky130_fd_sc_hd__clkbuf_16
X_27419_ _34093_/Q _27106_/X _27431_/S VGND VGND VPWR VPWR _27420_/A sky130_fd_sc_hd__mux2_1
X_28399_ _28399_/A VGND VGND VPWR VPWR _34526_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30430_ _30430_/A VGND VGND VPWR VPWR _35457_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18152_ _17859_/X _18150_/X _18151_/X _17862_/X VGND VGND VPWR VPWR _18152_/X sky130_fd_sc_hd__a22o_1
XFILLER_184_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17103_ _17059_/X _17101_/X _17102_/X _17065_/X VGND VGND VPWR VPWR _17103_/X sky130_fd_sc_hd__a22o_1
X_18083_ _35727_/Q _32238_/Q _35599_/Q _35535_/Q _15993_/X _15995_/X VGND VGND VPWR
+ VPWR _18083_/X sky130_fd_sc_hd__mux4_1
XFILLER_141_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30361_ _30361_/A VGND VGND VPWR VPWR _35424_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17034_ _16714_/X _17032_/X _17033_/X _16718_/X VGND VGND VPWR VPWR _17034_/X sky130_fd_sc_hd__a22o_1
X_32100_ _32356_/CLK _32100_/D VGND VGND VPWR VPWR _32100_/Q sky130_fd_sc_hd__dfxtp_1
X_33080_ _35768_/CLK _33080_/D VGND VGND VPWR VPWR _33080_/Q sky130_fd_sc_hd__dfxtp_1
X_30292_ _35392_/Q _29460_/X _30306_/S VGND VGND VPWR VPWR _30293_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32031_ _35677_/CLK _32031_/D VGND VGND VPWR VPWR _32031_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_341_CLK clkbuf_6_45__f_CLK/X VGND VGND VPWR VPWR _32894_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_124_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_891 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18985_ _18945_/X _18983_/X _18984_/X _18948_/X VGND VGND VPWR VPWR _18985_/X sky130_fd_sc_hd__a22o_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17936_ _17936_/A VGND VGND VPWR VPWR _17936_/X sky130_fd_sc_hd__buf_4
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33982_ _34174_/CLK _33982_/D VGND VGND VPWR VPWR _33982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35721_ _35721_/CLK _35721_/D VGND VGND VPWR VPWR _35721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32933_ _36005_/CLK _32933_/D VGND VGND VPWR VPWR _32933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17867_ _17867_/A VGND VGND VPWR VPWR _17867_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_94_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19606_ _33401_/Q _33337_/Q _33273_/Q _33209_/Q _19427_/X _19428_/X VGND VGND VPWR
+ VPWR _19606_/X sky130_fd_sc_hd__mux4_1
XFILLER_187_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35652_ _35716_/CLK _35652_/D VGND VGND VPWR VPWR _35652_/Q sky130_fd_sc_hd__dfxtp_1
X_16818_ _16493_/X _16816_/X _16817_/X _16498_/X VGND VGND VPWR VPWR _16818_/X sky130_fd_sc_hd__a22o_1
X_32864_ _35871_/CLK _32864_/D VGND VGND VPWR VPWR _32864_/Q sky130_fd_sc_hd__dfxtp_1
X_17798_ _33671_/Q _33607_/Q _33543_/Q _33479_/Q _17553_/X _17554_/X VGND VGND VPWR
+ VPWR _17798_/X sky130_fd_sc_hd__mux4_1
XFILLER_19_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34603_ _35754_/CLK _34603_/D VGND VGND VPWR VPWR _34603_/Q sky130_fd_sc_hd__dfxtp_1
X_31815_ _36114_/Q input57/X _31821_/S VGND VGND VPWR VPWR _31816_/A sky130_fd_sc_hd__mux2_1
X_19537_ _33655_/Q _33591_/Q _33527_/Q _33463_/Q _19500_/X _19501_/X VGND VGND VPWR
+ VPWR _19537_/X sky130_fd_sc_hd__mux4_1
X_35583_ _35713_/CLK _35583_/D VGND VGND VPWR VPWR _35583_/Q sky130_fd_sc_hd__dfxtp_1
X_16749_ _33129_/Q _36009_/Q _33001_/Q _32937_/Q _16709_/X _16710_/X VGND VGND VPWR
+ VPWR _16749_/X sky130_fd_sc_hd__mux4_1
X_32795_ _35669_/CLK _32795_/D VGND VGND VPWR VPWR _32795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_1052 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34534_ _36137_/CLK _34534_/D VGND VGND VPWR VPWR _34534_/Q sky130_fd_sc_hd__dfxtp_1
X_31746_ _36081_/Q input20/X _31750_/S VGND VGND VPWR VPWR _31747_/A sky130_fd_sc_hd__mux2_1
X_19468_ _19468_/A VGND VGND VPWR VPWR _32436_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_35_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_1085 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18419_ _18318_/X _18417_/X _18418_/X _18327_/X VGND VGND VPWR VPWR _18419_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34465_ _35297_/CLK _34465_/D VGND VGND VPWR VPWR _34465_/Q sky130_fd_sc_hd__dfxtp_1
X_31677_ _31677_/A VGND VGND VPWR VPWR _36048_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19399_ _19153_/X _19397_/X _19398_/X _19156_/X VGND VGND VPWR VPWR _19399_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36204_ _36207_/CLK _36204_/D VGND VGND VPWR VPWR _36204_/Q sky130_fd_sc_hd__dfxtp_1
X_33416_ _33673_/CLK _33416_/D VGND VGND VPWR VPWR _33416_/Q sky130_fd_sc_hd__dfxtp_1
X_21430_ _35691_/Q _32199_/Q _35563_/Q _35499_/Q _21211_/X _21212_/X VGND VGND VPWR
+ VPWR _21430_/X sky130_fd_sc_hd__mux4_1
X_30628_ _30628_/A VGND VGND VPWR VPWR _35551_/D sky130_fd_sc_hd__clkbuf_1
X_34396_ _36235_/CLK _34396_/D VGND VGND VPWR VPWR _34396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36135_ _36135_/CLK _36135_/D VGND VGND VPWR VPWR _36135_/Q sky130_fd_sc_hd__dfxtp_1
X_33347_ _33924_/CLK _33347_/D VGND VGND VPWR VPWR _33347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21361_ _21357_/X _21360_/X _21045_/X VGND VGND VPWR VPWR _21369_/C sky130_fd_sc_hd__o21ba_1
X_30559_ _30559_/A VGND VGND VPWR VPWR _35518_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23100_ _22900_/X _32090_/Q _23110_/S VGND VGND VPWR VPWR _23101_/A sky130_fd_sc_hd__mux2_1
X_20312_ _33421_/Q _33357_/Q _33293_/Q _33229_/Q _20133_/X _20134_/X VGND VGND VPWR
+ VPWR _20312_/X sky130_fd_sc_hd__mux4_1
Xinput70 R1[5] VGND VGND VPWR VPWR input70/X sky130_fd_sc_hd__clkbuf_4
X_24080_ _23033_/X _32581_/Q _24084_/S VGND VGND VPWR VPWR _24081_/A sky130_fd_sc_hd__mux2_1
X_36066_ _36066_/CLK _36066_/D VGND VGND VPWR VPWR _36066_/Q sky130_fd_sc_hd__dfxtp_1
Xinput81 R3[4] VGND VGND VPWR VPWR input81/X sky130_fd_sc_hd__buf_2
XFILLER_174_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33278_ _35711_/CLK _33278_/D VGND VGND VPWR VPWR _33278_/Q sky130_fd_sc_hd__dfxtp_1
X_21292_ _21047_/X _21290_/X _21291_/X _21050_/X VGND VGND VPWR VPWR _21292_/X sky130_fd_sc_hd__a22o_1
X_35017_ _35658_/CLK _35017_/D VGND VGND VPWR VPWR _35017_/Q sky130_fd_sc_hd__dfxtp_1
X_23031_ _23030_/X _32068_/Q _23040_/S VGND VGND VPWR VPWR _23032_/A sky130_fd_sc_hd__mux2_1
X_20243_ _33675_/Q _33611_/Q _33547_/Q _33483_/Q _20206_/X _20207_/X VGND VGND VPWR
+ VPWR _20243_/X sky130_fd_sc_hd__mux4_1
X_32229_ _35463_/CLK _32229_/D VGND VGND VPWR VPWR _32229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_332_CLK clkbuf_6_38__f_CLK/X VGND VGND VPWR VPWR _34485_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_190_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20174_ _20174_/A VGND VGND VPWR VPWR _32456_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_104_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24982_ input55/X VGND VGND VPWR VPWR _24982_/X sky130_fd_sc_hd__buf_4
X_27770_ input36/X VGND VGND VPWR VPWR _27770_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_130_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26721_ _26721_/A VGND VGND VPWR VPWR _33793_/D sky130_fd_sc_hd__clkbuf_1
X_23933_ _23933_/A VGND VGND VPWR VPWR _32511_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_245_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35919_ _35983_/CLK _35919_/D VGND VGND VPWR VPWR _35919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26652_ _26652_/A VGND VGND VPWR VPWR _33760_/D sky130_fd_sc_hd__clkbuf_1
X_29440_ _29440_/A VGND VGND VPWR VPWR _35001_/D sky130_fd_sc_hd__clkbuf_1
X_23864_ _22915_/X _32479_/Q _23864_/S VGND VGND VPWR VPWR _23865_/A sky130_fd_sc_hd__mux2_1
XTAP_3749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25603_ _25603_/A VGND VGND VPWR VPWR _33266_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22815_ _20660_/X _22813_/X _22814_/X _20672_/X VGND VGND VPWR VPWR _22815_/X sky130_fd_sc_hd__a22o_1
X_26583_ _24936_/X _33730_/Q _26593_/S VGND VGND VPWR VPWR _26584_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_399_CLK clkbuf_6_35__f_CLK/X VGND VGND VPWR VPWR _35765_/CLK sky130_fd_sc_hd__clkbuf_16
X_29371_ _34979_/Q _29370_/X _29389_/S VGND VGND VPWR VPWR _29372_/A sky130_fd_sc_hd__mux2_1
X_23795_ _23015_/X _32383_/Q _23811_/S VGND VGND VPWR VPWR _23796_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25534_ _24985_/X _33234_/Q _25540_/S VGND VGND VPWR VPWR _25535_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28322_ _27754_/X _34490_/Q _28328_/S VGND VGND VPWR VPWR _28323_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22746_ _35473_/Q _35409_/Q _35345_/Q _35281_/Q _22560_/X _22561_/X VGND VGND VPWR
+ VPWR _22746_/X sky130_fd_sc_hd__mux4_1
XFILLER_164_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28253_ _27652_/X _34457_/Q _28265_/S VGND VGND VPWR VPWR _28254_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25465_ _24883_/X _33201_/Q _25469_/S VGND VGND VPWR VPWR _25466_/A sky130_fd_sc_hd__mux2_1
X_22677_ _33167_/Q _36047_/Q _33039_/Q _32975_/Q _22368_/X _22369_/X VGND VGND VPWR
+ VPWR _22677_/X sky130_fd_sc_hd__mux4_1
XFILLER_201_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27204_ _27204_/A VGND VGND VPWR VPWR _33996_/D sky130_fd_sc_hd__clkbuf_1
X_24416_ _22922_/X _32737_/Q _24432_/S VGND VGND VPWR VPWR _24417_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_1314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21628_ _21622_/X _21627_/X _21379_/X VGND VGND VPWR VPWR _21650_/A sky130_fd_sc_hd__o21ba_1
X_28184_ _28184_/A VGND VGND VPWR VPWR _34424_/D sky130_fd_sc_hd__clkbuf_1
X_25396_ _25396_/A VGND VGND VPWR VPWR _33169_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27135_ _33974_/Q _27134_/X _27156_/S VGND VGND VPWR VPWR _27136_/A sky130_fd_sc_hd__mux2_1
X_24347_ _24347_/A VGND VGND VPWR VPWR _32704_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21559_ _21306_/X _21557_/X _21558_/X _21312_/X VGND VGND VPWR VPWR _21559_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27066_ _27230_/S VGND VGND VPWR VPWR _27094_/S sky130_fd_sc_hd__buf_6
XFILLER_4_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24278_ _24389_/S VGND VGND VPWR VPWR _24297_/S sky130_fd_sc_hd__buf_4
XFILLER_181_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26017_ _26017_/A VGND VGND VPWR VPWR _33462_/D sky130_fd_sc_hd__clkbuf_1
XTAP_7010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23229_ _23229_/A VGND VGND VPWR VPWR _30472_/A sky130_fd_sc_hd__buf_4
XTAP_7021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_323_CLK clkbuf_6_39__f_CLK/X VGND VGND VPWR VPWR _32905_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_7032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18770_ _32609_/Q _32545_/Q _32481_/Q _35937_/Q _18517_/X _18654_/X VGND VGND VPWR
+ VPWR _18770_/X sky130_fd_sc_hd__mux4_1
XFILLER_67_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15982_ input65/X VGND VGND VPWR VPWR _16061_/A sky130_fd_sc_hd__buf_8
X_27968_ _27968_/A VGND VGND VPWR VPWR _34322_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17721_ _34948_/Q _34884_/Q _34820_/Q _34756_/Q _17513_/X _17514_/X VGND VGND VPWR
+ VPWR _17721_/X sky130_fd_sc_hd__mux4_1
XTAP_5663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29707_ _29707_/A VGND VGND VPWR VPWR _35114_/D sky130_fd_sc_hd__clkbuf_1
X_26919_ _26919_/A VGND VGND VPWR VPWR _33887_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27899_ _27899_/A VGND VGND VPWR VPWR _34289_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17652_ _17511_/X _17650_/X _17651_/X _17516_/X VGND VGND VPWR VPWR _17652_/X sky130_fd_sc_hd__a22o_1
X_29638_ _35082_/Q _29491_/X _29652_/S VGND VGND VPWR VPWR _29639_/A sky130_fd_sc_hd__mux2_1
XTAP_4973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16603_ _16599_/X _16602_/X _16426_/X VGND VGND VPWR VPWR _16627_/A sky130_fd_sc_hd__o21ba_1
XFILLER_95_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17583_ _17936_/A VGND VGND VPWR VPWR _17583_/X sky130_fd_sc_hd__buf_4
XFILLER_28_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29569_ _29569_/A VGND VGND VPWR VPWR _35049_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19322_ _19146_/X _19320_/X _19321_/X _19151_/X VGND VGND VPWR VPWR _19322_/X sky130_fd_sc_hd__a22o_1
X_31600_ _31600_/A VGND VGND VPWR VPWR _36011_/D sky130_fd_sc_hd__clkbuf_1
X_16534_ _33379_/Q _33315_/Q _33251_/Q _33187_/Q _16421_/X _16422_/X VGND VGND VPWR
+ VPWR _16534_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32580_ _35973_/CLK _32580_/D VGND VGND VPWR VPWR _32580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_1206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31531_ _27807_/X _35979_/Q _31543_/S VGND VGND VPWR VPWR _31532_/A sky130_fd_sc_hd__mux2_1
X_19253_ _33391_/Q _33327_/Q _33263_/Q _33199_/Q _19074_/X _19075_/X VGND VGND VPWR
+ VPWR _19253_/X sky130_fd_sc_hd__mux4_1
XFILLER_31_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16465_ _16140_/X _16463_/X _16464_/X _16145_/X VGND VGND VPWR VPWR _16465_/X sky130_fd_sc_hd__a22o_1
XFILLER_188_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18204_ _35667_/Q _35027_/Q _34387_/Q _33747_/Q _16112_/X _16113_/X VGND VGND VPWR
+ VPWR _18204_/X sky130_fd_sc_hd__mux4_1
XPHY_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34250_ _34956_/CLK _34250_/D VGND VGND VPWR VPWR _34250_/Q sky130_fd_sc_hd__dfxtp_1
X_16396_ _33119_/Q _35999_/Q _32991_/Q _32927_/Q _16356_/X _16357_/X VGND VGND VPWR
+ VPWR _16396_/X sky130_fd_sc_hd__mux4_1
X_19184_ _33645_/Q _33581_/Q _33517_/Q _33453_/Q _19147_/X _19148_/X VGND VGND VPWR
+ VPWR _19184_/X sky130_fd_sc_hd__mux4_1
X_31462_ _27704_/X _35946_/Q _31480_/S VGND VGND VPWR VPWR _31463_/A sky130_fd_sc_hd__mux2_1
XPHY_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33201_ _33904_/CLK _33201_/D VGND VGND VPWR VPWR _33201_/Q sky130_fd_sc_hd__dfxtp_1
X_18135_ _18131_/X _18134_/X _17838_/X VGND VGND VPWR VPWR _18157_/A sky130_fd_sc_hd__o21ba_2
X_30413_ _30413_/A VGND VGND VPWR VPWR _35449_/D sky130_fd_sc_hd__clkbuf_1
X_34181_ _34183_/CLK _34181_/D VGND VGND VPWR VPWR _34181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31393_ _31393_/A VGND VGND VPWR VPWR _35913_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_1034 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33132_ _36013_/CLK _33132_/D VGND VGND VPWR VPWR _33132_/Q sky130_fd_sc_hd__dfxtp_1
X_30344_ _30344_/A VGND VGND VPWR VPWR _35416_/D sky130_fd_sc_hd__clkbuf_1
X_18066_ _18062_/X _18065_/X _17871_/X VGND VGND VPWR VPWR _18067_/D sky130_fd_sc_hd__o21ba_1
XFILLER_67_1310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17017_ _17013_/X _17016_/X _16812_/X VGND VGND VPWR VPWR _17018_/D sky130_fd_sc_hd__o21ba_1
Xclkbuf_6_5__f_CLK clkbuf_5_2_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_5__f_CLK/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_314_CLK clkbuf_6_48__f_CLK/X VGND VGND VPWR VPWR _35978_/CLK sky130_fd_sc_hd__clkbuf_16
X_30275_ _35384_/Q _29435_/X _30285_/S VGND VGND VPWR VPWR _30276_/A sky130_fd_sc_hd__mux2_1
X_33063_ _35755_/CLK _33063_/D VGND VGND VPWR VPWR _33063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32014_ _36202_/CLK _32014_/D VGND VGND VPWR VPWR _32014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18968_ _34151_/Q _34087_/Q _34023_/Q _33959_/Q _18687_/X _18688_/X VGND VGND VPWR
+ VPWR _18968_/X sky130_fd_sc_hd__mux4_2
XFILLER_26_1062 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17919_ _33162_/Q _36042_/Q _33034_/Q _32970_/Q _17768_/X _17769_/X VGND VGND VPWR
+ VPWR _17919_/X sky130_fd_sc_hd__mux4_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33965_ _35693_/CLK _33965_/D VGND VGND VPWR VPWR _33965_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18899_ _18793_/X _18897_/X _18898_/X _18798_/X VGND VGND VPWR VPWR _18899_/X sky130_fd_sc_hd__a22o_1
X_35704_ _35704_/CLK _35704_/D VGND VGND VPWR VPWR _35704_/Q sky130_fd_sc_hd__dfxtp_1
X_20930_ _35677_/Q _32183_/Q _35549_/Q _35485_/Q _20858_/X _20859_/X VGND VGND VPWR
+ VPWR _20930_/X sky130_fd_sc_hd__mux4_1
X_32916_ _35922_/CLK _32916_/D VGND VGND VPWR VPWR _32916_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_230_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33896_ _33897_/CLK _33896_/D VGND VGND VPWR VPWR _33896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35635_ _35635_/CLK _35635_/D VGND VGND VPWR VPWR _35635_/Q sky130_fd_sc_hd__dfxtp_1
X_20861_ _35611_/Q _34971_/Q _34331_/Q _33691_/Q _20653_/X _20655_/X VGND VGND VPWR
+ VPWR _20861_/X sky130_fd_sc_hd__mux4_1
XFILLER_148_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32847_ _32879_/CLK _32847_/D VGND VGND VPWR VPWR _32847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22600_ _34700_/Q _34636_/Q _34572_/Q _34508_/Q _22598_/X _22599_/X VGND VGND VPWR
+ VPWR _22600_/X sky130_fd_sc_hd__mux4_1
XFILLER_207_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23580_ _23580_/A VGND VGND VPWR VPWR _32282_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35566_ _35566_/CLK _35566_/D VGND VGND VPWR VPWR _35566_/Q sky130_fd_sc_hd__dfxtp_1
X_20792_ _35673_/Q _32179_/Q _35545_/Q _35481_/Q _20649_/X _20650_/X VGND VGND VPWR
+ VPWR _20792_/X sky130_fd_sc_hd__mux4_1
X_32778_ _32907_/CLK _32778_/D VGND VGND VPWR VPWR _32778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34517_ _36117_/CLK _34517_/D VGND VGND VPWR VPWR _34517_/Q sky130_fd_sc_hd__dfxtp_1
X_22531_ _22527_/X _22530_/X _22457_/X VGND VGND VPWR VPWR _22541_/C sky130_fd_sc_hd__o21ba_1
X_31729_ _36073_/Q input11/X _31729_/S VGND VGND VPWR VPWR _31730_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35497_ _35685_/CLK _35497_/D VGND VGND VPWR VPWR _35497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25250_ _25250_/A VGND VGND VPWR VPWR _33100_/D sky130_fd_sc_hd__clkbuf_1
X_34448_ _36176_/CLK _34448_/D VGND VGND VPWR VPWR _34448_/Q sky130_fd_sc_hd__dfxtp_1
X_22462_ _22462_/A VGND VGND VPWR VPWR _22462_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_167_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_950 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24201_ _32637_/Q _23417_/X _24201_/S VGND VGND VPWR VPWR _24202_/A sky130_fd_sc_hd__mux2_1
XFILLER_202_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21413_ _21404_/X _21411_/X _21412_/X VGND VGND VPWR VPWR _21414_/D sky130_fd_sc_hd__o21ba_1
X_25181_ _25181_/A VGND VGND VPWR VPWR _33067_/D sky130_fd_sc_hd__clkbuf_1
X_22393_ _34950_/Q _34886_/Q _34822_/Q _34758_/Q _22113_/X _22114_/X VGND VGND VPWR
+ VPWR _22393_/X sky130_fd_sc_hd__mux4_1
X_34379_ _35661_/CLK _34379_/D VGND VGND VPWR VPWR _34379_/Q sky130_fd_sc_hd__dfxtp_1
X_36118_ _36118_/CLK _36118_/D VGND VGND VPWR VPWR _36118_/Q sky130_fd_sc_hd__dfxtp_1
X_24132_ _32604_/Q _23249_/X _24138_/S VGND VGND VPWR VPWR _24133_/A sky130_fd_sc_hd__mux2_1
XFILLER_136_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21344_ _33385_/Q _33321_/Q _33257_/Q _33193_/Q _21021_/X _21022_/X VGND VGND VPWR
+ VPWR _21344_/X sky130_fd_sc_hd__mux4_1
XFILLER_108_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28940_ _28940_/A VGND VGND VPWR VPWR _34781_/D sky130_fd_sc_hd__clkbuf_1
X_36049_ _36049_/CLK _36049_/D VGND VGND VPWR VPWR _36049_/Q sky130_fd_sc_hd__dfxtp_1
X_24063_ _23008_/X _32573_/Q _24063_/S VGND VGND VPWR VPWR _24064_/A sky130_fd_sc_hd__mux2_1
XFILLER_235_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_305_CLK clkbuf_6_51__f_CLK/X VGND VGND VPWR VPWR _35847_/CLK sky130_fd_sc_hd__clkbuf_16
X_21275_ _21269_/X _21274_/X _21026_/X VGND VGND VPWR VPWR _21297_/A sky130_fd_sc_hd__o21ba_1
XFILLER_46_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23014_ _23014_/A VGND VGND VPWR VPWR _32062_/D sky130_fd_sc_hd__clkbuf_1
X_20226_ _35658_/Q _35018_/Q _34378_/Q _33738_/Q _20150_/X _20151_/X VGND VGND VPWR
+ VPWR _20226_/X sky130_fd_sc_hd__mux4_1
XFILLER_172_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28871_ _34749_/Q _27155_/X _28871_/S VGND VGND VPWR VPWR _28872_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27822_ input54/X VGND VGND VPWR VPWR _27822_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_49_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20157_ _20157_/A VGND VGND VPWR VPWR _20157_/X sky130_fd_sc_hd__buf_2
XFILLER_172_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_1421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_246_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24965_ _24964_/X _32971_/Q _24983_/S VGND VGND VPWR VPWR _24966_/A sky130_fd_sc_hd__mux2_1
XTAP_4225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27753_ _27753_/A VGND VGND VPWR VPWR _34233_/D sky130_fd_sc_hd__clkbuf_1
X_20088_ _20082_/X _20087_/X _19804_/X VGND VGND VPWR VPWR _20096_/C sky130_fd_sc_hd__o21ba_1
XTAP_4236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26704_ _26704_/A VGND VGND VPWR VPWR _33785_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23916_ _23916_/A VGND VGND VPWR VPWR _32503_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24896_ input25/X VGND VGND VPWR VPWR _24896_/X sky130_fd_sc_hd__clkbuf_4
X_27684_ _27683_/X _34211_/Q _27702_/S VGND VGND VPWR VPWR _27685_/A sky130_fd_sc_hd__mux2_1
XTAP_3546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29423_ _29525_/S VGND VGND VPWR VPWR _29451_/S sky130_fd_sc_hd__buf_6
XFILLER_72_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23847_ _23847_/A VGND VGND VPWR VPWR _32470_/D sky130_fd_sc_hd__clkbuf_1
X_26635_ _26635_/A VGND VGND VPWR VPWR _33752_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29354_ input63/X VGND VGND VPWR VPWR _29354_/X sky130_fd_sc_hd__buf_4
XFILLER_60_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26566_ _24911_/X _33722_/Q _26572_/S VGND VGND VPWR VPWR _26567_/A sky130_fd_sc_hd__mux2_1
X_23778_ _22990_/X _32375_/Q _23790_/S VGND VGND VPWR VPWR _23779_/A sky130_fd_sc_hd__mux2_1
XFILLER_220_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28305_ _27729_/X _34482_/Q _28307_/S VGND VGND VPWR VPWR _28306_/A sky130_fd_sc_hd__mux2_1
X_25517_ _25517_/A VGND VGND VPWR VPWR _33225_/D sky130_fd_sc_hd__clkbuf_1
X_22729_ _33681_/Q _33617_/Q _33553_/Q _33489_/Q _22506_/X _22507_/X VGND VGND VPWR
+ VPWR _22729_/X sky130_fd_sc_hd__mux4_1
XFILLER_241_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29285_ _34945_/Q _27168_/X _29297_/S VGND VGND VPWR VPWR _29286_/A sky130_fd_sc_hd__mux2_1
X_26497_ _24809_/X _33689_/Q _26509_/S VGND VGND VPWR VPWR _26498_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16250_ _16246_/X _16249_/X _16015_/X VGND VGND VPWR VPWR _16274_/A sky130_fd_sc_hd__o21ba_1
X_28236_ _28236_/A VGND VGND VPWR VPWR _34449_/D sky130_fd_sc_hd__clkbuf_1
X_25448_ _24858_/X _33193_/Q _25448_/S VGND VGND VPWR VPWR _25449_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16181_ _33369_/Q _33305_/Q _33241_/Q _33177_/Q _16002_/X _16003_/X VGND VGND VPWR
+ VPWR _16181_/X sky130_fd_sc_hd__mux4_1
XFILLER_142_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25379_ _33161_/Q _23460_/X _25395_/S VGND VGND VPWR VPWR _25380_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28167_ _28167_/A VGND VGND VPWR VPWR _34416_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27118_ input20/X VGND VGND VPWR VPWR _27118_/X sky130_fd_sc_hd__buf_2
X_28098_ _34384_/Q _27214_/X _28100_/S VGND VGND VPWR VPWR _28099_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27049_ _27049_/A VGND VGND VPWR VPWR _33946_/D sky130_fd_sc_hd__clkbuf_1
X_19940_ _19651_/X _19938_/X _19939_/X _19654_/X VGND VGND VPWR VPWR _19940_/X sky130_fd_sc_hd__a22o_1
XFILLER_181_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30060_ _30060_/A VGND VGND VPWR VPWR _35282_/D sky130_fd_sc_hd__clkbuf_1
X_19871_ _19867_/X _19870_/X _19793_/X _19794_/X VGND VGND VPWR VPWR _19888_/B sky130_fd_sc_hd__o211a_1
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1054 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18822_ _18747_/X _18820_/X _18821_/X _18750_/X VGND VGND VPWR VPWR _18822_/X sky130_fd_sc_hd__a22o_1
XTAP_6150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18753_ _34400_/Q _36128_/Q _34272_/Q _34208_/Q _18470_/X _18471_/X VGND VGND VPWR
+ VPWR _18753_/X sky130_fd_sc_hd__mux4_2
XFILLER_7_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17704_ _17859_/A VGND VGND VPWR VPWR _17704_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_110_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33750_ _36054_/CLK _33750_/D VGND VGND VPWR VPWR _33750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30962_ _31010_/S VGND VGND VPWR VPWR _30981_/S sky130_fd_sc_hd__buf_6
X_18684_ _18684_/A _18684_/B _18684_/C _18684_/D VGND VGND VPWR VPWR _18685_/A sky130_fd_sc_hd__or4_4
XFILLER_97_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32701_ _32891_/CLK _32701_/D VGND VGND VPWR VPWR _32701_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17635_ _32898_/Q _32834_/Q _32770_/Q _32706_/Q _17346_/X _17347_/X VGND VGND VPWR
+ VPWR _17635_/X sky130_fd_sc_hd__mux4_1
XFILLER_236_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33681_ _34441_/CLK _33681_/D VGND VGND VPWR VPWR _33681_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30893_ _35677_/Q input62/X _30897_/S VGND VGND VPWR VPWR _30894_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35420_ _35804_/CLK _35420_/D VGND VGND VPWR VPWR _35420_/Q sky130_fd_sc_hd__dfxtp_1
X_32632_ _36025_/CLK _32632_/D VGND VGND VPWR VPWR _32632_/Q sky130_fd_sc_hd__dfxtp_1
X_17566_ _33152_/Q _36032_/Q _33024_/Q _32960_/Q _17415_/X _17416_/X VGND VGND VPWR
+ VPWR _17566_/X sky130_fd_sc_hd__mux4_1
XFILLER_223_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19305_ _33072_/Q _32048_/Q _35824_/Q _35760_/Q _19025_/X _19026_/X VGND VGND VPWR
+ VPWR _19305_/X sky130_fd_sc_hd__mux4_2
X_35351_ _35799_/CLK _35351_/D VGND VGND VPWR VPWR _35351_/Q sky130_fd_sc_hd__dfxtp_1
X_16517_ _33058_/Q _32034_/Q _35810_/Q _35746_/Q _16372_/X _16373_/X VGND VGND VPWR
+ VPWR _16517_/X sky130_fd_sc_hd__mux4_1
X_32563_ _35955_/CLK _32563_/D VGND VGND VPWR VPWR _32563_/Q sky130_fd_sc_hd__dfxtp_1
X_17497_ _17850_/A VGND VGND VPWR VPWR _17497_/X sky130_fd_sc_hd__buf_4
XFILLER_147_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34302_ _36103_/CLK _34302_/D VGND VGND VPWR VPWR _34302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31514_ _27782_/X _35971_/Q _31522_/S VGND VGND VPWR VPWR _31515_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19236_ _33070_/Q _32046_/Q _35822_/Q _35758_/Q _19025_/X _19026_/X VGND VGND VPWR
+ VPWR _19236_/X sky130_fd_sc_hd__mux4_1
X_35282_ _35666_/CLK _35282_/D VGND VGND VPWR VPWR _35282_/Q sky130_fd_sc_hd__dfxtp_1
X_16448_ _34656_/Q _34592_/Q _34528_/Q _34464_/Q _16233_/X _16234_/X VGND VGND VPWR
+ VPWR _16448_/X sky130_fd_sc_hd__mux4_1
X_32494_ _35951_/CLK _32494_/D VGND VGND VPWR VPWR _32494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34233_ _36152_/CLK _34233_/D VGND VGND VPWR VPWR _34233_/Q sky130_fd_sc_hd__dfxtp_1
X_31445_ _27680_/X _35938_/Q _31459_/S VGND VGND VPWR VPWR _31446_/A sky130_fd_sc_hd__mux2_1
X_19167_ _35628_/Q _34988_/Q _34348_/Q _33708_/Q _19091_/X _19092_/X VGND VGND VPWR
+ VPWR _19167_/X sky130_fd_sc_hd__mux4_1
X_16379_ _16078_/X _16377_/X _16378_/X _16088_/X VGND VGND VPWR VPWR _16379_/X sky130_fd_sc_hd__a22o_1
XFILLER_30_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_91_CLK clkbuf_leaf_96_CLK/A VGND VGND VPWR VPWR _35551_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_219_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18118_ _16001_/X _18116_/X _18117_/X _16007_/X VGND VGND VPWR VPWR _18118_/X sky130_fd_sc_hd__a22o_1
XFILLER_121_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34164_ _34166_/CLK _34164_/D VGND VGND VPWR VPWR _34164_/Q sky130_fd_sc_hd__dfxtp_1
X_31376_ _31376_/A VGND VGND VPWR VPWR _35905_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19098_ _20157_/A VGND VGND VPWR VPWR _19098_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_69_1438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33115_ _35997_/CLK _33115_/D VGND VGND VPWR VPWR _33115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30327_ _35409_/Q _29512_/X _30327_/S VGND VGND VPWR VPWR _30328_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18049_ _32142_/Q _32334_/Q _32398_/Q _35918_/Q _17986_/X _17774_/X VGND VGND VPWR
+ VPWR _18049_/X sky130_fd_sc_hd__mux4_1
XFILLER_133_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34095_ _34991_/CLK _34095_/D VGND VGND VPWR VPWR _34095_/Q sky130_fd_sc_hd__dfxtp_1
X_33046_ _36119_/CLK _33046_/D VGND VGND VPWR VPWR _33046_/Q sky130_fd_sc_hd__dfxtp_1
X_21060_ _21051_/X _21058_/X _21059_/X VGND VGND VPWR VPWR _21061_/D sky130_fd_sc_hd__o21ba_1
X_30258_ _35376_/Q _29410_/X _30264_/S VGND VGND VPWR VPWR _30259_/A sky130_fd_sc_hd__mux2_1
XFILLER_235_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_904 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20011_ _33092_/Q _32068_/Q _35844_/Q _35780_/Q _19731_/X _19732_/X VGND VGND VPWR
+ VPWR _20011_/X sky130_fd_sc_hd__mux4_1
XFILLER_48_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1048 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30189_ _30189_/A VGND VGND VPWR VPWR _35343_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_235_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34997_ _35446_/CLK _34997_/D VGND VGND VPWR VPWR _34997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24750_ _24750_/A VGND VGND VPWR VPWR _32895_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33948_ _36211_/CLK _33948_/D VGND VGND VPWR VPWR _33948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21962_ _34682_/Q _34618_/Q _34554_/Q _34490_/Q _21892_/X _21893_/X VGND VGND VPWR
+ VPWR _21962_/X sky130_fd_sc_hd__mux4_1
XFILLER_55_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23701_ _23701_/A VGND VGND VPWR VPWR _32340_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_227_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20913_ _20913_/A VGND VGND VPWR VPWR _36188_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24681_ _22915_/X _32863_/Q _24681_/S VGND VGND VPWR VPWR _24682_/A sky130_fd_sc_hd__mux2_1
X_33879_ _34007_/CLK _33879_/D VGND VGND VPWR VPWR _33879_/Q sky130_fd_sc_hd__dfxtp_1
X_21893_ _22599_/A VGND VGND VPWR VPWR _21893_/X sky130_fd_sc_hd__buf_6
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26420_ _33653_/Q _23393_/X _26436_/S VGND VGND VPWR VPWR _26421_/A sky130_fd_sc_hd__mux2_1
X_35618_ _35618_/CLK _35618_/D VGND VGND VPWR VPWR _35618_/Q sky130_fd_sc_hd__dfxtp_1
X_23632_ _23632_/A VGND VGND VPWR VPWR _32307_/D sky130_fd_sc_hd__clkbuf_1
X_20844_ _33627_/Q _33563_/Q _33499_/Q _33435_/Q _20741_/X _20742_/X VGND VGND VPWR
+ VPWR _20844_/X sky130_fd_sc_hd__mux4_1
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_20_0_CLK clkbuf_2_2_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_20_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_54_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_214_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26351_ _26351_/A VGND VGND VPWR VPWR _33621_/D sky130_fd_sc_hd__clkbuf_1
X_23563_ _32276_/Q _23495_/X _23565_/S VGND VGND VPWR VPWR _23564_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35549_ _35613_/CLK _35549_/D VGND VGND VPWR VPWR _35549_/Q sky130_fd_sc_hd__dfxtp_1
X_20775_ _20769_/X _20774_/X _20704_/X VGND VGND VPWR VPWR _20776_/D sky130_fd_sc_hd__o21ba_1
XFILLER_39_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25302_ _25302_/A VGND VGND VPWR VPWR _33124_/D sky130_fd_sc_hd__clkbuf_1
X_22514_ _33930_/Q _33866_/Q _33802_/Q _36106_/Q _22330_/X _22331_/X VGND VGND VPWR
+ VPWR _22514_/X sky130_fd_sc_hd__mux4_1
X_29070_ _34843_/Q _27050_/X _29078_/S VGND VGND VPWR VPWR _29071_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26282_ _24892_/X _33588_/Q _26300_/S VGND VGND VPWR VPWR _26283_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23494_ _23494_/A VGND VGND VPWR VPWR _32243_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25233_ _25233_/A VGND VGND VPWR VPWR _33092_/D sky130_fd_sc_hd__clkbuf_1
X_28021_ _34347_/Q _27100_/X _28037_/S VGND VGND VPWR VPWR _28022_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22445_ _22373_/X _22443_/X _22444_/X _22377_/X VGND VGND VPWR VPWR _22445_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_82_CLK clkbuf_leaf_88_CLK/A VGND VGND VPWR VPWR _35805_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_13_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25164_ _25164_/A VGND VGND VPWR VPWR _33059_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22376_ _32902_/Q _32838_/Q _32774_/Q _32710_/Q _22299_/X _22300_/X VGND VGND VPWR
+ VPWR _22376_/X sky130_fd_sc_hd__mux4_1
XFILLER_100_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24115_ _31418_/A VGND VGND VPWR VPWR _24118_/A sky130_fd_sc_hd__inv_2
XFILLER_151_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21327_ _33064_/Q _32040_/Q _35816_/Q _35752_/Q _21325_/X _21326_/X VGND VGND VPWR
+ VPWR _21327_/X sky130_fd_sc_hd__mux4_1
X_25095_ _24942_/X _33028_/Q _25101_/S VGND VGND VPWR VPWR _25096_/A sky130_fd_sc_hd__mux2_1
X_29972_ _29972_/A VGND VGND VPWR VPWR _35240_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28923_ _29797_/A _31147_/B VGND VGND VPWR VPWR _29056_/S sky130_fd_sc_hd__nor2_8
X_24046_ _24046_/A VGND VGND VPWR VPWR _32564_/D sky130_fd_sc_hd__clkbuf_1
X_21258_ _21611_/A VGND VGND VPWR VPWR _21258_/X sky130_fd_sc_hd__buf_4
XFILLER_81_1104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_1224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20209_ _34186_/Q _34122_/Q _34058_/Q _33994_/Q _20099_/X _20100_/X VGND VGND VPWR
+ VPWR _20209_/X sky130_fd_sc_hd__mux4_1
X_28854_ _28854_/A VGND VGND VPWR VPWR _34740_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21189_ _35172_/Q _35108_/Q _35044_/Q _32164_/Q _20904_/X _20905_/X VGND VGND VPWR
+ VPWR _21189_/X sky130_fd_sc_hd__mux4_1
XFILLER_172_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27805_ _27804_/X _34250_/Q _27826_/S VGND VGND VPWR VPWR _27806_/A sky130_fd_sc_hd__mux2_1
XFILLER_131_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28785_ _28785_/A VGND VGND VPWR VPWR _34709_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25997_ _24871_/X _33453_/Q _26009_/S VGND VGND VPWR VPWR _25998_/A sky130_fd_sc_hd__mux2_1
XTAP_4033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27736_ _27838_/S VGND VGND VPWR VPWR _27764_/S sky130_fd_sc_hd__clkbuf_8
XTAP_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24948_ input43/X VGND VGND VPWR VPWR _24948_/X sky130_fd_sc_hd__buf_4
XTAP_4066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_246_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_935 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27667_ input63/X VGND VGND VPWR VPWR _27667_/X sky130_fd_sc_hd__buf_4
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24879_ _24879_/A VGND VGND VPWR VPWR _32943_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17420_ _17912_/A VGND VGND VPWR VPWR _17420_/X sky130_fd_sc_hd__clkbuf_4
X_29406_ _29406_/A VGND VGND VPWR VPWR _34990_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26618_ _24988_/X _33747_/Q _26622_/S VGND VGND VPWR VPWR _26619_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27598_ _34178_/Q _27171_/X _27608_/S VGND VGND VPWR VPWR _27599_/A sky130_fd_sc_hd__mux2_1
XFILLER_205_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29337_ _34968_/Q _29336_/X _29358_/S VGND VGND VPWR VPWR _29338_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17351_ _17859_/A VGND VGND VPWR VPWR _17351_/X sky130_fd_sc_hd__buf_6
X_26549_ _24886_/X _33714_/Q _26551_/S VGND VGND VPWR VPWR _26550_/A sky130_fd_sc_hd__mux2_1
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ _16296_/X _16301_/X _16075_/X VGND VGND VPWR VPWR _16312_/C sky130_fd_sc_hd__o21ba_1
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29268_ _34937_/Q _27143_/X _29276_/S VGND VGND VPWR VPWR _29269_/A sky130_fd_sc_hd__mux2_1
X_17282_ _32888_/Q _32824_/Q _32760_/Q _32696_/Q _16993_/X _16994_/X VGND VGND VPWR
+ VPWR _17282_/X sky130_fd_sc_hd__mux4_1
XFILLER_158_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19021_ _35688_/Q _32195_/Q _35560_/Q _35496_/Q _18911_/X _18912_/X VGND VGND VPWR
+ VPWR _19021_/X sky130_fd_sc_hd__mux4_1
X_28219_ _27801_/X _34441_/Q _28235_/S VGND VGND VPWR VPWR _28220_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16233_ _17998_/A VGND VGND VPWR VPWR _16233_/X sky130_fd_sc_hd__buf_6
X_29199_ _34904_/Q _27041_/X _29213_/S VGND VGND VPWR VPWR _29200_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_73_CLK clkbuf_leaf_73_CLK/A VGND VGND VPWR VPWR _36053_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_10_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31230_ _31230_/A VGND VGND VPWR VPWR _35836_/D sky130_fd_sc_hd__clkbuf_1
X_16164_ _33048_/Q _32024_/Q _35800_/Q _35736_/Q _16067_/X _16069_/X VGND VGND VPWR
+ VPWR _16164_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_6_18__f_CLK clkbuf_5_9_0_CLK/X VGND VGND VPWR VPWR clkbuf_leaf_88_CLK/A sky130_fd_sc_hd__clkbuf_16
XFILLER_126_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16095_ _34390_/Q _36118_/Q _34262_/Q _34198_/Q _16092_/X _16094_/X VGND VGND VPWR
+ VPWR _16095_/X sky130_fd_sc_hd__mux4_1
XFILLER_182_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31161_ _31161_/A VGND VGND VPWR VPWR _35803_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19923_ _34178_/Q _34114_/Q _34050_/Q _33986_/Q _19746_/X _19747_/X VGND VGND VPWR
+ VPWR _19923_/X sky130_fd_sc_hd__mux4_1
XFILLER_181_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30112_ _30112_/A VGND VGND VPWR VPWR _35306_/D sky130_fd_sc_hd__clkbuf_1
X_31092_ _31092_/A VGND VGND VPWR VPWR _35771_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30043_ _35274_/Q _29491_/X _30057_/S VGND VGND VPWR VPWR _30044_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_1414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34920_ _34920_/CLK _34920_/D VGND VGND VPWR VPWR _34920_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19854_ _20207_/A VGND VGND VPWR VPWR _19854_/X sky130_fd_sc_hd__buf_4
XFILLER_68_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18805_ _18799_/X _18804_/X _18726_/X VGND VGND VPWR VPWR _18829_/A sky130_fd_sc_hd__o21ba_1
XFILLER_95_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34851_ _34918_/CLK _34851_/D VGND VGND VPWR VPWR _34851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19785_ _20138_/A VGND VGND VPWR VPWR _19785_/X sky130_fd_sc_hd__clkbuf_4
X_16997_ _16991_/X _16996_/X _16787_/X _16788_/X VGND VGND VPWR VPWR _17018_/B sky130_fd_sc_hd__o211a_1
X_33802_ _36105_/CLK _33802_/D VGND VGND VPWR VPWR _33802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18736_ _18730_/X _18733_/X _18734_/X _18735_/X VGND VGND VPWR VPWR _18761_/B sky130_fd_sc_hd__o211a_1
XFILLER_3_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34782_ _36242_/CLK _34782_/D VGND VGND VPWR VPWR _34782_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31994_ _34405_/CLK _31994_/D VGND VGND VPWR VPWR _31994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33733_ _35717_/CLK _33733_/D VGND VGND VPWR VPWR _33733_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_1103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18667_ _18660_/X _18666_/X _18344_/X _18346_/X VGND VGND VPWR VPWR _18684_/B sky130_fd_sc_hd__o211a_1
X_30945_ _30945_/A VGND VGND VPWR VPWR _35701_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17618_ _17511_/X _17616_/X _17617_/X _17516_/X VGND VGND VPWR VPWR _17618_/X sky130_fd_sc_hd__a22o_1
XFILLER_240_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33664_ _33984_/CLK _33664_/D VGND VGND VPWR VPWR _33664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30876_ _30876_/A VGND VGND VPWR VPWR _35669_/D sky130_fd_sc_hd__clkbuf_1
X_18598_ _35420_/Q _35356_/Q _35292_/Q _35228_/Q _18495_/X _18496_/X VGND VGND VPWR
+ VPWR _18598_/X sky130_fd_sc_hd__mux4_1
X_35403_ _35596_/CLK _35403_/D VGND VGND VPWR VPWR _35403_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32615_ _35943_/CLK _32615_/D VGND VGND VPWR VPWR _32615_/Q sky130_fd_sc_hd__dfxtp_1
X_17549_ _17545_/X _17548_/X _17518_/X VGND VGND VPWR VPWR _17550_/D sky130_fd_sc_hd__o21ba_1
XFILLER_189_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33595_ _36093_/CLK _33595_/D VGND VGND VPWR VPWR _33595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35334_ _35466_/CLK _35334_/D VGND VGND VPWR VPWR _35334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_225_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20560_ _32917_/Q _32853_/Q _32789_/Q _32725_/Q _18284_/X _18287_/X VGND VGND VPWR
+ VPWR _20560_/X sky130_fd_sc_hd__mux4_1
X_32546_ _33119_/CLK _32546_/D VGND VGND VPWR VPWR _32546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19219_ _33390_/Q _33326_/Q _33262_/Q _33198_/Q _19074_/X _19075_/X VGND VGND VPWR
+ VPWR _19219_/X sky130_fd_sc_hd__mux4_1
X_35265_ _35458_/CLK _35265_/D VGND VGND VPWR VPWR _35265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20491_ _20205_/X _20489_/X _20490_/X _20210_/X VGND VGND VPWR VPWR _20491_/X sky130_fd_sc_hd__a22o_1
X_32477_ _35998_/CLK _32477_/D VGND VGND VPWR VPWR _32477_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_508_CLK clkbuf_leaf_2_CLK/A VGND VGND VPWR VPWR _34148_/CLK sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_64_CLK clkbuf_leaf_65_CLK/A VGND VGND VPWR VPWR _35922_/CLK sky130_fd_sc_hd__clkbuf_16
X_22230_ _32642_/Q _32578_/Q _32514_/Q _35970_/Q _22229_/X _22013_/X VGND VGND VPWR
+ VPWR _22230_/X sky130_fd_sc_hd__mux4_1
X_34216_ _36136_/CLK _34216_/D VGND VGND VPWR VPWR _34216_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31428_ _27655_/X _35930_/Q _31438_/S VGND VGND VPWR VPWR _31429_/A sky130_fd_sc_hd__mux2_1
X_35196_ _35645_/CLK _35196_/D VGND VGND VPWR VPWR _35196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22161_ _33920_/Q _33856_/Q _33792_/Q _36096_/Q _21977_/X _21978_/X VGND VGND VPWR
+ VPWR _22161_/X sky130_fd_sc_hd__mux4_1
X_34147_ _34148_/CLK _34147_/D VGND VGND VPWR VPWR _34147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31359_ _31359_/A VGND VGND VPWR VPWR _35897_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21112_ _21108_/X _21111_/X _21034_/X _21035_/X VGND VGND VPWR VPWR _21129_/B sky130_fd_sc_hd__o211a_1
XTAP_6908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34078_ _36205_/CLK _34078_/D VGND VGND VPWR VPWR _34078_/Q sky130_fd_sc_hd__dfxtp_1
X_22092_ _22020_/X _22090_/X _22091_/X _22024_/X VGND VGND VPWR VPWR _22092_/X sky130_fd_sc_hd__a22o_1
XTAP_6919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_1004 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25920_ _25920_/A VGND VGND VPWR VPWR _33416_/D sky130_fd_sc_hd__clkbuf_1
X_33029_ _35779_/CLK _33029_/D VGND VGND VPWR VPWR _33029_/Q sky130_fd_sc_hd__dfxtp_1
X_21043_ _33056_/Q _32032_/Q _35808_/Q _35744_/Q _20972_/X _20973_/X VGND VGND VPWR
+ VPWR _21043_/X sky130_fd_sc_hd__mux4_1
XFILLER_115_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25851_ _24855_/X _33384_/Q _25853_/S VGND VGND VPWR VPWR _25852_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24802_ _24802_/A VGND VGND VPWR VPWR _32918_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_189_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28570_ _28570_/A VGND VGND VPWR VPWR _34607_/D sky130_fd_sc_hd__clkbuf_1
X_25782_ _25782_/A VGND VGND VPWR VPWR _33351_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22994_ _22993_/X _32056_/Q _23009_/S VGND VGND VPWR VPWR _22995_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27521_ _27521_/A VGND VGND VPWR VPWR _34141_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21945_ _32122_/Q _32314_/Q _32378_/Q _35898_/Q _21880_/X _21668_/X VGND VGND VPWR
+ VPWR _21945_/X sky130_fd_sc_hd__mux4_1
X_24733_ _24733_/A VGND VGND VPWR VPWR _32887_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24664_ _24664_/A VGND VGND VPWR VPWR _32854_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27452_ _34109_/Q _27155_/X _27452_/S VGND VGND VPWR VPWR _27453_/A sky130_fd_sc_hd__mux2_1
XFILLER_242_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21876_ _22582_/A VGND VGND VPWR VPWR _21876_/X sky130_fd_sc_hd__buf_6
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26403_ _33645_/Q _23302_/X _26415_/S VGND VGND VPWR VPWR _26404_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23615_ _22953_/X _32299_/Q _23631_/S VGND VGND VPWR VPWR _23616_/A sky130_fd_sc_hd__mux2_1
X_20827_ _35610_/Q _34970_/Q _34330_/Q _33690_/Q _20653_/X _20655_/X VGND VGND VPWR
+ VPWR _20827_/X sky130_fd_sc_hd__mux4_1
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27383_ _34076_/Q _27053_/X _27389_/S VGND VGND VPWR VPWR _27384_/A sky130_fd_sc_hd__mux2_1
X_24595_ _22987_/X _32822_/Q _24609_/S VGND VGND VPWR VPWR _24596_/A sky130_fd_sc_hd__mux2_1
XFILLER_202_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29122_ _29191_/S VGND VGND VPWR VPWR _29141_/S sky130_fd_sc_hd__buf_4
X_26334_ _24970_/X _33613_/Q _26342_/S VGND VGND VPWR VPWR _26335_/A sky130_fd_sc_hd__mux2_1
X_23546_ _23546_/A VGND VGND VPWR VPWR _32267_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20758_ _20630_/X _20756_/X _20757_/X _20641_/X VGND VGND VPWR VPWR _20758_/X sky130_fd_sc_hd__a22o_1
XFILLER_211_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29053_ _29053_/A VGND VGND VPWR VPWR _34835_/D sky130_fd_sc_hd__clkbuf_1
X_26265_ _24868_/X _33580_/Q _26279_/S VGND VGND VPWR VPWR _26266_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23477_ _23477_/A VGND VGND VPWR VPWR _32237_/D sky130_fd_sc_hd__clkbuf_1
X_20689_ _20678_/X _20681_/X _20686_/X _20688_/X VGND VGND VPWR VPWR _20689_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_55_CLK clkbuf_leaf_57_CLK/A VGND VGND VPWR VPWR _32871_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_137_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28004_ _34339_/Q _27075_/X _28016_/S VGND VGND VPWR VPWR _28005_/A sky130_fd_sc_hd__mux2_1
X_25216_ _25216_/A VGND VGND VPWR VPWR _33084_/D sky130_fd_sc_hd__clkbuf_1
X_22428_ _22428_/A _22428_/B _22428_/C _22428_/D VGND VGND VPWR VPWR _22429_/A sky130_fd_sc_hd__or4_4
XFILLER_137_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26196_ _26196_/A VGND VGND VPWR VPWR _33547_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25147_ _25147_/A VGND VGND VPWR VPWR _33051_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22359_ _34182_/Q _34118_/Q _34054_/Q _33990_/Q _22046_/X _22047_/X VGND VGND VPWR
+ VPWR _22359_/X sky130_fd_sc_hd__mux4_1
XFILLER_178_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25078_ _24917_/X _33020_/Q _25080_/S VGND VGND VPWR VPWR _25079_/A sky130_fd_sc_hd__mux2_1
X_29955_ _35232_/Q _29360_/X _29973_/S VGND VGND VPWR VPWR _29956_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28906_ _28906_/A VGND VGND VPWR VPWR _34765_/D sky130_fd_sc_hd__clkbuf_1
X_16920_ _33902_/Q _33838_/Q _33774_/Q _36078_/Q _16671_/X _16672_/X VGND VGND VPWR
+ VPWR _16920_/X sky130_fd_sc_hd__mux4_1
X_24029_ _24029_/A VGND VGND VPWR VPWR _32556_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_219_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29886_ _29886_/A VGND VGND VPWR VPWR _35199_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16851_ _17910_/A VGND VGND VPWR VPWR _16851_/X sky130_fd_sc_hd__clkbuf_4
X_28837_ _28837_/A VGND VGND VPWR VPWR _34732_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19570_ _34168_/Q _34104_/Q _34040_/Q _33976_/Q _19393_/X _19394_/X VGND VGND VPWR
+ VPWR _19570_/X sky130_fd_sc_hd__mux4_1
XFILLER_213_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28768_ _34701_/Q _27205_/X _28776_/S VGND VGND VPWR VPWR _28769_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16782_ _33130_/Q _36010_/Q _33002_/Q _32938_/Q _16709_/X _16710_/X VGND VGND VPWR
+ VPWR _16782_/X sky130_fd_sc_hd__mux4_1
XFILLER_234_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18521_ _20286_/A VGND VGND VPWR VPWR _18521_/X sky130_fd_sc_hd__buf_6
X_27719_ _27719_/A VGND VGND VPWR VPWR _34222_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28699_ _34668_/Q _27103_/X _28713_/S VGND VGND VPWR VPWR _28700_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30730_ _35600_/Q _29509_/X _30732_/S VGND VGND VPWR VPWR _30731_/A sky130_fd_sc_hd__mux2_1
X_18452_ _18446_/X _18451_/X _18315_/X VGND VGND VPWR VPWR _18476_/A sky130_fd_sc_hd__o21ba_1
XFILLER_111_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17403_ _17403_/A _17403_/B _17403_/C _17403_/D VGND VGND VPWR VPWR _17404_/A sky130_fd_sc_hd__or4_4
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18383_ _20016_/A VGND VGND VPWR VPWR _18383_/X sky130_fd_sc_hd__clkbuf_8
X_30661_ _35567_/Q _29407_/X _30669_/S VGND VGND VPWR VPWR _30662_/A sky130_fd_sc_hd__mux2_1
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32400_ _35985_/CLK _32400_/D VGND VGND VPWR VPWR _32400_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ _17334_/A VGND VGND VPWR VPWR _31993_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_222_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33380_ _33828_/CLK _33380_/D VGND VGND VPWR VPWR _33380_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30592_ _30592_/A VGND VGND VPWR VPWR _35534_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32331_ _35980_/CLK _32331_/D VGND VGND VPWR VPWR _32331_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17265_ _17158_/X _17263_/X _17264_/X _17163_/X VGND VGND VPWR VPWR _17265_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_46_CLK clkbuf_leaf_49_CLK/A VGND VGND VPWR VPWR _35817_/CLK sky130_fd_sc_hd__clkbuf_16
X_19004_ _18800_/X _19002_/X _19003_/X _18803_/X VGND VGND VPWR VPWR _19004_/X sky130_fd_sc_hd__a22o_1
XFILLER_31_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16216_ _16212_/X _16215_/X _16015_/X VGND VGND VPWR VPWR _16242_/A sky130_fd_sc_hd__o21ba_1
X_35050_ _35434_/CLK _35050_/D VGND VGND VPWR VPWR _35050_/Q sky130_fd_sc_hd__dfxtp_1
X_32262_ _35718_/CLK _32262_/D VGND VGND VPWR VPWR _32262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17196_ _17192_/X _17195_/X _17165_/X VGND VGND VPWR VPWR _17197_/D sky130_fd_sc_hd__o21ba_1
XFILLER_128_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34001_ _34193_/CLK _34001_/D VGND VGND VPWR VPWR _34001_/Q sky130_fd_sc_hd__dfxtp_1
X_31213_ _27735_/X _35828_/Q _31231_/S VGND VGND VPWR VPWR _31214_/A sky130_fd_sc_hd__mux2_1
X_16147_ _17864_/A VGND VGND VPWR VPWR _16147_/X sky130_fd_sc_hd__buf_6
XFILLER_182_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32193_ _35687_/CLK _32193_/D VGND VGND VPWR VPWR _32193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31144_ _31144_/A VGND VGND VPWR VPWR _35796_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16078_ _17153_/A VGND VGND VPWR VPWR _16078_/X sky130_fd_sc_hd__buf_4
XFILLER_68_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19906_ _19651_/X _19904_/X _19905_/X _19654_/X VGND VGND VPWR VPWR _19906_/X sky130_fd_sc_hd__a22o_1
XFILLER_9_1324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31075_ _31075_/A VGND VGND VPWR VPWR _35763_/D sky130_fd_sc_hd__clkbuf_1
X_35952_ _35952_/CLK _35952_/D VGND VGND VPWR VPWR _35952_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34903_ _34903_/CLK _34903_/D VGND VGND VPWR VPWR _34903_/Q sky130_fd_sc_hd__dfxtp_1
X_30026_ _35266_/Q _29466_/X _30036_/S VGND VGND VPWR VPWR _30027_/A sky130_fd_sc_hd__mux2_1
X_19837_ _35647_/Q _35007_/Q _34367_/Q _33727_/Q _19797_/X _19798_/X VGND VGND VPWR
+ VPWR _19837_/X sky130_fd_sc_hd__mux4_1
XFILLER_69_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35883_ _35883_/CLK _35883_/D VGND VGND VPWR VPWR _35883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34834_ _34964_/CLK _34834_/D VGND VGND VPWR VPWR _34834_/Q sky130_fd_sc_hd__dfxtp_1
Xinput2 DW[10] VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__buf_6
X_19768_ _34685_/Q _34621_/Q _34557_/Q _34493_/Q _19592_/X _19593_/X VGND VGND VPWR
+ VPWR _19768_/X sky130_fd_sc_hd__mux4_1
XFILLER_209_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18719_ _34144_/Q _34080_/Q _34016_/Q _33952_/Q _18687_/X _18688_/X VGND VGND VPWR
+ VPWR _18719_/X sky130_fd_sc_hd__mux4_1
X_34765_ _34957_/CLK _34765_/D VGND VGND VPWR VPWR _34765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_232_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31977_ _34790_/CLK _31977_/D VGND VGND VPWR VPWR _31977_/Q sky130_fd_sc_hd__dfxtp_1
X_19699_ _34427_/Q _36155_/Q _34299_/Q _34235_/Q _19529_/X _19530_/X VGND VGND VPWR
+ VPWR _19699_/X sky130_fd_sc_hd__mux4_1
XFILLER_36_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21730_ _33908_/Q _33844_/Q _33780_/Q _36084_/Q _21624_/X _21625_/X VGND VGND VPWR
+ VPWR _21730_/X sky130_fd_sc_hd__mux4_1
X_33716_ _35701_/CLK _33716_/D VGND VGND VPWR VPWR _33716_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30928_ _30928_/A VGND VGND VPWR VPWR _35693_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34696_ _36113_/CLK _34696_/D VGND VGND VPWR VPWR _34696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33647_ _34035_/CLK _33647_/D VGND VGND VPWR VPWR _33647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21661_ _32626_/Q _32562_/Q _32498_/Q _35954_/Q _21523_/X _21660_/X VGND VGND VPWR
+ VPWR _21661_/X sky130_fd_sc_hd__mux4_1
X_30859_ _35661_/Q input51/X _30867_/S VGND VGND VPWR VPWR _30860_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23400_ _32212_/Q _23399_/X _23418_/S VGND VGND VPWR VPWR _23401_/A sky130_fd_sc_hd__mux2_1
X_20612_ _33878_/Q _33814_/Q _33750_/Q _36054_/Q _20609_/X _20611_/X VGND VGND VPWR
+ VPWR _20612_/X sky130_fd_sc_hd__mux4_1
XFILLER_36_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24380_ _24380_/A VGND VGND VPWR VPWR _32720_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_240_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33578_ _34153_/CLK _33578_/D VGND VGND VPWR VPWR _33578_/Q sky130_fd_sc_hd__dfxtp_1
X_21592_ _32112_/Q _32304_/Q _32368_/Q _35888_/Q _21527_/X _21315_/X VGND VGND VPWR
+ VPWR _21592_/X sky130_fd_sc_hd__mux4_1
XFILLER_193_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_1267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23331_ _32183_/Q _23252_/X _23335_/S VGND VGND VPWR VPWR _23332_/A sky130_fd_sc_hd__mux2_1
X_35317_ _35446_/CLK _35317_/D VGND VGND VPWR VPWR _35317_/Q sky130_fd_sc_hd__dfxtp_1
X_20543_ _34452_/Q _36180_/Q _34324_/Q _34260_/Q _18367_/X _18369_/X VGND VGND VPWR
+ VPWR _20543_/X sky130_fd_sc_hd__mux4_1
XFILLER_162_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32529_ _36049_/CLK _32529_/D VGND VGND VPWR VPWR _32529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_37_CLK clkbuf_6_7__f_CLK/X VGND VGND VPWR VPWR _35938_/CLK sky130_fd_sc_hd__clkbuf_16
X_26050_ _26050_/A VGND VGND VPWR VPWR _33478_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35248_ _35634_/CLK _35248_/D VGND VGND VPWR VPWR _35248_/Q sky130_fd_sc_hd__dfxtp_1
X_23262_ _23565_/S VGND VGND VPWR VPWR _23290_/S sky130_fd_sc_hd__buf_6
X_20474_ _35666_/Q _35026_/Q _34386_/Q _33746_/Q _18412_/X _18413_/X VGND VGND VPWR
+ VPWR _20474_/X sky130_fd_sc_hd__mux4_1
X_25001_ _24803_/X _32983_/Q _25017_/S VGND VGND VPWR VPWR _25002_/A sky130_fd_sc_hd__mux2_1
X_22213_ _34689_/Q _34625_/Q _34561_/Q _34497_/Q _21892_/X _21893_/X VGND VGND VPWR
+ VPWR _22213_/X sky130_fd_sc_hd__mux4_1
XFILLER_119_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_934 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23193_ _23193_/A VGND VGND VPWR VPWR _32134_/D sky130_fd_sc_hd__clkbuf_1
X_35179_ _35180_/CLK _35179_/D VGND VGND VPWR VPWR _35179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22144_ _35199_/Q _35135_/Q _35071_/Q _32255_/Q _21963_/X _21964_/X VGND VGND VPWR
+ VPWR _22144_/X sky130_fd_sc_hd__mux4_1
XFILLER_10_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29740_ _29740_/A VGND VGND VPWR VPWR _35130_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26952_ _33903_/Q _23316_/X _26960_/S VGND VGND VPWR VPWR _26953_/A sky130_fd_sc_hd__mux2_1
X_22075_ _22075_/A _22075_/B _22075_/C _22075_/D VGND VGND VPWR VPWR _22076_/A sky130_fd_sc_hd__or4_4
XTAP_6749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25903_ _25903_/A VGND VGND VPWR VPWR _33408_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21026_ _22438_/A VGND VGND VPWR VPWR _21026_/X sky130_fd_sc_hd__buf_4
XFILLER_86_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29671_ _29671_/A VGND VGND VPWR VPWR _35097_/D sky130_fd_sc_hd__clkbuf_1
X_26883_ _26883_/A VGND VGND VPWR VPWR _33870_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28622_ _27797_/X _34632_/Q _28640_/S VGND VGND VPWR VPWR _28623_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25834_ _25945_/S VGND VGND VPWR VPWR _25853_/S sky130_fd_sc_hd__buf_4
XFILLER_132_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28553_ _28553_/A VGND VGND VPWR VPWR _34599_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25765_ _24927_/X _33343_/Q _25781_/S VGND VGND VPWR VPWR _25766_/A sky130_fd_sc_hd__mux2_1
X_22977_ input22/X VGND VGND VPWR VPWR _22977_/X sky130_fd_sc_hd__buf_2
XFILLER_243_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27504_ _30877_/B _31688_/B VGND VGND VPWR VPWR _27637_/S sky130_fd_sc_hd__nor2_8
XFILLER_28_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24716_ _24716_/A VGND VGND VPWR VPWR _32879_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_215_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28484_ _27794_/X _34567_/Q _28484_/S VGND VGND VPWR VPWR _28485_/A sky130_fd_sc_hd__mux2_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21928_ _21753_/X _21926_/X _21927_/X _21756_/X VGND VGND VPWR VPWR _21928_/X sky130_fd_sc_hd__a22o_1
XFILLER_243_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25696_ _25696_/A VGND VGND VPWR VPWR _33310_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27435_ _27435_/A VGND VGND VPWR VPWR _34100_/D sky130_fd_sc_hd__clkbuf_1
X_24647_ _23064_/X _32847_/Q _24651_/S VGND VGND VPWR VPWR _24648_/A sky130_fd_sc_hd__mux2_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21859_ _21853_/X _21858_/X _21751_/X VGND VGND VPWR VPWR _21867_/C sky130_fd_sc_hd__o21ba_1
XFILLER_163_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27366_ _27366_/A VGND VGND VPWR VPWR _34068_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24578_ _22962_/X _32814_/Q _24588_/S VGND VGND VPWR VPWR _24579_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_875 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29105_ _29105_/A VGND VGND VPWR VPWR _34859_/D sky130_fd_sc_hd__clkbuf_1
X_26317_ _24945_/X _33605_/Q _26321_/S VGND VGND VPWR VPWR _26318_/A sky130_fd_sc_hd__mux2_1
X_23529_ _23529_/A VGND VGND VPWR VPWR _32259_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27297_ _27297_/A VGND VGND VPWR VPWR _34035_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_28_CLK clkbuf_6_5__f_CLK/X VGND VGND VPWR VPWR _36209_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_184_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29036_ _34827_/Q _27199_/X _29048_/S VGND VGND VPWR VPWR _29037_/A sky130_fd_sc_hd__mux2_1
X_17050_ _17050_/A _17050_/B _17050_/C _17050_/D VGND VGND VPWR VPWR _17051_/A sky130_fd_sc_hd__or4_4
X_26248_ _24843_/X _33572_/Q _26258_/S VGND VGND VPWR VPWR _26249_/A sky130_fd_sc_hd__mux2_1
X_16001_ _17864_/A VGND VGND VPWR VPWR _16001_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_87_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26179_ _26179_/A VGND VGND VPWR VPWR _33539_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_978 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29938_ _35224_/Q _29336_/X _29952_/S VGND VGND VPWR VPWR _29939_/A sky130_fd_sc_hd__mux2_1
X_17952_ _17765_/X _17950_/X _17951_/X _17771_/X VGND VGND VPWR VPWR _17952_/X sky130_fd_sc_hd__a22o_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16903_ _35437_/Q _35373_/Q _35309_/Q _35245_/Q _16901_/X _16902_/X VGND VGND VPWR
+ VPWR _16903_/X sky130_fd_sc_hd__mux4_1
XFILLER_239_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17883_ _33161_/Q _36041_/Q _33033_/Q _32969_/Q _17768_/X _17769_/X VGND VGND VPWR
+ VPWR _17883_/X sky130_fd_sc_hd__mux4_1
XFILLER_113_1406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29869_ _29869_/A VGND VGND VPWR VPWR _35191_/D sky130_fd_sc_hd__clkbuf_1
X_19622_ _35449_/Q _35385_/Q _35321_/Q _35257_/Q _19554_/X _19555_/X VGND VGND VPWR
+ VPWR _19622_/X sky130_fd_sc_hd__mux4_1
X_31900_ _23408_/X _36154_/Q _31906_/S VGND VGND VPWR VPWR _31901_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16834_ _33067_/Q _32043_/Q _35819_/Q _35755_/Q _16725_/X _16726_/X VGND VGND VPWR
+ VPWR _16834_/X sky130_fd_sc_hd__mux4_1
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32880_ _32906_/CLK _32880_/D VGND VGND VPWR VPWR _32880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31831_ _23240_/X _36121_/Q _31843_/S VGND VGND VPWR VPWR _31832_/A sky130_fd_sc_hd__mux2_1
X_19553_ _19298_/X _19551_/X _19552_/X _19301_/X VGND VGND VPWR VPWR _19553_/X sky130_fd_sc_hd__a22o_1
X_16765_ _34409_/Q _36137_/Q _34281_/Q _34217_/Q _16523_/X _16524_/X VGND VGND VPWR
+ VPWR _16765_/X sky130_fd_sc_hd__mux4_1
XFILLER_18_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18504_ _34393_/Q _36121_/Q _34265_/Q _34201_/Q _18470_/X _18471_/X VGND VGND VPWR
+ VPWR _18504_/X sky130_fd_sc_hd__mux4_1
XFILLER_18_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34550_ _36024_/CLK _34550_/D VGND VGND VPWR VPWR _34550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31762_ _31762_/A VGND VGND VPWR VPWR _36088_/D sky130_fd_sc_hd__clkbuf_1
X_19484_ _35637_/Q _34997_/Q _34357_/Q _33717_/Q _19444_/X _19445_/X VGND VGND VPWR
+ VPWR _19484_/X sky130_fd_sc_hd__mux4_1
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16696_ _16692_/X _16695_/X _16459_/X VGND VGND VPWR VPWR _16697_/D sky130_fd_sc_hd__o21ba_1
XFILLER_61_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33501_ _36191_/CLK _33501_/D VGND VGND VPWR VPWR _33501_/Q sky130_fd_sc_hd__dfxtp_1
X_18435_ _34903_/Q _34839_/Q _34775_/Q _34711_/Q _18396_/X _18398_/X VGND VGND VPWR
+ VPWR _18435_/X sky130_fd_sc_hd__mux4_1
XFILLER_206_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30713_ _30740_/S VGND VGND VPWR VPWR _30732_/S sky130_fd_sc_hd__buf_4
XFILLER_181_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34481_ _36143_/CLK _34481_/D VGND VGND VPWR VPWR _34481_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31693_ _31693_/A VGND VGND VPWR VPWR _36055_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36220_ _36223_/CLK _36220_/D VGND VGND VPWR VPWR _36220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33432_ _34009_/CLK _33432_/D VGND VGND VPWR VPWR _33432_/Q sky130_fd_sc_hd__dfxtp_1
X_18366_ _20282_/A VGND VGND VPWR VPWR _20235_/A sky130_fd_sc_hd__buf_12
X_30644_ _35559_/Q _29382_/X _30648_/S VGND VGND VPWR VPWR _30645_/A sky130_fd_sc_hd__mux2_1
XFILLER_222_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17317_ _17799_/A VGND VGND VPWR VPWR _17317_/X sky130_fd_sc_hd__buf_6
X_36151_ _36151_/CLK _36151_/D VGND VGND VPWR VPWR _36151_/Q sky130_fd_sc_hd__dfxtp_1
X_33363_ _36179_/CLK _33363_/D VGND VGND VPWR VPWR _33363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18297_ _18281_/X _18288_/X _18291_/X _18296_/X VGND VGND VPWR VPWR _18297_/X sky130_fd_sc_hd__a22o_1
X_30575_ _30575_/A VGND VGND VPWR VPWR _35526_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_19_CLK clkbuf_6_4__f_CLK/X VGND VGND VPWR VPWR _35490_/CLK sky130_fd_sc_hd__clkbuf_16
X_35102_ _36223_/CLK _35102_/D VGND VGND VPWR VPWR _35102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32314_ _35962_/CLK _32314_/D VGND VGND VPWR VPWR _32314_/Q sky130_fd_sc_hd__dfxtp_1
X_36082_ _36082_/CLK _36082_/D VGND VGND VPWR VPWR _36082_/Q sky130_fd_sc_hd__dfxtp_1
X_17248_ _32887_/Q _32823_/Q _32759_/Q _32695_/Q _16993_/X _16994_/X VGND VGND VPWR
+ VPWR _17248_/X sky130_fd_sc_hd__mux4_1
X_33294_ _36105_/CLK _33294_/D VGND VGND VPWR VPWR _33294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35033_ _35160_/CLK _35033_/D VGND VGND VPWR VPWR _35033_/Q sky130_fd_sc_hd__dfxtp_1
X_32245_ _35733_/CLK _32245_/D VGND VGND VPWR VPWR _32245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17179_ _32117_/Q _32309_/Q _32373_/Q _35893_/Q _16927_/X _17068_/X VGND VGND VPWR
+ VPWR _17179_/X sky130_fd_sc_hd__mux4_1
XFILLER_66_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20190_ _35657_/Q _35017_/Q _34377_/Q _33737_/Q _20150_/X _20151_/X VGND VGND VPWR
+ VPWR _20190_/X sky130_fd_sc_hd__mux4_1
XFILLER_157_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32176_ _34926_/CLK _32176_/D VGND VGND VPWR VPWR _32176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31127_ _35788_/Q input50/X _31137_/S VGND VGND VPWR VPWR _31128_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35935_ _35998_/CLK _35935_/D VGND VGND VPWR VPWR _35935_/Q sky130_fd_sc_hd__dfxtp_1
X_31058_ _35755_/Q input14/X _31074_/S VGND VGND VPWR VPWR _31059_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22900_ input45/X VGND VGND VPWR VPWR _22900_/X sky130_fd_sc_hd__buf_2
X_30009_ _35258_/Q _29441_/X _30015_/S VGND VGND VPWR VPWR _30010_/A sky130_fd_sc_hd__mux2_1
X_23880_ _23880_/A VGND VGND VPWR VPWR _32486_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_229_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35866_ _35994_/CLK _35866_/D VGND VGND VPWR VPWR _35866_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22831_ _21758_/A _22829_/X _22830_/X _21763_/A VGND VGND VPWR VPWR _22831_/X sky130_fd_sc_hd__a22o_1
XFILLER_72_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34817_ _36163_/CLK _34817_/D VGND VGND VPWR VPWR _34817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_244_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35797_ _36052_/CLK _35797_/D VGND VGND VPWR VPWR _35797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22762_ _33426_/Q _33362_/Q _33298_/Q _33234_/Q _20637_/X _20639_/X VGND VGND VPWR
+ VPWR _22762_/X sky130_fd_sc_hd__mux4_1
X_25550_ _24809_/X _33241_/Q _25562_/S VGND VGND VPWR VPWR _25551_/A sky130_fd_sc_hd__mux2_1
X_34748_ _36154_/CLK _34748_/D VGND VGND VPWR VPWR _34748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24501_ _24501_/A VGND VGND VPWR VPWR _32777_/D sky130_fd_sc_hd__clkbuf_1
X_21713_ _21603_/X _21711_/X _21712_/X _21606_/X VGND VGND VPWR VPWR _21713_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25481_ _25481_/A VGND VGND VPWR VPWR _33208_/D sky130_fd_sc_hd__clkbuf_1
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22693_ _34447_/Q _36175_/Q _34319_/Q _34255_/Q _22535_/X _22536_/X VGND VGND VPWR
+ VPWR _22693_/X sky130_fd_sc_hd__mux4_1
XFILLER_129_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34679_ _36150_/CLK _34679_/D VGND VGND VPWR VPWR _34679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_244_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27220_ input57/X VGND VGND VPWR VPWR _27220_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_52_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21644_ _35185_/Q _35121_/Q _35057_/Q _32198_/Q _21610_/X _21611_/X VGND VGND VPWR
+ VPWR _21644_/X sky130_fd_sc_hd__mux4_1
X_24432_ _22946_/X _32745_/Q _24432_/S VGND VGND VPWR VPWR _24433_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24363_ _23042_/X _32712_/Q _24381_/S VGND VGND VPWR VPWR _24364_/A sky130_fd_sc_hd__mux2_1
X_27151_ _27151_/A VGND VGND VPWR VPWR _33979_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21575_ _21400_/X _21573_/X _21574_/X _21403_/X VGND VGND VPWR VPWR _21575_/X sky130_fd_sc_hd__a22o_1
XFILLER_227_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23314_ _32175_/Q _23225_/X _23335_/S VGND VGND VPWR VPWR _23315_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26102_ _24827_/X _33503_/Q _26102_/S VGND VGND VPWR VPWR _26103_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20526_ _32660_/Q _32596_/Q _32532_/Q _35988_/Q _20282_/X _19177_/A VGND VGND VPWR
+ VPWR _20526_/X sky130_fd_sc_hd__mux4_1
X_27082_ _33957_/Q _27081_/X _27094_/S VGND VGND VPWR VPWR _27083_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24294_ _24294_/A VGND VGND VPWR VPWR _32679_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23245_ _23245_/A VGND VGND VPWR VPWR _32154_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26033_ _24923_/X _33470_/Q _26051_/S VGND VGND VPWR VPWR _26034_/A sky130_fd_sc_hd__mux2_1
XFILLER_238_1110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20457_ _20457_/A _20457_/B _20457_/C _20457_/D VGND VGND VPWR VPWR _20458_/A sky130_fd_sc_hd__or4_1
XFILLER_21_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23176_ _23011_/X _32126_/Q _23194_/S VGND VGND VPWR VPWR _23177_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20388_ _18301_/X _20386_/X _20387_/X _18307_/X VGND VGND VPWR VPWR _20388_/X sky130_fd_sc_hd__a22o_1
XFILLER_238_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22127_ _21806_/X _22125_/X _22126_/X _21809_/X VGND VGND VPWR VPWR _22127_/X sky130_fd_sc_hd__a22o_1
XTAP_6524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27984_ _27984_/A VGND VGND VPWR VPWR _34329_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput180 _36215_/Q VGND VGND VPWR VPWR D2[33] sky130_fd_sc_hd__buf_2
XFILLER_248_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput191 _36225_/Q VGND VGND VPWR VPWR D2[43] sky130_fd_sc_hd__buf_2
XTAP_5812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29723_ _29723_/A VGND VGND VPWR VPWR _35122_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22058_ _32893_/Q _32829_/Q _32765_/Q _32701_/Q _21946_/X _21947_/X VGND VGND VPWR
+ VPWR _22058_/X sky130_fd_sc_hd__mux4_1
X_26935_ _33895_/Q _23283_/X _26939_/S VGND VGND VPWR VPWR _26936_/A sky130_fd_sc_hd__mux2_1
XTAP_6579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21009_ _34655_/Q _34591_/Q _34527_/Q _34463_/Q _20833_/X _20834_/X VGND VGND VPWR
+ VPWR _21009_/X sky130_fd_sc_hd__mux4_1
XTAP_5867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29654_ _35090_/Q _29515_/X _29660_/S VGND VGND VPWR VPWR _29655_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26866_ _26866_/A VGND VGND VPWR VPWR _33862_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28605_ _27773_/X _34624_/Q _28619_/S VGND VGND VPWR VPWR _28606_/A sky130_fd_sc_hd__mux2_1
XFILLER_235_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25817_ _25817_/A VGND VGND VPWR VPWR _33367_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29585_ _35057_/Q _29413_/X _29589_/S VGND VGND VPWR VPWR _29586_/A sky130_fd_sc_hd__mux2_1
X_26797_ _26797_/A VGND VGND VPWR VPWR _33829_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28536_ _28536_/A VGND VGND VPWR VPWR _34591_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16550_ _35427_/Q _35363_/Q _35299_/Q _35235_/Q _16548_/X _16549_/X VGND VGND VPWR
+ VPWR _16550_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25748_ _24902_/X _33335_/Q _25760_/S VGND VGND VPWR VPWR _25749_/A sky130_fd_sc_hd__mux2_1
XFILLER_216_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_243_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28467_ _28467_/A VGND VGND VPWR VPWR _34558_/D sky130_fd_sc_hd__clkbuf_1
X_16481_ _33057_/Q _32033_/Q _35809_/Q _35745_/Q _16372_/X _16373_/X VGND VGND VPWR
+ VPWR _16481_/X sky130_fd_sc_hd__mux4_1
XFILLER_204_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25679_ _24796_/X _33302_/Q _25697_/S VGND VGND VPWR VPWR _25680_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18220_ _34196_/Q _34132_/Q _34068_/Q _34004_/Q _16049_/X _16050_/X VGND VGND VPWR
+ VPWR _18220_/X sky130_fd_sc_hd__mux4_1
XFILLER_223_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27418_ _27418_/A VGND VGND VPWR VPWR _34092_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_1120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28398_ _27667_/X _34526_/Q _28400_/S VGND VGND VPWR VPWR _28399_/A sky130_fd_sc_hd__mux2_1
XFILLER_203_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18151_ _35217_/Q _35153_/Q _35089_/Q _32273_/Q _16092_/X _16094_/X VGND VGND VPWR
+ VPWR _18151_/X sky130_fd_sc_hd__mux4_1
X_27349_ _34060_/Q _27202_/X _27359_/S VGND VGND VPWR VPWR _27350_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17102_ _33139_/Q _36019_/Q _33011_/Q _32947_/Q _17062_/X _17063_/X VGND VGND VPWR
+ VPWR _17102_/X sky130_fd_sc_hd__mux4_1
XFILLER_172_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18082_ _18078_/X _18081_/X _17846_/X _17847_/X VGND VGND VPWR VPWR _18097_/B sky130_fd_sc_hd__o211a_1
XFILLER_129_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30360_ _35424_/Q _29360_/X _30378_/S VGND VGND VPWR VPWR _30361_/A sky130_fd_sc_hd__mux2_1
XFILLER_200_996 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29019_ _34819_/Q _27174_/X _29027_/S VGND VGND VPWR VPWR _29020_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17033_ _32881_/Q _32817_/Q _32753_/Q _32689_/Q _16993_/X _16994_/X VGND VGND VPWR
+ VPWR _17033_/X sky130_fd_sc_hd__mux4_1
XFILLER_156_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30291_ _30291_/A VGND VGND VPWR VPWR _35391_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32030_ _35805_/CLK _32030_/D VGND VGND VPWR VPWR _32030_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18984_ _35623_/Q _34983_/Q _34343_/Q _33703_/Q _18738_/X _18739_/X VGND VGND VPWR
+ VPWR _18984_/X sky130_fd_sc_hd__mux4_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17935_ _17935_/A VGND VGND VPWR VPWR _17935_/X sky130_fd_sc_hd__buf_6
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33981_ _34877_/CLK _33981_/D VGND VGND VPWR VPWR _33981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_230_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35720_ _35721_/CLK _35720_/D VGND VGND VPWR VPWR _35720_/Q sky130_fd_sc_hd__dfxtp_1
X_32932_ _36005_/CLK _32932_/D VGND VGND VPWR VPWR _32932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17866_ _17866_/A VGND VGND VPWR VPWR _17866_/X sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_8_CLK clkbuf_leaf_9_CLK/A VGND VGND VPWR VPWR _34913_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_26_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19605_ _19499_/X _19603_/X _19604_/X _19504_/X VGND VGND VPWR VPWR _19605_/X sky130_fd_sc_hd__a22o_1
X_16817_ _34155_/Q _34091_/Q _34027_/Q _33963_/Q _16740_/X _16741_/X VGND VGND VPWR
+ VPWR _16817_/X sky130_fd_sc_hd__mux4_1
XFILLER_238_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35651_ _35651_/CLK _35651_/D VGND VGND VPWR VPWR _35651_/Q sky130_fd_sc_hd__dfxtp_1
X_32863_ _35870_/CLK _32863_/D VGND VGND VPWR VPWR _32863_/Q sky130_fd_sc_hd__dfxtp_1
X_17797_ _17797_/A VGND VGND VPWR VPWR _32006_/D sky130_fd_sc_hd__buf_4
XFILLER_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31814_ _31814_/A VGND VGND VPWR VPWR _36113_/D sky130_fd_sc_hd__clkbuf_1
X_19536_ _19536_/A VGND VGND VPWR VPWR _32438_/D sky130_fd_sc_hd__buf_2
X_34602_ _36140_/CLK _34602_/D VGND VGND VPWR VPWR _34602_/Q sky130_fd_sc_hd__dfxtp_1
X_35582_ _35713_/CLK _35582_/D VGND VGND VPWR VPWR _35582_/Q sky130_fd_sc_hd__dfxtp_1
X_16748_ _32617_/Q _32553_/Q _32489_/Q _35945_/Q _16570_/X _16707_/X VGND VGND VPWR
+ VPWR _16748_/X sky130_fd_sc_hd__mux4_1
X_32794_ _34070_/CLK _32794_/D VGND VGND VPWR VPWR _32794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34533_ _36136_/CLK _34533_/D VGND VGND VPWR VPWR _34533_/Q sky130_fd_sc_hd__dfxtp_1
X_31745_ _31745_/A VGND VGND VPWR VPWR _36080_/D sky130_fd_sc_hd__clkbuf_1
X_19467_ _19467_/A _19467_/B _19467_/C _19467_/D VGND VGND VPWR VPWR _19468_/A sky130_fd_sc_hd__or4_1
X_16679_ _32103_/Q _32295_/Q _32359_/Q _35879_/Q _16574_/X _16362_/X VGND VGND VPWR
+ VPWR _16679_/X sky130_fd_sc_hd__mux4_1
XFILLER_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1097 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18418_ _33111_/Q _35991_/Q _32983_/Q _32919_/Q _18324_/X _18325_/X VGND VGND VPWR
+ VPWR _18418_/X sky130_fd_sc_hd__mux4_1
X_34464_ _34594_/CLK _34464_/D VGND VGND VPWR VPWR _34464_/Q sky130_fd_sc_hd__dfxtp_1
X_31676_ _27822_/X _36048_/Q _31678_/S VGND VGND VPWR VPWR _31677_/A sky130_fd_sc_hd__mux2_1
X_19398_ _33907_/Q _33843_/Q _33779_/Q _36083_/Q _19324_/X _19325_/X VGND VGND VPWR
+ VPWR _19398_/X sky130_fd_sc_hd__mux4_1
XFILLER_72_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33415_ _33415_/CLK _33415_/D VGND VGND VPWR VPWR _33415_/Q sky130_fd_sc_hd__dfxtp_1
X_36203_ _36210_/CLK _36203_/D VGND VGND VPWR VPWR _36203_/Q sky130_fd_sc_hd__dfxtp_1
X_18349_ _20099_/A VGND VGND VPWR VPWR _18349_/X sky130_fd_sc_hd__buf_6
X_30627_ _35551_/Q _29357_/X _30627_/S VGND VGND VPWR VPWR _30628_/A sky130_fd_sc_hd__mux2_1
X_34395_ _35162_/CLK _34395_/D VGND VGND VPWR VPWR _34395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36134_ _36136_/CLK _36134_/D VGND VGND VPWR VPWR _36134_/Q sky130_fd_sc_hd__dfxtp_1
X_33346_ _36097_/CLK _33346_/D VGND VGND VPWR VPWR _33346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21360_ _21250_/X _21358_/X _21359_/X _21253_/X VGND VGND VPWR VPWR _21360_/X sky130_fd_sc_hd__a22o_1
XFILLER_175_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30558_ _35518_/Q _29453_/X _30576_/S VGND VGND VPWR VPWR _30559_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_826 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20311_ _20205_/X _20309_/X _20310_/X _20210_/X VGND VGND VPWR VPWR _20311_/X sky130_fd_sc_hd__a22o_1
XFILLER_107_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36065_ _36065_/CLK _36065_/D VGND VGND VPWR VPWR _36065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33277_ _33531_/CLK _33277_/D VGND VGND VPWR VPWR _33277_/Q sky130_fd_sc_hd__dfxtp_1
Xinput60 DW[63] VGND VGND VPWR VPWR input60/X sky130_fd_sc_hd__clkbuf_16
X_21291_ _35175_/Q _35111_/Q _35047_/Q _32167_/Q _21257_/X _21258_/X VGND VGND VPWR
+ VPWR _21291_/X sky130_fd_sc_hd__mux4_1
Xinput71 R2[0] VGND VGND VPWR VPWR input71/X sky130_fd_sc_hd__clkbuf_1
XFILLER_190_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30489_ _30489_/A VGND VGND VPWR VPWR _35485_/D sky130_fd_sc_hd__clkbuf_1
Xinput82 R3[5] VGND VGND VPWR VPWR input82/X sky130_fd_sc_hd__clkbuf_4
X_35016_ _35658_/CLK _35016_/D VGND VGND VPWR VPWR _35016_/Q sky130_fd_sc_hd__dfxtp_1
X_23030_ input41/X VGND VGND VPWR VPWR _23030_/X sky130_fd_sc_hd__buf_2
X_20242_ _20242_/A VGND VGND VPWR VPWR _32458_/D sky130_fd_sc_hd__clkbuf_4
X_32228_ _35721_/CLK _32228_/D VGND VGND VPWR VPWR _32228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32159_ _35609_/CLK _32159_/D VGND VGND VPWR VPWR _32159_/Q sky130_fd_sc_hd__dfxtp_1
X_20173_ _20173_/A _20173_/B _20173_/C _20173_/D VGND VGND VPWR VPWR _20174_/A sky130_fd_sc_hd__or4_2
XFILLER_130_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24981_ _24981_/A VGND VGND VPWR VPWR _32976_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26720_ _33793_/Q _23432_/X _26732_/S VGND VGND VPWR VPWR _26721_/A sky130_fd_sc_hd__mux2_1
XTAP_4418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35918_ _35982_/CLK _35918_/D VGND VGND VPWR VPWR _35918_/Q sky130_fd_sc_hd__dfxtp_1
X_23932_ _23015_/X _32511_/Q _23948_/S VGND VGND VPWR VPWR _23933_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26651_ _33760_/Q _23261_/X _26669_/S VGND VGND VPWR VPWR _26652_/A sky130_fd_sc_hd__mux2_1
X_35849_ _35849_/CLK _35849_/D VGND VGND VPWR VPWR _35849_/Q sky130_fd_sc_hd__dfxtp_1
X_23863_ _23863_/A VGND VGND VPWR VPWR _32478_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25602_ _24886_/X _33266_/Q _25604_/S VGND VGND VPWR VPWR _25603_/A sky130_fd_sc_hd__mux2_1
X_22814_ _34963_/Q _34899_/Q _34835_/Q _34771_/Q _20683_/X _20685_/X VGND VGND VPWR
+ VPWR _22814_/X sky130_fd_sc_hd__mux4_1
X_29370_ input5/X VGND VGND VPWR VPWR _29370_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_244_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26582_ _26582_/A VGND VGND VPWR VPWR _33729_/D sky130_fd_sc_hd__clkbuf_1
X_23794_ _23794_/A VGND VGND VPWR VPWR _32382_/D sky130_fd_sc_hd__clkbuf_1
X_28321_ _28321_/A VGND VGND VPWR VPWR _34489_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_241_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25533_ _25533_/A VGND VGND VPWR VPWR _33233_/D sky130_fd_sc_hd__clkbuf_1
X_22745_ _20581_/X _22743_/X _22744_/X _20591_/X VGND VGND VPWR VPWR _22745_/X sky130_fd_sc_hd__a22o_1
XFILLER_38_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28252_ _28252_/A VGND VGND VPWR VPWR _34456_/D sky130_fd_sc_hd__clkbuf_1
X_22676_ _32655_/Q _32591_/Q _32527_/Q _35983_/Q _22582_/X _22366_/X VGND VGND VPWR
+ VPWR _22676_/X sky130_fd_sc_hd__mux4_1
X_25464_ _25464_/A VGND VGND VPWR VPWR _33200_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_213_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27203_ _33996_/Q _27202_/X _27218_/S VGND VGND VPWR VPWR _27204_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24415_ _24415_/A VGND VGND VPWR VPWR _32736_/D sky130_fd_sc_hd__clkbuf_1
X_21627_ _21453_/X _21623_/X _21626_/X _21456_/X VGND VGND VPWR VPWR _21627_/X sky130_fd_sc_hd__a22o_1
XFILLER_240_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28183_ _27748_/X _34424_/Q _28193_/S VGND VGND VPWR VPWR _28184_/A sky130_fd_sc_hd__mux2_1
X_25395_ _33169_/Q _23484_/X _25395_/S VGND VGND VPWR VPWR _25396_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27134_ input26/X VGND VGND VPWR VPWR _27134_/X sky130_fd_sc_hd__buf_2
XFILLER_194_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24346_ _23018_/X _32704_/Q _24360_/S VGND VGND VPWR VPWR _24347_/A sky130_fd_sc_hd__mux2_1
X_21558_ _33135_/Q _36015_/Q _33007_/Q _32943_/Q _21309_/X _21310_/X VGND VGND VPWR
+ VPWR _21558_/X sky130_fd_sc_hd__mux4_1
XFILLER_20_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20509_ _20505_/X _20508_/X _20157_/A VGND VGND VPWR VPWR _20517_/C sky130_fd_sc_hd__o21ba_1
X_24277_ _24277_/A VGND VGND VPWR VPWR _32671_/D sky130_fd_sc_hd__clkbuf_1
X_27065_ input2/X VGND VGND VPWR VPWR _27065_/X sky130_fd_sc_hd__clkbuf_4
X_21489_ _21453_/X _21487_/X _21488_/X _21456_/X VGND VGND VPWR VPWR _21489_/X sky130_fd_sc_hd__a22o_1
XTAP_7000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23228_ _28786_/A _27232_/B input84/X VGND VGND VPWR VPWR _23229_/A sky130_fd_sc_hd__or3b_1
X_26016_ _24899_/X _33462_/Q _26030_/S VGND VGND VPWR VPWR _26017_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23159_ _22987_/X _32118_/Q _23173_/S VGND VGND VPWR VPWR _23160_/A sky130_fd_sc_hd__mux2_1
XTAP_7055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_778 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27967_ _27828_/X _34322_/Q _27973_/S VGND VGND VPWR VPWR _27968_/A sky130_fd_sc_hd__mux2_1
XTAP_6365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15981_ _17859_/A VGND VGND VPWR VPWR _15981_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_79_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17720_ _34436_/Q _36164_/Q _34308_/Q _34244_/Q _17582_/X _17583_/X VGND VGND VPWR
+ VPWR _17720_/X sky130_fd_sc_hd__mux4_1
XTAP_5642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29706_ _35114_/Q _29391_/X _29724_/S VGND VGND VPWR VPWR _29707_/A sky130_fd_sc_hd__mux2_1
XTAP_6398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26918_ _33887_/Q _23258_/X _26918_/S VGND VGND VPWR VPWR _26919_/A sky130_fd_sc_hd__mux2_1
XTAP_5664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27898_ _27726_/X _34289_/Q _27902_/S VGND VGND VPWR VPWR _27899_/A sky130_fd_sc_hd__mux2_1
XTAP_4941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17651_ _34946_/Q _34882_/Q _34818_/Q _34754_/Q _17513_/X _17514_/X VGND VGND VPWR
+ VPWR _17651_/X sky130_fd_sc_hd__mux4_1
X_29637_ _29637_/A VGND VGND VPWR VPWR _35081_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26849_ _33854_/Q _23420_/X _26867_/S VGND VGND VPWR VPWR _26850_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_1360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16602_ _16500_/X _16600_/X _16601_/X _16503_/X VGND VGND VPWR VPWR _16602_/X sky130_fd_sc_hd__a22o_1
X_17582_ _17935_/A VGND VGND VPWR VPWR _17582_/X sky130_fd_sc_hd__buf_6
X_29568_ _35049_/Q _29388_/X _29568_/S VGND VGND VPWR VPWR _29569_/A sky130_fd_sc_hd__mux2_1
XFILLER_235_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19321_ _34161_/Q _34097_/Q _34033_/Q _33969_/Q _19040_/X _19041_/X VGND VGND VPWR
+ VPWR _19321_/X sky130_fd_sc_hd__mux4_1
XFILLER_244_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28519_ _27646_/X _34583_/Q _28535_/S VGND VGND VPWR VPWR _28520_/A sky130_fd_sc_hd__mux2_1
XFILLER_216_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16533_ _16493_/X _16531_/X _16532_/X _16498_/X VGND VGND VPWR VPWR _16533_/X sky130_fd_sc_hd__a22o_1
XFILLER_216_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29499_ _29499_/A VGND VGND VPWR VPWR _35020_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31530_ _31530_/A VGND VGND VPWR VPWR _35978_/D sky130_fd_sc_hd__clkbuf_1
X_19252_ _19146_/X _19250_/X _19251_/X _19151_/X VGND VGND VPWR VPWR _19252_/X sky130_fd_sc_hd__a22o_1
XFILLER_189_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16464_ _34145_/Q _34081_/Q _34017_/Q _33953_/Q _16387_/X _16388_/X VGND VGND VPWR
+ VPWR _16464_/X sky130_fd_sc_hd__mux4_1
XFILLER_31_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18203_ _35731_/Q _32243_/Q _35603_/Q _35539_/Q _15993_/X _15995_/X VGND VGND VPWR
+ VPWR _18203_/X sky130_fd_sc_hd__mux4_1
XFILLER_182_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19183_ _19183_/A VGND VGND VPWR VPWR _32428_/D sky130_fd_sc_hd__clkbuf_1
X_31461_ _31551_/S VGND VGND VPWR VPWR _31480_/S sky130_fd_sc_hd__buf_4
XPHY_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16395_ _32607_/Q _32543_/Q _32479_/Q _35935_/Q _16217_/X _16354_/X VGND VGND VPWR
+ VPWR _16395_/X sky130_fd_sc_hd__mux4_1
XPHY_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33200_ _36080_/CLK _33200_/D VGND VGND VPWR VPWR _33200_/Q sky130_fd_sc_hd__dfxtp_1
X_18134_ _17912_/X _18132_/X _18133_/X _17915_/X VGND VGND VPWR VPWR _18134_/X sky130_fd_sc_hd__a22o_1
XFILLER_223_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30412_ _35449_/Q _29438_/X _30420_/S VGND VGND VPWR VPWR _30413_/A sky130_fd_sc_hd__mux2_1
X_34180_ _34180_/CLK _34180_/D VGND VGND VPWR VPWR _34180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31392_ _27801_/X _35913_/Q _31408_/S VGND VGND VPWR VPWR _31393_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33131_ _36010_/CLK _33131_/D VGND VGND VPWR VPWR _33131_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18065_ _17864_/X _18063_/X _18064_/X _17869_/X VGND VGND VPWR VPWR _18065_/X sky130_fd_sc_hd__a22o_1
X_30343_ _35416_/Q _29336_/X _30357_/S VGND VGND VPWR VPWR _30344_/A sky130_fd_sc_hd__mux2_1
XFILLER_208_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17016_ _16805_/X _17014_/X _17015_/X _16810_/X VGND VGND VPWR VPWR _17016_/X sky130_fd_sc_hd__a22o_1
XFILLER_67_1322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33062_ _35755_/CLK _33062_/D VGND VGND VPWR VPWR _33062_/Q sky130_fd_sc_hd__dfxtp_1
X_30274_ _30274_/A VGND VGND VPWR VPWR _35383_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32013_ _36202_/CLK _32013_/D VGND VGND VPWR VPWR _32013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18967_ _33639_/Q _33575_/Q _33511_/Q _33447_/Q _18794_/X _18795_/X VGND VGND VPWR
+ VPWR _18967_/X sky130_fd_sc_hd__mux4_1
XFILLER_224_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17918_ _32650_/Q _32586_/Q _32522_/Q _35978_/Q _17629_/X _17766_/X VGND VGND VPWR
+ VPWR _17918_/X sky130_fd_sc_hd__mux4_1
XFILLER_26_1074 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33964_ _35627_/CLK _33964_/D VGND VGND VPWR VPWR _33964_/Q sky130_fd_sc_hd__dfxtp_1
X_18898_ _34149_/Q _34085_/Q _34021_/Q _33957_/Q _18687_/X _18688_/X VGND VGND VPWR
+ VPWR _18898_/X sky130_fd_sc_hd__mux4_1
XFILLER_113_1044 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35703_ _35703_/CLK _35703_/D VGND VGND VPWR VPWR _35703_/Q sky130_fd_sc_hd__dfxtp_1
X_17849_ _35720_/Q _32230_/Q _35592_/Q _35528_/Q _17670_/X _17671_/X VGND VGND VPWR
+ VPWR _17849_/X sky130_fd_sc_hd__mux4_1
X_32915_ _35985_/CLK _32915_/D VGND VGND VPWR VPWR _32915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33895_ _33895_/CLK _33895_/D VGND VGND VPWR VPWR _33895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20860_ _35675_/Q _32181_/Q _35547_/Q _35483_/Q _20858_/X _20859_/X VGND VGND VPWR
+ VPWR _20860_/X sky130_fd_sc_hd__mux4_1
X_32846_ _32911_/CLK _32846_/D VGND VGND VPWR VPWR _32846_/Q sky130_fd_sc_hd__dfxtp_1
X_35634_ _35634_/CLK _35634_/D VGND VGND VPWR VPWR _35634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19519_ _35702_/Q _32211_/Q _35574_/Q _35510_/Q _19264_/X _19265_/X VGND VGND VPWR
+ VPWR _19519_/X sky130_fd_sc_hd__mux4_1
X_20791_ _20787_/X _20790_/X _20644_/X _20646_/X VGND VGND VPWR VPWR _20808_/B sky130_fd_sc_hd__o211a_1
X_32777_ _32907_/CLK _32777_/D VGND VGND VPWR VPWR _32777_/Q sky130_fd_sc_hd__dfxtp_1
X_35565_ _35693_/CLK _35565_/D VGND VGND VPWR VPWR _35565_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_250_CLK clkbuf_6_63__f_CLK/X VGND VGND VPWR VPWR _34945_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_39_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22530_ _22309_/X _22528_/X _22529_/X _22312_/X VGND VGND VPWR VPWR _22530_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_1186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34516_ _36117_/CLK _34516_/D VGND VGND VPWR VPWR _34516_/Q sky130_fd_sc_hd__dfxtp_1
X_31728_ _31728_/A VGND VGND VPWR VPWR _36072_/D sky130_fd_sc_hd__clkbuf_1
X_35496_ _35687_/CLK _35496_/D VGND VGND VPWR VPWR _35496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22461_ _35208_/Q _35144_/Q _35080_/Q _32264_/Q _22316_/X _22317_/X VGND VGND VPWR
+ VPWR _22461_/X sky130_fd_sc_hd__mux4_1
X_34447_ _36175_/CLK _34447_/D VGND VGND VPWR VPWR _34447_/Q sky130_fd_sc_hd__dfxtp_1
X_31659_ _31686_/S VGND VGND VPWR VPWR _31678_/S sky130_fd_sc_hd__buf_4
XFILLER_33_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21412_ _22471_/A VGND VGND VPWR VPWR _21412_/X sky130_fd_sc_hd__buf_2
X_24200_ _24200_/A VGND VGND VPWR VPWR _32636_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_176_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25180_ _33067_/Q _23296_/X _25196_/S VGND VGND VPWR VPWR _25181_/A sky130_fd_sc_hd__mux2_1
X_22392_ _34438_/Q _36166_/Q _34310_/Q _34246_/Q _22182_/X _22183_/X VGND VGND VPWR
+ VPWR _22392_/X sky130_fd_sc_hd__mux4_1
X_34378_ _35210_/CLK _34378_/D VGND VGND VPWR VPWR _34378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24131_ _24131_/A VGND VGND VPWR VPWR _32603_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36117_ _36117_/CLK _36117_/D VGND VGND VPWR VPWR _36117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21343_ _21093_/X _21339_/X _21342_/X _21098_/X VGND VGND VPWR VPWR _21343_/X sky130_fd_sc_hd__a22o_1
X_33329_ _33393_/CLK _33329_/D VGND VGND VPWR VPWR _33329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24062_ _24062_/A VGND VGND VPWR VPWR _32572_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36048_ _36049_/CLK _36048_/D VGND VGND VPWR VPWR _36048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21274_ _21100_/X _21270_/X _21273_/X _21103_/X VGND VGND VPWR VPWR _21274_/X sky130_fd_sc_hd__a22o_1
XFILLER_2_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23013_ _23011_/X _32062_/Q _23040_/S VGND VGND VPWR VPWR _23014_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20225_ _35722_/Q _32233_/Q _35594_/Q _35530_/Q _19970_/X _19971_/X VGND VGND VPWR
+ VPWR _20225_/X sky130_fd_sc_hd__mux4_1
XFILLER_172_1414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28870_ _28870_/A VGND VGND VPWR VPWR _34748_/D sky130_fd_sc_hd__clkbuf_1
X_27821_ _27821_/A VGND VGND VPWR VPWR _34255_/D sky130_fd_sc_hd__clkbuf_1
X_20156_ _20009_/X _20154_/X _20155_/X _20012_/X VGND VGND VPWR VPWR _20156_/X sky130_fd_sc_hd__a22o_1
XFILLER_89_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27752_ _27751_/X _34233_/Q _27764_/S VGND VGND VPWR VPWR _27753_/A sky130_fd_sc_hd__mux2_1
X_24964_ input49/X VGND VGND VPWR VPWR _24964_/X sky130_fd_sc_hd__buf_4
X_20087_ _20009_/X _20083_/X _20086_/X _20012_/X VGND VGND VPWR VPWR _20087_/X sky130_fd_sc_hd__a22o_1
XFILLER_40_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26703_ _33785_/Q _23405_/X _26711_/S VGND VGND VPWR VPWR _26704_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23915_ _22990_/X _32503_/Q _23927_/S VGND VGND VPWR VPWR _23916_/A sky130_fd_sc_hd__mux2_1
XFILLER_218_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27683_ input5/X VGND VGND VPWR VPWR _27683_/X sky130_fd_sc_hd__buf_4
XFILLER_217_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24895_ _24895_/A VGND VGND VPWR VPWR _32948_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29422_ input24/X VGND VGND VPWR VPWR _29422_/X sky130_fd_sc_hd__buf_2
XFILLER_246_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26634_ _33752_/Q _23237_/X _26648_/S VGND VGND VPWR VPWR _26635_/A sky130_fd_sc_hd__mux2_1
XTAP_3558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23846_ _22879_/X _32470_/Q _23864_/S VGND VGND VPWR VPWR _23847_/A sky130_fd_sc_hd__mux2_1
XTAP_3569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29353_ _29353_/A VGND VGND VPWR VPWR _34973_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26565_ _26565_/A VGND VGND VPWR VPWR _33721_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20989_ _34143_/Q _34079_/Q _34015_/Q _33951_/Q _20987_/X _20988_/X VGND VGND VPWR
+ VPWR _20989_/X sky130_fd_sc_hd__mux4_1
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23777_ _23777_/A VGND VGND VPWR VPWR _32374_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_241_CLK clkbuf_6_60__f_CLK/X VGND VGND VPWR VPWR _36163_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_53_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28304_ _28304_/A VGND VGND VPWR VPWR _34481_/D sky130_fd_sc_hd__clkbuf_1
X_25516_ _24958_/X _33225_/Q _25532_/S VGND VGND VPWR VPWR _25517_/A sky130_fd_sc_hd__mux2_1
X_22728_ _22728_/A VGND VGND VPWR VPWR _36240_/D sky130_fd_sc_hd__clkbuf_1
X_29284_ _29284_/A VGND VGND VPWR VPWR _34944_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_213_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26496_ _26496_/A VGND VGND VPWR VPWR _33688_/D sky130_fd_sc_hd__clkbuf_1
X_28235_ _27825_/X _34449_/Q _28235_/S VGND VGND VPWR VPWR _28236_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25447_ _25447_/A VGND VGND VPWR VPWR _33192_/D sky130_fd_sc_hd__clkbuf_1
X_22659_ _22655_/X _22658_/X _22457_/X VGND VGND VPWR VPWR _22667_/C sky130_fd_sc_hd__o21ba_1
XFILLER_51_1134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16180_ _16140_/X _16178_/X _16179_/X _16145_/X VGND VGND VPWR VPWR _16180_/X sky130_fd_sc_hd__a22o_1
XFILLER_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28166_ _27723_/X _34416_/Q _28172_/S VGND VGND VPWR VPWR _28167_/A sky130_fd_sc_hd__mux2_1
X_25378_ _25378_/A VGND VGND VPWR VPWR _33160_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27117_ _27117_/A VGND VGND VPWR VPWR _33968_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24329_ _22993_/X _32696_/Q _24339_/S VGND VGND VPWR VPWR _24330_/A sky130_fd_sc_hd__mux2_1
X_28097_ _28097_/A VGND VGND VPWR VPWR _34383_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27048_ _33946_/Q _27047_/X _27063_/S VGND VGND VPWR VPWR _27049_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19870_ _19720_/X _19868_/X _19869_/X _19724_/X VGND VGND VPWR VPWR _19870_/X sky130_fd_sc_hd__a22o_1
XFILLER_122_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18821_ _35170_/Q _35106_/Q _35042_/Q _32162_/Q _18604_/X _18605_/X VGND VGND VPWR
+ VPWR _18821_/X sky130_fd_sc_hd__mux4_1
XTAP_6140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1066 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28999_ _28999_/A VGND VGND VPWR VPWR _34809_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18752_ _19458_/A VGND VGND VPWR VPWR _18752_/X sky130_fd_sc_hd__clkbuf_4
XTAP_5450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17703_ _17697_/X _17702_/X _17493_/X _17494_/X VGND VGND VPWR VPWR _17724_/B sky130_fd_sc_hd__o211a_1
XFILLER_114_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18683_ _18679_/X _18682_/X _18404_/X VGND VGND VPWR VPWR _18684_/D sky130_fd_sc_hd__o21ba_2
XTAP_5494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30961_ _30961_/A VGND VGND VPWR VPWR _35709_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32700_ _32895_/CLK _32700_/D VGND VGND VPWR VPWR _32700_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_480_CLK clkbuf_6_10__f_CLK/X VGND VGND VPWR VPWR _35627_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_76_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17634_ _32130_/Q _32322_/Q _32386_/Q _35906_/Q _17633_/X _17421_/X VGND VGND VPWR
+ VPWR _17634_/X sky130_fd_sc_hd__mux4_1
XFILLER_84_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33680_ _34064_/CLK _33680_/D VGND VGND VPWR VPWR _33680_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30892_ _30892_/A VGND VGND VPWR VPWR _35676_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32631_ _34485_/CLK _32631_/D VGND VGND VPWR VPWR _32631_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17565_ _32640_/Q _32576_/Q _32512_/Q _35968_/Q _17276_/X _17413_/X VGND VGND VPWR
+ VPWR _17565_/X sky130_fd_sc_hd__mux4_1
XFILLER_189_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_232_CLK clkbuf_6_55__f_CLK/X VGND VGND VPWR VPWR _36109_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_182_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19304_ _35440_/Q _35376_/Q _35312_/Q _35248_/Q _19201_/X _19202_/X VGND VGND VPWR
+ VPWR _19304_/X sky130_fd_sc_hd__mux4_1
X_35350_ _36118_/CLK _35350_/D VGND VGND VPWR VPWR _35350_/Q sky130_fd_sc_hd__dfxtp_1
X_16516_ _35426_/Q _35362_/Q _35298_/Q _35234_/Q _16195_/X _16196_/X VGND VGND VPWR
+ VPWR _16516_/X sky130_fd_sc_hd__mux4_1
X_32562_ _32882_/CLK _32562_/D VGND VGND VPWR VPWR _32562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17496_ _35710_/Q _32219_/Q _35582_/Q _35518_/Q _17317_/X _17318_/X VGND VGND VPWR
+ VPWR _17496_/X sky130_fd_sc_hd__mux4_1
XFILLER_17_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_833 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31513_ _31513_/A VGND VGND VPWR VPWR _35970_/D sky130_fd_sc_hd__clkbuf_1
X_19235_ _35438_/Q _35374_/Q _35310_/Q _35246_/Q _19201_/X _19202_/X VGND VGND VPWR
+ VPWR _19235_/X sky130_fd_sc_hd__mux4_1
X_34301_ _36154_/CLK _34301_/D VGND VGND VPWR VPWR _34301_/Q sky130_fd_sc_hd__dfxtp_1
X_35281_ _35859_/CLK _35281_/D VGND VGND VPWR VPWR _35281_/Q sky130_fd_sc_hd__dfxtp_1
X_16447_ _17153_/A VGND VGND VPWR VPWR _16447_/X sky130_fd_sc_hd__buf_4
XFILLER_182_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32493_ _35883_/CLK _32493_/D VGND VGND VPWR VPWR _32493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_899 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34232_ _35192_/CLK _34232_/D VGND VGND VPWR VPWR _34232_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31444_ _31444_/A VGND VGND VPWR VPWR _35937_/D sky130_fd_sc_hd__clkbuf_1
X_19166_ _35692_/Q _32200_/Q _35564_/Q _35500_/Q _18911_/X _18912_/X VGND VGND VPWR
+ VPWR _19166_/X sky130_fd_sc_hd__mux4_1
X_16378_ _35166_/Q _35102_/Q _35038_/Q _32158_/Q _16304_/X _16305_/X VGND VGND VPWR
+ VPWR _16378_/X sky130_fd_sc_hd__mux4_1
XFILLER_160_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18117_ _33104_/Q _32080_/Q _35856_/Q _35792_/Q _16079_/X _16080_/X VGND VGND VPWR
+ VPWR _18117_/X sky130_fd_sc_hd__mux4_1
X_34163_ _35697_/CLK _34163_/D VGND VGND VPWR VPWR _34163_/Q sky130_fd_sc_hd__dfxtp_1
X_31375_ _27776_/X _35905_/Q _31387_/S VGND VGND VPWR VPWR _31376_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19097_ _18950_/X _19095_/X _19096_/X _18953_/X VGND VGND VPWR VPWR _19097_/X sky130_fd_sc_hd__a22o_1
XFILLER_69_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33114_ _34007_/CLK _33114_/D VGND VGND VPWR VPWR _33114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_219_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30326_ _30326_/A VGND VGND VPWR VPWR _35408_/D sky130_fd_sc_hd__clkbuf_1
X_18048_ _17765_/X _18046_/X _18047_/X _17771_/X VGND VGND VPWR VPWR _18048_/X sky130_fd_sc_hd__a22o_1
XFILLER_105_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34094_ _35630_/CLK _34094_/D VGND VGND VPWR VPWR _34094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_299_CLK clkbuf_6_57__f_CLK/X VGND VGND VPWR VPWR _35651_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_99_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33045_ _36053_/CLK _33045_/D VGND VGND VPWR VPWR _33045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_236_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30257_ _30257_/A VGND VGND VPWR VPWR _35375_/D sky130_fd_sc_hd__clkbuf_1
X_20010_ _35460_/Q _35396_/Q _35332_/Q _35268_/Q _19907_/X _19908_/X VGND VGND VPWR
+ VPWR _20010_/X sky130_fd_sc_hd__mux4_1
XFILLER_8_1219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30188_ _35343_/Q _29506_/X _30192_/S VGND VGND VPWR VPWR _30189_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19999_ _20133_/A VGND VGND VPWR VPWR _19999_/X sky130_fd_sc_hd__buf_4
XFILLER_41_1303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34996_ _35446_/CLK _34996_/D VGND VGND VPWR VPWR _34996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33947_ _36212_/CLK _33947_/D VGND VGND VPWR VPWR _33947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21961_ _21955_/X _21960_/X _21751_/X VGND VGND VPWR VPWR _21971_/C sky130_fd_sc_hd__o21ba_1
XFILLER_95_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23700_ _23079_/X _32340_/Q _23702_/S VGND VGND VPWR VPWR _23701_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_471_CLK clkbuf_6_11__f_CLK/X VGND VGND VPWR VPWR _35566_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20912_ _20912_/A _20912_/B _20912_/C _20912_/D VGND VGND VPWR VPWR _20913_/A sky130_fd_sc_hd__or4_1
X_24680_ _24680_/A VGND VGND VPWR VPWR _32862_/D sky130_fd_sc_hd__clkbuf_1
X_21892_ _22598_/A VGND VGND VPWR VPWR _21892_/X sky130_fd_sc_hd__buf_8
X_33878_ _36055_/CLK _33878_/D VGND VGND VPWR VPWR _33878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20843_ _20843_/A VGND VGND VPWR VPWR _36186_/D sky130_fd_sc_hd__clkbuf_2
X_35617_ _35620_/CLK _35617_/D VGND VGND VPWR VPWR _35617_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23631_ _22977_/X _32307_/Q _23631_/S VGND VGND VPWR VPWR _23632_/A sky130_fd_sc_hd__mux2_1
X_32829_ _32891_/CLK _32829_/D VGND VGND VPWR VPWR _32829_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_223_CLK clkbuf_6_53__f_CLK/X VGND VGND VPWR VPWR _34954_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_74_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_1254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26350_ _24994_/X _33621_/Q _26350_/S VGND VGND VPWR VPWR _26351_/A sky130_fd_sc_hd__mux2_1
X_20774_ _20691_/X _20772_/X _20773_/X _20701_/X VGND VGND VPWR VPWR _20774_/X sky130_fd_sc_hd__a22o_1
X_23562_ _23562_/A VGND VGND VPWR VPWR _32275_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35548_ _36058_/CLK _35548_/D VGND VGND VPWR VPWR _35548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25301_ _33124_/Q _23274_/X _25311_/S VGND VGND VPWR VPWR _25302_/A sky130_fd_sc_hd__mux2_1
X_22513_ _33418_/Q _33354_/Q _33290_/Q _33226_/Q _22433_/X _22434_/X VGND VGND VPWR
+ VPWR _22513_/X sky130_fd_sc_hd__mux4_1
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23493_ _32243_/Q _23492_/X _23499_/S VGND VGND VPWR VPWR _23494_/A sky130_fd_sc_hd__mux2_1
X_26281_ _26350_/S VGND VGND VPWR VPWR _26300_/S sky130_fd_sc_hd__buf_4
XFILLER_50_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35479_ _35735_/CLK _35479_/D VGND VGND VPWR VPWR _35479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28020_ _28020_/A VGND VGND VPWR VPWR _34346_/D sky130_fd_sc_hd__clkbuf_1
X_25232_ _33092_/Q _23441_/X _25238_/S VGND VGND VPWR VPWR _25233_/A sky130_fd_sc_hd__mux2_1
X_22444_ _32904_/Q _32840_/Q _32776_/Q _32712_/Q _22299_/X _22300_/X VGND VGND VPWR
+ VPWR _22444_/X sky130_fd_sc_hd__mux4_1
XFILLER_109_804 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22375_ _32134_/Q _32326_/Q _32390_/Q _35910_/Q _22233_/X _22374_/X VGND VGND VPWR
+ VPWR _22375_/X sky130_fd_sc_hd__mux4_1
X_25163_ _33059_/Q _23271_/X _25175_/S VGND VGND VPWR VPWR _25164_/A sky130_fd_sc_hd__mux2_1
XFILLER_136_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24114_ _24114_/A VGND VGND VPWR VPWR _32597_/D sky130_fd_sc_hd__clkbuf_1
X_21326_ _22536_/A VGND VGND VPWR VPWR _21326_/X sky130_fd_sc_hd__buf_4
X_25094_ _25094_/A VGND VGND VPWR VPWR _33027_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29971_ _35240_/Q _29385_/X _29973_/S VGND VGND VPWR VPWR _29972_/A sky130_fd_sc_hd__mux2_1
X_28922_ _28922_/A VGND VGND VPWR VPWR _34773_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21257_ _22316_/A VGND VGND VPWR VPWR _21257_/X sky130_fd_sc_hd__buf_6
X_24045_ _22980_/X _32564_/Q _24063_/S VGND VGND VPWR VPWR _24046_/A sky130_fd_sc_hd__mux2_1
XFILLER_176_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20208_ _33674_/Q _33610_/Q _33546_/Q _33482_/Q _20206_/X _20207_/X VGND VGND VPWR
+ VPWR _20208_/X sky130_fd_sc_hd__mux4_1
XFILLER_137_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28853_ _34740_/Q _27127_/X _28871_/S VGND VGND VPWR VPWR _28854_/A sky130_fd_sc_hd__mux2_1
X_21188_ _34660_/Q _34596_/Q _34532_/Q _34468_/Q _21186_/X _21187_/X VGND VGND VPWR
+ VPWR _21188_/X sky130_fd_sc_hd__mux4_1
XFILLER_133_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27804_ input48/X VGND VGND VPWR VPWR _27804_/X sky130_fd_sc_hd__clkbuf_4
X_20139_ _20132_/X _20137_/X _20138_/X VGND VGND VPWR VPWR _20173_/A sky130_fd_sc_hd__o21ba_2
XFILLER_38_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28784_ _34709_/Q _27229_/X _28784_/S VGND VGND VPWR VPWR _28785_/A sky130_fd_sc_hd__mux2_1
XTAP_4001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25996_ _25996_/A VGND VGND VPWR VPWR _33452_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27735_ input24/X VGND VGND VPWR VPWR _27735_/X sky130_fd_sc_hd__buf_2
XFILLER_86_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24947_ _24947_/A VGND VGND VPWR VPWR _32965_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_462_CLK clkbuf_6_9__f_CLK/X VGND VGND VPWR VPWR _35180_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27666_ _27666_/A VGND VGND VPWR VPWR _34205_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24878_ _24877_/X _32943_/Q _24890_/S VGND VGND VPWR VPWR _24879_/A sky130_fd_sc_hd__mux2_1
XTAP_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29405_ _34990_/Q _29404_/X _29420_/S VGND VGND VPWR VPWR _29406_/A sky130_fd_sc_hd__mux2_1
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26617_ _26617_/A VGND VGND VPWR VPWR _33746_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23829_ _23829_/A VGND VGND VPWR VPWR _32399_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27597_ _27597_/A VGND VGND VPWR VPWR _34177_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_214_CLK clkbuf_6_52__f_CLK/X VGND VGND VPWR VPWR _35663_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_26_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29336_ input23/X VGND VGND VPWR VPWR _29336_/X sky130_fd_sc_hd__buf_2
XFILLER_57_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17350_ _17344_/X _17349_/X _17140_/X _17141_/X VGND VGND VPWR VPWR _17371_/B sky130_fd_sc_hd__o211a_1
X_26548_ _26548_/A VGND VGND VPWR VPWR _33713_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_884 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _16297_/X _16298_/X _16299_/X _16300_/X VGND VGND VPWR VPWR _16301_/X sky130_fd_sc_hd__a22o_1
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29267_ _29267_/A VGND VGND VPWR VPWR _34936_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17281_ _32120_/Q _32312_/Q _32376_/Q _35896_/Q _17280_/X _17068_/X VGND VGND VPWR
+ VPWR _17281_/X sky130_fd_sc_hd__mux4_1
X_26479_ _26479_/A VGND VGND VPWR VPWR _33681_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19020_ _19013_/X _19019_/X _18734_/X _18735_/X VGND VGND VPWR VPWR _19037_/B sky130_fd_sc_hd__o211a_2
X_28218_ _28218_/A VGND VGND VPWR VPWR _34440_/D sky130_fd_sc_hd__clkbuf_1
X_16232_ _16228_/X _16231_/X _16075_/X VGND VGND VPWR VPWR _16242_/C sky130_fd_sc_hd__o21ba_1
XFILLER_13_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29198_ _29198_/A VGND VGND VPWR VPWR _34903_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16163_ _35416_/Q _35352_/Q _35288_/Q _35224_/Q _16062_/X _16064_/X VGND VGND VPWR
+ VPWR _16163_/X sky130_fd_sc_hd__mux4_1
X_28149_ _27698_/X _34408_/Q _28151_/S VGND VGND VPWR VPWR _28150_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31160_ _27658_/X _35803_/Q _31168_/S VGND VGND VPWR VPWR _31161_/A sky130_fd_sc_hd__mux2_1
X_16094_ _16877_/A VGND VGND VPWR VPWR _16094_/X sky130_fd_sc_hd__buf_4
XFILLER_55_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30111_ _35306_/Q _29391_/X _30129_/S VGND VGND VPWR VPWR _30112_/A sky130_fd_sc_hd__mux2_1
X_19922_ _33666_/Q _33602_/Q _33538_/Q _33474_/Q _19853_/X _19854_/X VGND VGND VPWR
+ VPWR _19922_/X sky130_fd_sc_hd__mux4_1
XFILLER_138_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31091_ _35771_/Q input31/X _31095_/S VGND VGND VPWR VPWR _31092_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30042_ _30042_/A VGND VGND VPWR VPWR _35273_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19853_ _20206_/A VGND VGND VPWR VPWR _19853_/X sky130_fd_sc_hd__buf_4
XFILLER_116_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18804_ _18800_/X _18801_/X _18802_/X _18803_/X VGND VGND VPWR VPWR _18804_/X sky130_fd_sc_hd__a22o_1
XFILLER_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34850_ _34914_/CLK _34850_/D VGND VGND VPWR VPWR _34850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19784_ _19506_/X _19782_/X _19783_/X _19509_/X VGND VGND VPWR VPWR _19784_/X sky130_fd_sc_hd__a22o_1
X_16996_ _16714_/X _16992_/X _16995_/X _16718_/X VGND VGND VPWR VPWR _16996_/X sky130_fd_sc_hd__a22o_1
XFILLER_209_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33801_ _36105_/CLK _33801_/D VGND VGND VPWR VPWR _33801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18735_ _20147_/A VGND VGND VPWR VPWR _18735_/X sky130_fd_sc_hd__buf_2
X_34781_ _36242_/CLK _34781_/D VGND VGND VPWR VPWR _34781_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31993_ _34405_/CLK _31993_/D VGND VGND VPWR VPWR _31993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_453_CLK clkbuf_6_14__f_CLK/X VGND VGND VPWR VPWR _34413_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_76_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33732_ _35525_/CLK _33732_/D VGND VGND VPWR VPWR _33732_/Q sky130_fd_sc_hd__dfxtp_1
X_18666_ _18661_/X _18663_/X _18664_/X _18665_/X VGND VGND VPWR VPWR _18666_/X sky130_fd_sc_hd__a22o_1
X_30944_ _35701_/Q input25/X _30960_/S VGND VGND VPWR VPWR _30945_/A sky130_fd_sc_hd__mux2_1
XTAP_4590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17617_ _34945_/Q _34881_/Q _34817_/Q _34753_/Q _17513_/X _17514_/X VGND VGND VPWR
+ VPWR _17617_/X sky130_fd_sc_hd__mux4_1
XFILLER_51_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30875_ _35669_/Q input60/X _30875_/S VGND VGND VPWR VPWR _30876_/A sky130_fd_sc_hd__mux2_1
X_33663_ _35456_/CLK _33663_/D VGND VGND VPWR VPWR _33663_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18597_ _20164_/A VGND VGND VPWR VPWR _18597_/X sky130_fd_sc_hd__buf_4
XFILLER_149_1268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_205_CLK clkbuf_6_54__f_CLK/X VGND VGND VPWR VPWR _35718_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_75_1432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35402_ _35723_/CLK _35402_/D VGND VGND VPWR VPWR _35402_/Q sky130_fd_sc_hd__dfxtp_1
X_17548_ _17511_/X _17546_/X _17547_/X _17516_/X VGND VGND VPWR VPWR _17548_/X sky130_fd_sc_hd__a22o_1
XFILLER_205_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32614_ _35945_/CLK _32614_/D VGND VGND VPWR VPWR _32614_/Q sky130_fd_sc_hd__dfxtp_1
X_33594_ _33913_/CLK _33594_/D VGND VGND VPWR VPWR _33594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35333_ _35463_/CLK _35333_/D VGND VGND VPWR VPWR _35333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32545_ _35875_/CLK _32545_/D VGND VGND VPWR VPWR _32545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17479_ _17199_/X _17477_/X _17478_/X _17204_/X VGND VGND VPWR VPWR _17479_/X sky130_fd_sc_hd__a22o_1
XFILLER_221_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19218_ _19146_/X _19216_/X _19217_/X _19151_/X VGND VGND VPWR VPWR _19218_/X sky130_fd_sc_hd__a22o_1
X_20490_ _34195_/Q _34131_/Q _34067_/Q _34003_/Q _18349_/X _18350_/X VGND VGND VPWR
+ VPWR _20490_/X sky130_fd_sc_hd__mux4_1
X_32476_ _35998_/CLK _32476_/D VGND VGND VPWR VPWR _32476_/Q sky130_fd_sc_hd__dfxtp_1
X_35264_ _35839_/CLK _35264_/D VGND VGND VPWR VPWR _35264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31427_ _31427_/A VGND VGND VPWR VPWR _35929_/D sky130_fd_sc_hd__clkbuf_1
X_19149_ _33644_/Q _33580_/Q _33516_/Q _33452_/Q _19147_/X _19148_/X VGND VGND VPWR
+ VPWR _19149_/X sky130_fd_sc_hd__mux4_1
X_34215_ _35554_/CLK _34215_/D VGND VGND VPWR VPWR _34215_/Q sky130_fd_sc_hd__dfxtp_1
X_35195_ _35644_/CLK _35195_/D VGND VGND VPWR VPWR _35195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22160_ _33408_/Q _33344_/Q _33280_/Q _33216_/Q _22080_/X _22081_/X VGND VGND VPWR
+ VPWR _22160_/X sky130_fd_sc_hd__mux4_1
X_34146_ _34146_/CLK _34146_/D VGND VGND VPWR VPWR _34146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_1471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31358_ _27751_/X _35897_/Q _31366_/S VGND VGND VPWR VPWR _31359_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21111_ _20961_/X _21109_/X _21110_/X _20965_/X VGND VGND VPWR VPWR _21111_/X sky130_fd_sc_hd__a22o_1
XFILLER_12_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30309_ _35400_/Q _29484_/X _30327_/S VGND VGND VPWR VPWR _30310_/A sky130_fd_sc_hd__mux2_1
X_34077_ _36188_/CLK _34077_/D VGND VGND VPWR VPWR _34077_/Q sky130_fd_sc_hd__dfxtp_1
X_22091_ _32894_/Q _32830_/Q _32766_/Q _32702_/Q _21946_/X _21947_/X VGND VGND VPWR
+ VPWR _22091_/X sky130_fd_sc_hd__mux4_1
XTAP_6909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31289_ _27649_/X _35864_/Q _31303_/S VGND VGND VPWR VPWR _31290_/A sky130_fd_sc_hd__mux2_1
X_33028_ _36038_/CLK _33028_/D VGND VGND VPWR VPWR _33028_/Q sky130_fd_sc_hd__dfxtp_1
X_21042_ _35424_/Q _35360_/Q _35296_/Q _35232_/Q _20795_/X _20796_/X VGND VGND VPWR
+ VPWR _21042_/X sky130_fd_sc_hd__mux4_1
XFILLER_141_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25850_ _25850_/A VGND VGND VPWR VPWR _33383_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24801_ _24796_/X _32918_/Q _24828_/S VGND VGND VPWR VPWR _24802_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25781_ _24951_/X _33351_/Q _25781_/S VGND VGND VPWR VPWR _25782_/A sky130_fd_sc_hd__mux2_1
X_22993_ input28/X VGND VGND VPWR VPWR _22993_/X sky130_fd_sc_hd__clkbuf_4
X_34979_ _35176_/CLK _34979_/D VGND VGND VPWR VPWR _34979_/Q sky130_fd_sc_hd__dfxtp_1
X_27520_ _34141_/Q _27056_/X _27524_/S VGND VGND VPWR VPWR _27521_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_444_CLK clkbuf_leaf_61_CLK/A VGND VGND VPWR VPWR _32911_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_41_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24732_ _22990_/X _32887_/Q _24744_/S VGND VGND VPWR VPWR _24733_/A sky130_fd_sc_hd__mux2_1
X_21944_ _21659_/X _21942_/X _21943_/X _21665_/X VGND VGND VPWR VPWR _21944_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27451_ _27451_/A VGND VGND VPWR VPWR _34108_/D sky130_fd_sc_hd__clkbuf_1
X_24663_ _22879_/X _32854_/Q _24681_/S VGND VGND VPWR VPWR _24664_/A sky130_fd_sc_hd__mux2_1
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_24__f_CLK clkbuf_5_12_0_CLK/X VGND VGND VPWR VPWR clkbuf_leaf_73_CLK/A sky130_fd_sc_hd__clkbuf_16
XFILLER_27_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21875_ _21871_/X _21874_/X _21732_/X VGND VGND VPWR VPWR _21901_/A sky130_fd_sc_hd__o21ba_1
XFILLER_54_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_890 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26402_ _26402_/A VGND VGND VPWR VPWR _33644_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23614_ _23614_/A VGND VGND VPWR VPWR _32298_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_247_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20826_ _35674_/Q _32180_/Q _35546_/Q _35482_/Q _20649_/X _20650_/X VGND VGND VPWR
+ VPWR _20826_/X sky130_fd_sc_hd__mux4_1
X_27382_ _27382_/A VGND VGND VPWR VPWR _34075_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24594_ _24594_/A VGND VGND VPWR VPWR _32821_/D sky130_fd_sc_hd__clkbuf_1
X_29121_ _29121_/A VGND VGND VPWR VPWR _34867_/D sky130_fd_sc_hd__clkbuf_1
X_26333_ _26333_/A VGND VGND VPWR VPWR _33612_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23545_ _32267_/Q _23466_/X _23557_/S VGND VGND VPWR VPWR _23546_/A sky130_fd_sc_hd__mux2_1
X_20757_ _32856_/Q _32792_/Q _32728_/Q _32664_/Q _20637_/X _20639_/X VGND VGND VPWR
+ VPWR _20757_/X sky130_fd_sc_hd__mux4_1
XFILLER_10_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29052_ _34835_/Q _27223_/X _29056_/S VGND VGND VPWR VPWR _29053_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26264_ _26264_/A VGND VGND VPWR VPWR _33579_/D sky130_fd_sc_hd__clkbuf_1
X_20688_ _21756_/A VGND VGND VPWR VPWR _20688_/X sky130_fd_sc_hd__buf_4
XFILLER_195_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23476_ _32237_/Q _23475_/X _23485_/S VGND VGND VPWR VPWR _23477_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28003_ _28003_/A VGND VGND VPWR VPWR _34338_/D sky130_fd_sc_hd__clkbuf_1
X_25215_ _33084_/Q _23414_/X _25217_/S VGND VGND VPWR VPWR _25216_/A sky130_fd_sc_hd__mux2_1
X_22427_ _22423_/X _22426_/X _22118_/X VGND VGND VPWR VPWR _22428_/D sky130_fd_sc_hd__o21ba_1
X_26195_ _24964_/X _33547_/Q _26207_/S VGND VGND VPWR VPWR _26196_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25146_ _33051_/Q _23246_/X _25154_/S VGND VGND VPWR VPWR _25147_/A sky130_fd_sc_hd__mux2_1
X_22358_ _33670_/Q _33606_/Q _33542_/Q _33478_/Q _22153_/X _22154_/X VGND VGND VPWR
+ VPWR _22358_/X sky130_fd_sc_hd__mux4_1
XFILLER_174_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21309_ _22506_/A VGND VGND VPWR VPWR _21309_/X sky130_fd_sc_hd__buf_4
X_22289_ _34180_/Q _34116_/Q _34052_/Q _33988_/Q _22046_/X _22047_/X VGND VGND VPWR
+ VPWR _22289_/X sky130_fd_sc_hd__mux4_1
X_29954_ _30065_/S VGND VGND VPWR VPWR _29973_/S sky130_fd_sc_hd__buf_4
X_25077_ _25077_/A VGND VGND VPWR VPWR _33019_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28905_ _34765_/Q _27205_/X _28913_/S VGND VGND VPWR VPWR _28906_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24028_ _22956_/X _32556_/Q _24042_/S VGND VGND VPWR VPWR _24029_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29885_ _35199_/Q _29457_/X _29901_/S VGND VGND VPWR VPWR _29886_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16850_ _34156_/Q _34092_/Q _34028_/Q _33964_/Q _16740_/X _16741_/X VGND VGND VPWR
+ VPWR _16850_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28836_ _34732_/Q _27103_/X _28850_/S VGND VGND VPWR VPWR _28837_/A sky130_fd_sc_hd__mux2_1
XFILLER_219_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28767_ _28767_/A VGND VGND VPWR VPWR _34700_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16781_ _32618_/Q _32554_/Q _32490_/Q _35946_/Q _16570_/X _16707_/X VGND VGND VPWR
+ VPWR _16781_/X sky130_fd_sc_hd__mux4_1
X_25979_ _25979_/A VGND VGND VPWR VPWR _33444_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18520_ _18318_/X _18518_/X _18519_/X _18327_/X VGND VGND VPWR VPWR _18520_/X sky130_fd_sc_hd__a22o_1
XFILLER_20_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_435_CLK clkbuf_6_36__f_CLK/X VGND VGND VPWR VPWR _34611_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_219_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27718_ _27717_/X _34222_/Q _27733_/S VGND VGND VPWR VPWR _27719_/A sky130_fd_sc_hd__mux2_1
XTAP_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28698_ _28698_/A VGND VGND VPWR VPWR _34667_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18451_ _18447_/X _18448_/X _18449_/X _18450_/X VGND VGND VPWR VPWR _18451_/X sky130_fd_sc_hd__a22o_1
XTAP_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27649_ input23/X VGND VGND VPWR VPWR _27649_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_18_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17402_ _17398_/X _17401_/X _17165_/X VGND VGND VPWR VPWR _17403_/D sky130_fd_sc_hd__o21ba_1
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18382_ _20282_/A VGND VGND VPWR VPWR _20016_/A sky130_fd_sc_hd__buf_12
X_30660_ _30660_/A VGND VGND VPWR VPWR _35566_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29319_ _29319_/A VGND VGND VPWR VPWR _34961_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17333_ _17333_/A _17333_/B _17333_/C _17333_/D VGND VGND VPWR VPWR _17334_/A sky130_fd_sc_hd__or4_4
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30591_ _35534_/Q _29503_/X _30597_/S VGND VGND VPWR VPWR _30592_/A sky130_fd_sc_hd__mux2_1
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32330_ _32907_/CLK _32330_/D VGND VGND VPWR VPWR _32330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17264_ _34935_/Q _34871_/Q _34807_/Q _34743_/Q _17160_/X _17161_/X VGND VGND VPWR
+ VPWR _17264_/X sky130_fd_sc_hd__mux4_1
XFILLER_105_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19003_ _33896_/Q _33832_/Q _33768_/Q _36072_/Q _18971_/X _18972_/X VGND VGND VPWR
+ VPWR _19003_/X sky130_fd_sc_hd__mux4_1
X_16215_ _16147_/X _16213_/X _16214_/X _16150_/X VGND VGND VPWR VPWR _16215_/X sky130_fd_sc_hd__a22o_1
XFILLER_70_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32261_ _35718_/CLK _32261_/D VGND VGND VPWR VPWR _32261_/Q sky130_fd_sc_hd__dfxtp_1
X_17195_ _17158_/X _17193_/X _17194_/X _17163_/X VGND VGND VPWR VPWR _17195_/X sky130_fd_sc_hd__a22o_1
X_34000_ _34192_/CLK _34000_/D VGND VGND VPWR VPWR _34000_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31212_ _31281_/S VGND VGND VPWR VPWR _31231_/S sky130_fd_sc_hd__buf_6
X_16146_ _16140_/X _16143_/X _16144_/X _16145_/X VGND VGND VPWR VPWR _16146_/X sky130_fd_sc_hd__a22o_1
XFILLER_128_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32192_ _35559_/CLK _32192_/D VGND VGND VPWR VPWR _32192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31143_ _35796_/Q input59/X _31145_/S VGND VGND VPWR VPWR _31144_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16077_ _17765_/A VGND VGND VPWR VPWR _17153_/A sky130_fd_sc_hd__buf_8
X_19905_ _35649_/Q _35009_/Q _34369_/Q _33729_/Q _19797_/X _19798_/X VGND VGND VPWR
+ VPWR _19905_/X sky130_fd_sc_hd__mux4_1
XFILLER_130_618 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31074_ _35763_/Q input22/X _31074_/S VGND VGND VPWR VPWR _31075_/A sky130_fd_sc_hd__mux2_1
X_35951_ _35951_/CLK _35951_/D VGND VGND VPWR VPWR _35951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_216_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34902_ _34903_/CLK _34902_/D VGND VGND VPWR VPWR _34902_/Q sky130_fd_sc_hd__dfxtp_1
X_30025_ _30025_/A VGND VGND VPWR VPWR _35265_/D sky130_fd_sc_hd__clkbuf_1
X_19836_ _35711_/Q _32221_/Q _35583_/Q _35519_/Q _19617_/X _19618_/X VGND VGND VPWR
+ VPWR _19836_/X sky130_fd_sc_hd__mux4_1
XFILLER_9_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35882_ _35883_/CLK _35882_/D VGND VGND VPWR VPWR _35882_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34833_ _34897_/CLK _34833_/D VGND VGND VPWR VPWR _34833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19767_ _19763_/X _19766_/X _19451_/X VGND VGND VPWR VPWR _19775_/C sky130_fd_sc_hd__o21ba_1
Xinput3 DW[11] VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__buf_6
X_16979_ _16975_/X _16978_/X _16812_/X VGND VGND VPWR VPWR _16980_/D sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_426_CLK clkbuf_6_35__f_CLK/X VGND VGND VPWR VPWR _35124_/CLK sky130_fd_sc_hd__clkbuf_16
X_18718_ _33632_/Q _33568_/Q _33504_/Q _33440_/Q _18441_/X _18442_/X VGND VGND VPWR
+ VPWR _18718_/X sky130_fd_sc_hd__mux4_1
X_34764_ _34957_/CLK _34764_/D VGND VGND VPWR VPWR _34764_/Q sky130_fd_sc_hd__dfxtp_1
X_31976_ _34790_/CLK _31976_/D VGND VGND VPWR VPWR _31976_/Q sky130_fd_sc_hd__dfxtp_1
X_19698_ _19453_/X _19696_/X _19697_/X _19456_/X VGND VGND VPWR VPWR _19698_/X sky130_fd_sc_hd__a22o_1
XFILLER_225_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33715_ _35635_/CLK _33715_/D VGND VGND VPWR VPWR _33715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18649_ _33374_/Q _33310_/Q _33246_/Q _33182_/Q _18302_/X _18303_/X VGND VGND VPWR
+ VPWR _18649_/X sky130_fd_sc_hd__mux4_1
X_30927_ _35693_/Q input16/X _30939_/S VGND VGND VPWR VPWR _30928_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34695_ _35657_/CLK _34695_/D VGND VGND VPWR VPWR _34695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_939 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30858_ _30858_/A VGND VGND VPWR VPWR _35660_/D sky130_fd_sc_hd__clkbuf_1
X_33646_ _33902_/CLK _33646_/D VGND VGND VPWR VPWR _33646_/Q sky130_fd_sc_hd__dfxtp_1
X_21660_ _22366_/A VGND VGND VPWR VPWR _21660_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_178_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20611_ _22561_/A VGND VGND VPWR VPWR _20611_/X sky130_fd_sc_hd__buf_4
X_21591_ _21306_/X _21589_/X _21590_/X _21312_/X VGND VGND VPWR VPWR _21591_/X sky130_fd_sc_hd__a22o_1
XFILLER_127_1363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30789_ _30789_/A VGND VGND VPWR VPWR _35627_/D sky130_fd_sc_hd__clkbuf_1
X_33577_ _33897_/CLK _33577_/D VGND VGND VPWR VPWR _33577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20542_ _18348_/X _20540_/X _20541_/X _18358_/X VGND VGND VPWR VPWR _20542_/X sky130_fd_sc_hd__a22o_1
X_23330_ _23330_/A VGND VGND VPWR VPWR _32182_/D sky130_fd_sc_hd__clkbuf_1
X_35316_ _35698_/CLK _35316_/D VGND VGND VPWR VPWR _35316_/Q sky130_fd_sc_hd__dfxtp_1
X_32528_ _35985_/CLK _32528_/D VGND VGND VPWR VPWR _32528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20473_ _35730_/Q _32241_/Q _35602_/Q _35538_/Q _18293_/X _18295_/X VGND VGND VPWR
+ VPWR _20473_/X sky130_fd_sc_hd__mux4_1
X_35247_ _35438_/CLK _35247_/D VGND VGND VPWR VPWR _35247_/Q sky130_fd_sc_hd__dfxtp_1
X_23261_ input2/X VGND VGND VPWR VPWR _23261_/X sky130_fd_sc_hd__buf_4
X_32459_ _36079_/CLK _32459_/D VGND VGND VPWR VPWR _32459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25000_ _25000_/A VGND VGND VPWR VPWR _32982_/D sky130_fd_sc_hd__clkbuf_1
X_22212_ _22206_/X _22211_/X _22104_/X VGND VGND VPWR VPWR _22220_/C sky130_fd_sc_hd__o21ba_1
XFILLER_152_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23192_ _23036_/X _32134_/Q _23194_/S VGND VGND VPWR VPWR _23193_/A sky130_fd_sc_hd__mux2_1
X_35178_ _35564_/CLK _35178_/D VGND VGND VPWR VPWR _35178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22143_ _34687_/Q _34623_/Q _34559_/Q _34495_/Q _21892_/X _21893_/X VGND VGND VPWR
+ VPWR _22143_/X sky130_fd_sc_hd__mux4_1
X_34129_ _34193_/CLK _34129_/D VGND VGND VPWR VPWR _34129_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26951_ _26951_/A VGND VGND VPWR VPWR _33902_/D sky130_fd_sc_hd__clkbuf_1
X_22074_ _22070_/X _22073_/X _21765_/X VGND VGND VPWR VPWR _22075_/D sky130_fd_sc_hd__o21ba_1
XTAP_6739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25902_ _24930_/X _33408_/Q _25916_/S VGND VGND VPWR VPWR _25903_/A sky130_fd_sc_hd__mux2_1
X_21025_ _20747_/X _21023_/X _21024_/X _20750_/X VGND VGND VPWR VPWR _21025_/X sky130_fd_sc_hd__a22o_1
XFILLER_87_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_247_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29670_ _35097_/Q _29339_/X _29682_/S VGND VGND VPWR VPWR _29671_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26882_ _33870_/Q _23475_/X _26888_/S VGND VGND VPWR VPWR _26883_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_908 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_248_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28621_ _28648_/S VGND VGND VPWR VPWR _28640_/S sky130_fd_sc_hd__buf_4
XFILLER_47_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25833_ _25833_/A VGND VGND VPWR VPWR _33375_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_417_CLK clkbuf_6_32__f_CLK/X VGND VGND VPWR VPWR _35567_/CLK sky130_fd_sc_hd__clkbuf_16
X_28552_ _27695_/X _34599_/Q _28556_/S VGND VGND VPWR VPWR _28553_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25764_ _25764_/A VGND VGND VPWR VPWR _33342_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22976_ _22976_/A VGND VGND VPWR VPWR _32050_/D sky130_fd_sc_hd__clkbuf_1
X_27503_ _27503_/A VGND VGND VPWR VPWR _34133_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_215_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24715_ _22965_/X _32879_/Q _24723_/S VGND VGND VPWR VPWR _24716_/A sky130_fd_sc_hd__mux2_1
XFILLER_243_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28483_ _28483_/A VGND VGND VPWR VPWR _34566_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21927_ _35193_/Q _35129_/Q _35065_/Q _32249_/Q _21610_/X _21611_/X VGND VGND VPWR
+ VPWR _21927_/X sky130_fd_sc_hd__mux4_1
X_25695_ _24824_/X _33310_/Q _25697_/S VGND VGND VPWR VPWR _25696_/A sky130_fd_sc_hd__mux2_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_607 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27434_ _34100_/Q _27127_/X _27452_/S VGND VGND VPWR VPWR _27435_/A sky130_fd_sc_hd__mux2_1
X_24646_ _24646_/A VGND VGND VPWR VPWR _32846_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21858_ _21603_/X _21856_/X _21857_/X _21606_/X VGND VGND VPWR VPWR _21858_/X sky130_fd_sc_hd__a22o_1
XFILLER_187_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27365_ _34068_/Q _27226_/X _27367_/S VGND VGND VPWR VPWR _27366_/A sky130_fd_sc_hd__mux2_1
XFILLER_208_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20809_ _20809_/A VGND VGND VPWR VPWR _36185_/D sky130_fd_sc_hd__clkbuf_2
X_24577_ _24577_/A VGND VGND VPWR VPWR _32813_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_208_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21789_ _21785_/X _21788_/X _21751_/X VGND VGND VPWR VPWR _21797_/C sky130_fd_sc_hd__o21ba_1
XFILLER_23_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29104_ _34859_/Q _27100_/X _29120_/S VGND VGND VPWR VPWR _29105_/A sky130_fd_sc_hd__mux2_1
X_26316_ _26316_/A VGND VGND VPWR VPWR _33604_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_204_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23528_ _32259_/Q _23438_/X _23536_/S VGND VGND VPWR VPWR _23529_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27296_ _34035_/Q _27124_/X _27296_/S VGND VGND VPWR VPWR _27297_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29035_ _29035_/A VGND VGND VPWR VPWR _34826_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_587 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26247_ _26247_/A VGND VGND VPWR VPWR _33571_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23459_ _23459_/A VGND VGND VPWR VPWR _32231_/D sky130_fd_sc_hd__clkbuf_1
X_16000_ _17773_/A VGND VGND VPWR VPWR _17864_/A sky130_fd_sc_hd__buf_12
XFILLER_221_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26178_ _24939_/X _33539_/Q _26186_/S VGND VGND VPWR VPWR _26179_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_1057 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25129_ _25129_/A VGND VGND VPWR VPWR _33044_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29937_ _29937_/A VGND VGND VPWR VPWR _35223_/D sky130_fd_sc_hd__clkbuf_1
X_17951_ _33163_/Q _36043_/Q _33035_/Q _32971_/Q _17768_/X _17769_/X VGND VGND VPWR
+ VPWR _17951_/X sky130_fd_sc_hd__mux4_1
XFILLER_124_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16902_ _17961_/A VGND VGND VPWR VPWR _16902_/X sky130_fd_sc_hd__buf_4
X_17882_ _32649_/Q _32585_/Q _32521_/Q _35977_/Q _17629_/X _17766_/X VGND VGND VPWR
+ VPWR _17882_/X sky130_fd_sc_hd__mux4_1
XFILLER_26_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29868_ _35191_/Q _29432_/X _29880_/S VGND VGND VPWR VPWR _29869_/A sky130_fd_sc_hd__mux2_1
X_19621_ _19298_/X _19619_/X _19620_/X _19301_/X VGND VGND VPWR VPWR _19621_/X sky130_fd_sc_hd__a22o_1
XFILLER_38_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28819_ _34724_/Q _27078_/X _28829_/S VGND VGND VPWR VPWR _28820_/A sky130_fd_sc_hd__mux2_1
X_16833_ _35435_/Q _35371_/Q _35307_/Q _35243_/Q _16548_/X _16549_/X VGND VGND VPWR
+ VPWR _16833_/X sky130_fd_sc_hd__mux4_1
XFILLER_226_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29799_ _35158_/Q _29328_/X _29817_/S VGND VGND VPWR VPWR _29800_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_408_CLK clkbuf_6_34__f_CLK/X VGND VGND VPWR VPWR _34099_/CLK sky130_fd_sc_hd__clkbuf_16
X_31830_ _31830_/A VGND VGND VPWR VPWR _36120_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19552_ _35639_/Q _34999_/Q _34359_/Q _33719_/Q _19444_/X _19445_/X VGND VGND VPWR
+ VPWR _19552_/X sky130_fd_sc_hd__mux4_1
X_16764_ _16447_/X _16762_/X _16763_/X _16450_/X VGND VGND VPWR VPWR _16764_/X sky130_fd_sc_hd__a22o_1
XFILLER_65_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_1240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18503_ _18378_/X _18501_/X _18502_/X _18388_/X VGND VGND VPWR VPWR _18503_/X sky130_fd_sc_hd__a22o_1
XFILLER_18_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31761_ _36088_/Q input28/X _31771_/S VGND VGND VPWR VPWR _31762_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19483_ _35701_/Q _32210_/Q _35573_/Q _35509_/Q _19264_/X _19265_/X VGND VGND VPWR
+ VPWR _19483_/X sky130_fd_sc_hd__mux4_1
X_16695_ _16452_/X _16693_/X _16694_/X _16457_/X VGND VGND VPWR VPWR _16695_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30712_ _30712_/A VGND VGND VPWR VPWR _35591_/D sky130_fd_sc_hd__clkbuf_1
X_33500_ _36211_/CLK _33500_/D VGND VGND VPWR VPWR _33500_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18434_ _34391_/Q _36119_/Q _34263_/Q _34199_/Q _18392_/X _18394_/X VGND VGND VPWR
+ VPWR _18434_/X sky130_fd_sc_hd__mux4_1
XFILLER_178_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31692_ _36055_/Q input12/X _31708_/S VGND VGND VPWR VPWR _31693_/A sky130_fd_sc_hd__mux2_1
X_34480_ _34927_/CLK _34480_/D VGND VGND VPWR VPWR _34480_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18365_ _35414_/Q _35350_/Q _35286_/Q _35222_/Q _18362_/X _18364_/X VGND VGND VPWR
+ VPWR _18365_/X sky130_fd_sc_hd__mux4_1
X_33431_ _35995_/CLK _33431_/D VGND VGND VPWR VPWR _33431_/Q sky130_fd_sc_hd__dfxtp_1
X_30643_ _30643_/A VGND VGND VPWR VPWR _35558_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17316_ _17312_/X _17315_/X _17140_/X _17141_/X VGND VGND VPWR VPWR _17333_/B sky130_fd_sc_hd__o211a_1
X_33362_ _36179_/CLK _33362_/D VGND VGND VPWR VPWR _33362_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36150_ _36150_/CLK _36150_/D VGND VGND VPWR VPWR _36150_/Q sky130_fd_sc_hd__dfxtp_1
X_18296_ _34134_/Q _34070_/Q _34006_/Q _33942_/Q _18293_/X _18295_/X VGND VGND VPWR
+ VPWR _18296_/X sky130_fd_sc_hd__mux4_1
X_30574_ _35526_/Q _29478_/X _30576_/S VGND VGND VPWR VPWR _30575_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35101_ _36219_/CLK _35101_/D VGND VGND VPWR VPWR _35101_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_857 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17247_ _32119_/Q _32311_/Q _32375_/Q _35895_/Q _16927_/X _17068_/X VGND VGND VPWR
+ VPWR _17247_/X sky130_fd_sc_hd__mux4_1
X_32313_ _32889_/CLK _32313_/D VGND VGND VPWR VPWR _32313_/Q sky130_fd_sc_hd__dfxtp_1
X_33293_ _34186_/CLK _33293_/D VGND VGND VPWR VPWR _33293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36081_ _36082_/CLK _36081_/D VGND VGND VPWR VPWR _36081_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35032_ _35162_/CLK _35032_/D VGND VGND VPWR VPWR _35032_/Q sky130_fd_sc_hd__dfxtp_1
X_32244_ _35733_/CLK _32244_/D VGND VGND VPWR VPWR _32244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17178_ _17059_/X _17176_/X _17177_/X _17065_/X VGND VGND VPWR VPWR _17178_/X sky130_fd_sc_hd__a22o_1
XFILLER_157_1312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16129_ _16060_/X _16127_/X _16128_/X _16072_/X VGND VGND VPWR VPWR _16129_/X sky130_fd_sc_hd__a22o_1
X_32175_ _35735_/CLK _32175_/D VGND VGND VPWR VPWR _32175_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31126_ _31126_/A VGND VGND VPWR VPWR _35787_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35934_ _35998_/CLK _35934_/D VGND VGND VPWR VPWR _35934_/Q sky130_fd_sc_hd__dfxtp_1
X_31057_ _31057_/A VGND VGND VPWR VPWR _35754_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30008_ _30008_/A VGND VGND VPWR VPWR _35257_/D sky130_fd_sc_hd__clkbuf_1
X_19819_ _19810_/X _19817_/X _19818_/X VGND VGND VPWR VPWR _19820_/D sky130_fd_sc_hd__o21ba_1
XFILLER_110_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35865_ _35865_/CLK _35865_/D VGND VGND VPWR VPWR _35865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34816_ _36104_/CLK _34816_/D VGND VGND VPWR VPWR _34816_/Q sky130_fd_sc_hd__dfxtp_1
X_22830_ _32916_/Q _32852_/Q _32788_/Q _32724_/Q _20584_/X _20587_/X VGND VGND VPWR
+ VPWR _22830_/X sky130_fd_sc_hd__mux4_1
XFILLER_56_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35796_ _35860_/CLK _35796_/D VGND VGND VPWR VPWR _35796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22761_ _22505_/X _22759_/X _22760_/X _22510_/X VGND VGND VPWR VPWR _22761_/X sky130_fd_sc_hd__a22o_1
X_34747_ _34877_/CLK _34747_/D VGND VGND VPWR VPWR _34747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31959_ _34148_/CLK _31959_/D VGND VGND VPWR VPWR _31959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24500_ _23046_/X _32777_/Q _24516_/S VGND VGND VPWR VPWR _24501_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21712_ _33075_/Q _32051_/Q _35827_/Q _35763_/Q _21678_/X _21679_/X VGND VGND VPWR
+ VPWR _21712_/X sky130_fd_sc_hd__mux4_1
XFILLER_225_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25480_ _24905_/X _33208_/Q _25490_/S VGND VGND VPWR VPWR _25481_/A sky130_fd_sc_hd__mux2_1
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_747 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22692_ _22459_/X _22690_/X _22691_/X _22462_/X VGND VGND VPWR VPWR _22692_/X sky130_fd_sc_hd__a22o_1
X_34678_ _35126_/CLK _34678_/D VGND VGND VPWR VPWR _34678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24431_ _24431_/A VGND VGND VPWR VPWR _32744_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33629_ _36205_/CLK _33629_/D VGND VGND VPWR VPWR _33629_/Q sky130_fd_sc_hd__dfxtp_1
X_21643_ _34673_/Q _34609_/Q _34545_/Q _34481_/Q _21539_/X _21540_/X VGND VGND VPWR
+ VPWR _21643_/X sky130_fd_sc_hd__mux4_1
XFILLER_244_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27150_ _33979_/Q _27149_/X _27156_/S VGND VGND VPWR VPWR _27151_/A sky130_fd_sc_hd__mux2_1
X_24362_ _24389_/S VGND VGND VPWR VPWR _24381_/S sky130_fd_sc_hd__buf_4
X_21574_ _35183_/Q _35119_/Q _35055_/Q _32176_/Q _21257_/X _21258_/X VGND VGND VPWR
+ VPWR _21574_/X sky130_fd_sc_hd__mux4_1
XFILLER_138_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26101_ _26101_/A VGND VGND VPWR VPWR _33502_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23313_ _23499_/S VGND VGND VPWR VPWR _23335_/S sky130_fd_sc_hd__buf_6
X_20525_ _20521_/X _20524_/X _20138_/A VGND VGND VPWR VPWR _20547_/A sky130_fd_sc_hd__o21ba_1
X_27081_ input7/X VGND VGND VPWR VPWR _27081_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_20_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24293_ _22940_/X _32679_/Q _24297_/S VGND VGND VPWR VPWR _24294_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26032_ _26080_/S VGND VGND VPWR VPWR _26051_/S sky130_fd_sc_hd__buf_6
XFILLER_10_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23244_ _32154_/Q _23243_/X _23259_/S VGND VGND VPWR VPWR _23245_/A sky130_fd_sc_hd__mux2_1
X_20456_ _20452_/X _20455_/X _20171_/X VGND VGND VPWR VPWR _20457_/D sky130_fd_sc_hd__o21ba_1
XFILLER_140_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20387_ _33103_/Q _32079_/Q _35855_/Q _35791_/Q _20084_/X _20085_/X VGND VGND VPWR
+ VPWR _20387_/X sky130_fd_sc_hd__mux4_1
X_23175_ _23223_/S VGND VGND VPWR VPWR _23194_/S sky130_fd_sc_hd__buf_4
XFILLER_122_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22126_ _33919_/Q _33855_/Q _33791_/Q _36095_/Q _21977_/X _21978_/X VGND VGND VPWR
+ VPWR _22126_/X sky130_fd_sc_hd__mux4_1
XFILLER_136_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27983_ _34329_/Q _27044_/X _27995_/S VGND VGND VPWR VPWR _27984_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput170 _36206_/Q VGND VGND VPWR VPWR D2[24] sky130_fd_sc_hd__buf_2
XFILLER_121_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput181 _36216_/Q VGND VGND VPWR VPWR D2[34] sky130_fd_sc_hd__buf_2
XFILLER_82_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput192 _36226_/Q VGND VGND VPWR VPWR D2[44] sky130_fd_sc_hd__buf_2
XTAP_5802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26934_ _26934_/A VGND VGND VPWR VPWR _33894_/D sky130_fd_sc_hd__clkbuf_1
X_29722_ _35122_/Q _29416_/X _29724_/S VGND VGND VPWR VPWR _29723_/A sky130_fd_sc_hd__mux2_1
XTAP_6569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22057_ _32125_/Q _32317_/Q _32381_/Q _35901_/Q _21880_/X _22021_/X VGND VGND VPWR
+ VPWR _22057_/X sky130_fd_sc_hd__mux4_1
XFILLER_82_1063 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21008_ _21004_/X _21007_/X _20675_/X VGND VGND VPWR VPWR _21016_/C sky130_fd_sc_hd__o21ba_1
XFILLER_102_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29653_ _29653_/A VGND VGND VPWR VPWR _35089_/D sky130_fd_sc_hd__clkbuf_1
X_26865_ _33862_/Q _23447_/X _26867_/S VGND VGND VPWR VPWR _26866_/A sky130_fd_sc_hd__mux2_1
XTAP_5868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28604_ _28604_/A VGND VGND VPWR VPWR _34623_/D sky130_fd_sc_hd__clkbuf_1
X_25816_ _24803_/X _33367_/Q _25832_/S VGND VGND VPWR VPWR _25817_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29584_ _29584_/A VGND VGND VPWR VPWR _35056_/D sky130_fd_sc_hd__clkbuf_1
X_26796_ _33829_/Q _23277_/X _26804_/S VGND VGND VPWR VPWR _26797_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28535_ _27670_/X _34591_/Q _28535_/S VGND VGND VPWR VPWR _28536_/A sky130_fd_sc_hd__mux2_1
X_25747_ _25747_/A VGND VGND VPWR VPWR _33334_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_216_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22959_ input16/X VGND VGND VPWR VPWR _22959_/X sky130_fd_sc_hd__buf_2
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_243_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28466_ _27766_/X _34558_/Q _28484_/S VGND VGND VPWR VPWR _28467_/A sky130_fd_sc_hd__mux2_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16480_ _35425_/Q _35361_/Q _35297_/Q _35233_/Q _16195_/X _16196_/X VGND VGND VPWR
+ VPWR _16480_/X sky130_fd_sc_hd__mux4_1
XFILLER_189_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25678_ _25810_/S VGND VGND VPWR VPWR _25697_/S sky130_fd_sc_hd__buf_4
XFILLER_243_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27417_ _34092_/Q _27103_/X _27431_/S VGND VGND VPWR VPWR _27418_/A sky130_fd_sc_hd__mux2_1
X_24629_ _24629_/A VGND VGND VPWR VPWR _32838_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_223_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28397_ _28397_/A VGND VGND VPWR VPWR _34525_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_1132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18150_ _34705_/Q _34641_/Q _34577_/Q _34513_/Q _17998_/X _17999_/X VGND VGND VPWR
+ VPWR _18150_/X sky130_fd_sc_hd__mux4_1
X_27348_ _27348_/A VGND VGND VPWR VPWR _34059_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17101_ _32627_/Q _32563_/Q _32499_/Q _35955_/Q _16923_/X _17060_/X VGND VGND VPWR
+ VPWR _17101_/X sky130_fd_sc_hd__mux4_1
XFILLER_50_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18081_ _17773_/X _18079_/X _18080_/X _17777_/X VGND VGND VPWR VPWR _18081_/X sky130_fd_sc_hd__a22o_1
XFILLER_7_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27279_ _27279_/A VGND VGND VPWR VPWR _34026_/D sky130_fd_sc_hd__clkbuf_1
X_29018_ _29018_/A VGND VGND VPWR VPWR _34818_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_1463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17032_ _32113_/Q _32305_/Q _32369_/Q _35889_/Q _16927_/X _16715_/X VGND VGND VPWR
+ VPWR _17032_/X sky130_fd_sc_hd__mux4_1
XFILLER_156_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30290_ _35391_/Q _29457_/X _30306_/S VGND VGND VPWR VPWR _30291_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18983_ _35687_/Q _32194_/Q _35559_/Q _35495_/Q _18911_/X _18912_/X VGND VGND VPWR
+ VPWR _18983_/X sky130_fd_sc_hd__mux4_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17934_ _17859_/X _17932_/X _17933_/X _17862_/X VGND VGND VPWR VPWR _17934_/X sky130_fd_sc_hd__a22o_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33980_ _35449_/CLK _33980_/D VGND VGND VPWR VPWR _33980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32931_ _36005_/CLK _32931_/D VGND VGND VPWR VPWR _32931_/Q sky130_fd_sc_hd__dfxtp_1
X_17865_ _34440_/Q _36168_/Q _34312_/Q _34248_/Q _17582_/X _17583_/X VGND VGND VPWR
+ VPWR _17865_/X sky130_fd_sc_hd__mux4_1
XFILLER_26_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19604_ _34169_/Q _34105_/Q _34041_/Q _33977_/Q _19393_/X _19394_/X VGND VGND VPWR
+ VPWR _19604_/X sky130_fd_sc_hd__mux4_1
XFILLER_4_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35650_ _35777_/CLK _35650_/D VGND VGND VPWR VPWR _35650_/Q sky130_fd_sc_hd__dfxtp_1
X_16816_ _33643_/Q _33579_/Q _33515_/Q _33451_/Q _16494_/X _16495_/X VGND VGND VPWR
+ VPWR _16816_/X sky130_fd_sc_hd__mux4_1
X_32862_ _35989_/CLK _32862_/D VGND VGND VPWR VPWR _32862_/Q sky130_fd_sc_hd__dfxtp_1
X_17796_ _17796_/A _17796_/B _17796_/C _17796_/D VGND VGND VPWR VPWR _17797_/A sky130_fd_sc_hd__or4_1
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_219_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34601_ _34913_/CLK _34601_/D VGND VGND VPWR VPWR _34601_/Q sky130_fd_sc_hd__dfxtp_1
X_31813_ _36113_/Q input55/X _31813_/S VGND VGND VPWR VPWR _31814_/A sky130_fd_sc_hd__mux2_1
X_19535_ _19535_/A _19535_/B _19535_/C _19535_/D VGND VGND VPWR VPWR _19536_/A sky130_fd_sc_hd__or4_1
XFILLER_93_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16747_ _16743_/X _16746_/X _16426_/X VGND VGND VPWR VPWR _16769_/A sky130_fd_sc_hd__o21ba_1
X_35581_ _35581_/CLK _35581_/D VGND VGND VPWR VPWR _35581_/Q sky130_fd_sc_hd__dfxtp_1
X_32793_ _34070_/CLK _32793_/D VGND VGND VPWR VPWR _32793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34532_ _35490_/CLK _34532_/D VGND VGND VPWR VPWR _34532_/Q sky130_fd_sc_hd__dfxtp_1
X_31744_ _36080_/Q input19/X _31750_/S VGND VGND VPWR VPWR _31745_/A sky130_fd_sc_hd__mux2_1
X_19466_ _19457_/X _19464_/X _19465_/X VGND VGND VPWR VPWR _19467_/D sky130_fd_sc_hd__o21ba_1
X_16678_ _16353_/X _16676_/X _16677_/X _16359_/X VGND VGND VPWR VPWR _16678_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18417_ _32599_/Q _32535_/Q _32471_/Q _35927_/Q _20166_/A _20017_/A VGND VGND VPWR
+ VPWR _18417_/X sky130_fd_sc_hd__mux4_1
XFILLER_210_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34463_ _35544_/CLK _34463_/D VGND VGND VPWR VPWR _34463_/Q sky130_fd_sc_hd__dfxtp_1
X_31675_ _31675_/A VGND VGND VPWR VPWR _36047_/D sky130_fd_sc_hd__clkbuf_1
X_19397_ _33395_/Q _33331_/Q _33267_/Q _33203_/Q _19074_/X _19075_/X VGND VGND VPWR
+ VPWR _19397_/X sky130_fd_sc_hd__mux4_1
XFILLER_210_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36202_ _36202_/CLK _36202_/D VGND VGND VPWR VPWR _36202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33414_ _33415_/CLK _33414_/D VGND VGND VPWR VPWR _33414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18348_ _20159_/A VGND VGND VPWR VPWR _18348_/X sky130_fd_sc_hd__clkbuf_4
X_30626_ _30626_/A VGND VGND VPWR VPWR _35550_/D sky130_fd_sc_hd__clkbuf_1
X_34394_ _36235_/CLK _34394_/D VGND VGND VPWR VPWR _34394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36133_ _36136_/CLK _36133_/D VGND VGND VPWR VPWR _36133_/Q sky130_fd_sc_hd__dfxtp_1
X_33345_ _33924_/CLK _33345_/D VGND VGND VPWR VPWR _33345_/Q sky130_fd_sc_hd__dfxtp_1
X_30557_ _30605_/S VGND VGND VPWR VPWR _30576_/S sky130_fd_sc_hd__buf_6
X_18279_ input79/X input80/X VGND VGND VPWR VPWR _20065_/A sky130_fd_sc_hd__nor2b_4
X_20310_ _34189_/Q _34125_/Q _34061_/Q _33997_/Q _20099_/X _20100_/X VGND VGND VPWR
+ VPWR _20310_/X sky130_fd_sc_hd__mux4_1
XFILLER_200_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput50 DW[54] VGND VGND VPWR VPWR input50/X sky130_fd_sc_hd__buf_8
X_36064_ _36065_/CLK _36064_/D VGND VGND VPWR VPWR _36064_/Q sky130_fd_sc_hd__dfxtp_1
X_21290_ _34663_/Q _34599_/Q _34535_/Q _34471_/Q _21186_/X _21187_/X VGND VGND VPWR
+ VPWR _21290_/X sky130_fd_sc_hd__mux4_1
X_30488_ _35485_/Q _29351_/X _30492_/S VGND VGND VPWR VPWR _30489_/A sky130_fd_sc_hd__mux2_1
X_33276_ _33531_/CLK _33276_/D VGND VGND VPWR VPWR _33276_/Q sky130_fd_sc_hd__dfxtp_1
Xinput61 DW[6] VGND VGND VPWR VPWR input61/X sky130_fd_sc_hd__buf_6
Xinput72 R2[1] VGND VGND VPWR VPWR input72/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput83 RW[0] VGND VGND VPWR VPWR input83/X sky130_fd_sc_hd__clkbuf_4
X_20241_ _20241_/A _20241_/B _20241_/C _20241_/D VGND VGND VPWR VPWR _20242_/A sky130_fd_sc_hd__or4_2
X_35015_ _35715_/CLK _35015_/D VGND VGND VPWR VPWR _35015_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32227_ _35525_/CLK _32227_/D VGND VGND VPWR VPWR _32227_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20172_ _20163_/X _20170_/X _20171_/X VGND VGND VPWR VPWR _20173_/D sky130_fd_sc_hd__o21ba_1
X_32158_ _36223_/CLK _32158_/D VGND VGND VPWR VPWR _32158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31109_ _31109_/A VGND VGND VPWR VPWR _35779_/D sky130_fd_sc_hd__clkbuf_1
X_32089_ _35733_/CLK _32089_/D VGND VGND VPWR VPWR _32089_/Q sky130_fd_sc_hd__dfxtp_1
X_24980_ _24979_/X _32976_/Q _24983_/S VGND VGND VPWR VPWR _24981_/A sky130_fd_sc_hd__mux2_1
XFILLER_229_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_233_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35917_ _35983_/CLK _35917_/D VGND VGND VPWR VPWR _35917_/Q sky130_fd_sc_hd__dfxtp_1
X_23931_ _23931_/A VGND VGND VPWR VPWR _32510_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26650_ _26761_/S VGND VGND VPWR VPWR _26669_/S sky130_fd_sc_hd__buf_4
X_35848_ _35849_/CLK _35848_/D VGND VGND VPWR VPWR _35848_/Q sky130_fd_sc_hd__dfxtp_1
X_23862_ _22912_/X _32478_/Q _23864_/S VGND VGND VPWR VPWR _23863_/A sky130_fd_sc_hd__mux2_1
XTAP_3729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25601_ _25601_/A VGND VGND VPWR VPWR _33265_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22813_ _34451_/Q _36179_/Q _34323_/Q _34259_/Q _22535_/X _22536_/X VGND VGND VPWR
+ VPWR _22813_/X sky130_fd_sc_hd__mux4_1
XFILLER_26_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26581_ _24933_/X _33729_/Q _26593_/S VGND VGND VPWR VPWR _26582_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35779_ _35779_/CLK _35779_/D VGND VGND VPWR VPWR _35779_/Q sky130_fd_sc_hd__dfxtp_1
X_23793_ _23011_/X _32382_/Q _23811_/S VGND VGND VPWR VPWR _23794_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28320_ _27751_/X _34489_/Q _28328_/S VGND VGND VPWR VPWR _28321_/A sky130_fd_sc_hd__mux2_1
X_25532_ _24982_/X _33233_/Q _25532_/S VGND VGND VPWR VPWR _25533_/A sky130_fd_sc_hd__mux2_1
X_22744_ _35665_/Q _35025_/Q _34385_/Q _33745_/Q _22450_/X _22451_/X VGND VGND VPWR
+ VPWR _22744_/X sky130_fd_sc_hd__mux4_1
XFILLER_73_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28251_ _27649_/X _34456_/Q _28265_/S VGND VGND VPWR VPWR _28252_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25463_ _24880_/X _33200_/Q _25469_/S VGND VGND VPWR VPWR _25464_/A sky130_fd_sc_hd__mux2_1
X_22675_ _22671_/X _22674_/X _22438_/X VGND VGND VPWR VPWR _22697_/A sky130_fd_sc_hd__o21ba_1
XFILLER_12_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27202_ input50/X VGND VGND VPWR VPWR _27202_/X sky130_fd_sc_hd__buf_4
XFILLER_200_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24414_ _22918_/X _32736_/Q _24432_/S VGND VGND VPWR VPWR _24415_/A sky130_fd_sc_hd__mux2_1
X_21626_ _33905_/Q _33841_/Q _33777_/Q _36081_/Q _21624_/X _21625_/X VGND VGND VPWR
+ VPWR _21626_/X sky130_fd_sc_hd__mux4_1
XFILLER_40_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28182_ _28182_/A VGND VGND VPWR VPWR _34423_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_1192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25394_ _25394_/A VGND VGND VPWR VPWR _33168_/D sky130_fd_sc_hd__clkbuf_1
X_27133_ _27133_/A VGND VGND VPWR VPWR _33973_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_1018 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24345_ _24345_/A VGND VGND VPWR VPWR _32703_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21557_ _32623_/Q _32559_/Q _32495_/Q _35951_/Q _21523_/X _21307_/X VGND VGND VPWR
+ VPWR _21557_/X sky130_fd_sc_hd__mux4_1
X_20508_ _18301_/X _20506_/X _20507_/X _18307_/X VGND VGND VPWR VPWR _20508_/X sky130_fd_sc_hd__a22o_1
X_27064_ _27064_/A VGND VGND VPWR VPWR _33951_/D sky130_fd_sc_hd__clkbuf_1
X_24276_ _22915_/X _32671_/Q _24276_/S VGND VGND VPWR VPWR _24277_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21488_ _33901_/Q _33837_/Q _33773_/Q _36077_/Q _21271_/X _21272_/X VGND VGND VPWR
+ VPWR _21488_/X sky130_fd_sc_hd__mux4_1
X_26015_ _26015_/A VGND VGND VPWR VPWR _33461_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23227_ _23227_/A VGND VGND VPWR VPWR _29797_/A sky130_fd_sc_hd__buf_12
XFILLER_4_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20439_ _32145_/Q _32337_/Q _32401_/Q _35921_/Q _20286_/X _19311_/A VGND VGND VPWR
+ VPWR _20439_/X sky130_fd_sc_hd__mux4_1
XFILLER_10_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23158_ _23158_/A VGND VGND VPWR VPWR _32117_/D sky130_fd_sc_hd__clkbuf_1
XTAP_7056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22109_ _22462_/A VGND VGND VPWR VPWR _22109_/X sky130_fd_sc_hd__clkbuf_4
XTAP_7089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15980_ _17765_/A VGND VGND VPWR VPWR _17859_/A sky130_fd_sc_hd__buf_12
X_27966_ _27966_/A VGND VGND VPWR VPWR _34321_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23089_ _23089_/A VGND VGND VPWR VPWR _28110_/A sky130_fd_sc_hd__buf_6
XTAP_6366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29705_ _29795_/S VGND VGND VPWR VPWR _29724_/S sky130_fd_sc_hd__buf_6
XFILLER_76_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26917_ _26917_/A VGND VGND VPWR VPWR _33886_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27897_ _27897_/A VGND VGND VPWR VPWR _34288_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17650_ _34434_/Q _36162_/Q _34306_/Q _34242_/Q _17582_/X _17583_/X VGND VGND VPWR
+ VPWR _17650_/X sky130_fd_sc_hd__mux4_1
X_29636_ _35081_/Q _29488_/X _29652_/S VGND VGND VPWR VPWR _29637_/A sky130_fd_sc_hd__mux2_1
XTAP_5698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26848_ _26896_/S VGND VGND VPWR VPWR _26867_/S sky130_fd_sc_hd__buf_6
XTAP_4964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_1180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16601_ _33893_/Q _33829_/Q _33765_/Q _36069_/Q _16318_/X _16319_/X VGND VGND VPWR
+ VPWR _16601_/X sky130_fd_sc_hd__mux4_1
X_17581_ _17506_/X _17579_/X _17580_/X _17509_/X VGND VGND VPWR VPWR _17581_/X sky130_fd_sc_hd__a22o_1
XTAP_4997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26779_ _33821_/Q _23252_/X _26783_/S VGND VGND VPWR VPWR _26780_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29567_ _29567_/A VGND VGND VPWR VPWR _35048_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19320_ _33649_/Q _33585_/Q _33521_/Q _33457_/Q _19147_/X _19148_/X VGND VGND VPWR
+ VPWR _19320_/X sky130_fd_sc_hd__mux4_1
X_16532_ _34147_/Q _34083_/Q _34019_/Q _33955_/Q _16387_/X _16388_/X VGND VGND VPWR
+ VPWR _16532_/X sky130_fd_sc_hd__mux4_1
XFILLER_73_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28518_ _28518_/A VGND VGND VPWR VPWR _34582_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29498_ _35020_/Q _29497_/X _29513_/S VGND VGND VPWR VPWR _29499_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19251_ _34159_/Q _34095_/Q _34031_/Q _33967_/Q _19040_/X _19041_/X VGND VGND VPWR
+ VPWR _19251_/X sky130_fd_sc_hd__mux4_1
XFILLER_108_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16463_ _33633_/Q _33569_/Q _33505_/Q _33441_/Q _16141_/X _16142_/X VGND VGND VPWR
+ VPWR _16463_/X sky130_fd_sc_hd__mux4_1
X_28449_ _27742_/X _34550_/Q _28463_/S VGND VGND VPWR VPWR _28450_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_223_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18202_ _18198_/X _18201_/X _17846_/A _17847_/A VGND VGND VPWR VPWR _18217_/B sky130_fd_sc_hd__o211a_1
XFILLER_231_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19182_ _19182_/A _19182_/B _19182_/C _19182_/D VGND VGND VPWR VPWR _19183_/A sky130_fd_sc_hd__or4_4
X_31460_ _31460_/A VGND VGND VPWR VPWR _35945_/D sky130_fd_sc_hd__clkbuf_1
XPHY_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16394_ _16390_/X _16393_/X _16015_/X VGND VGND VPWR VPWR _16416_/A sky130_fd_sc_hd__o21ba_1
XPHY_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18133_ _33937_/Q _33873_/Q _33809_/Q _36113_/Q _16062_/X _16064_/X VGND VGND VPWR
+ VPWR _18133_/X sky130_fd_sc_hd__mux4_1
X_30411_ _30411_/A VGND VGND VPWR VPWR _35448_/D sky130_fd_sc_hd__clkbuf_1
X_31391_ _31391_/A VGND VGND VPWR VPWR _35912_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18064_ _34958_/Q _34894_/Q _34830_/Q _34766_/Q _17866_/X _17867_/X VGND VGND VPWR
+ VPWR _18064_/X sky130_fd_sc_hd__mux4_1
X_30342_ _30342_/A VGND VGND VPWR VPWR _35415_/D sky130_fd_sc_hd__clkbuf_1
X_33130_ _36141_/CLK _33130_/D VGND VGND VPWR VPWR _33130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_890 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17015_ _34928_/Q _34864_/Q _34800_/Q _34736_/Q _16807_/X _16808_/X VGND VGND VPWR
+ VPWR _17015_/X sky130_fd_sc_hd__mux4_1
XFILLER_208_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33061_ _35814_/CLK _33061_/D VGND VGND VPWR VPWR _33061_/Q sky130_fd_sc_hd__dfxtp_1
X_30273_ _35383_/Q _29432_/X _30285_/S VGND VGND VPWR VPWR _30274_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32012_ _36202_/CLK _32012_/D VGND VGND VPWR VPWR _32012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18966_ _18966_/A VGND VGND VPWR VPWR _32422_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_230_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17917_ _17911_/X _17916_/X _17838_/X VGND VGND VPWR VPWR _17941_/A sky130_fd_sc_hd__o21ba_2
XFILLER_113_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33963_ _34091_/CLK _33963_/D VGND VGND VPWR VPWR _33963_/Q sky130_fd_sc_hd__dfxtp_1
X_18897_ _33637_/Q _33573_/Q _33509_/Q _33445_/Q _18794_/X _18795_/X VGND VGND VPWR
+ VPWR _18897_/X sky130_fd_sc_hd__mux4_1
XFILLER_230_1247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35702_ _35703_/CLK _35702_/D VGND VGND VPWR VPWR _35702_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32914_ _32914_/CLK _32914_/D VGND VGND VPWR VPWR _32914_/Q sky130_fd_sc_hd__dfxtp_1
X_17848_ _17842_/X _17845_/X _17846_/X _17847_/X VGND VGND VPWR VPWR _17873_/B sky130_fd_sc_hd__o211a_1
XFILLER_113_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33894_ _36066_/CLK _33894_/D VGND VGND VPWR VPWR _33894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35633_ _35633_/CLK _35633_/D VGND VGND VPWR VPWR _35633_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32845_ _32909_/CLK _32845_/D VGND VGND VPWR VPWR _32845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17779_ _17772_/X _17778_/X _17493_/X _17494_/X VGND VGND VPWR VPWR _17796_/B sky130_fd_sc_hd__o211a_1
XFILLER_54_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19518_ _19514_/X _19517_/X _19440_/X _19441_/X VGND VGND VPWR VPWR _19535_/B sky130_fd_sc_hd__o211a_1
X_35564_ _35564_/CLK _35564_/D VGND VGND VPWR VPWR _35564_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20790_ _20630_/X _20788_/X _20789_/X _20641_/X VGND VGND VPWR VPWR _20790_/X sky130_fd_sc_hd__a22o_1
XFILLER_165_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32776_ _32906_/CLK _32776_/D VGND VGND VPWR VPWR _32776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34515_ _36115_/CLK _34515_/D VGND VGND VPWR VPWR _34515_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31727_ _36072_/Q input10/X _31729_/S VGND VGND VPWR VPWR _31728_/A sky130_fd_sc_hd__mux2_1
X_19449_ _33076_/Q _32052_/Q _35828_/Q _35764_/Q _19378_/X _19379_/X VGND VGND VPWR
+ VPWR _19449_/X sky130_fd_sc_hd__mux4_1
XFILLER_62_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35495_ _35624_/CLK _35495_/D VGND VGND VPWR VPWR _35495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34446_ _36176_/CLK _34446_/D VGND VGND VPWR VPWR _34446_/Q sky130_fd_sc_hd__dfxtp_1
X_22460_ _34696_/Q _34632_/Q _34568_/Q _34504_/Q _22245_/X _22246_/X VGND VGND VPWR
+ VPWR _22460_/X sky130_fd_sc_hd__mux4_1
XFILLER_195_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31658_ _31658_/A VGND VGND VPWR VPWR _36039_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21411_ _21405_/X _21406_/X _21409_/X _21410_/X VGND VGND VPWR VPWR _21411_/X sky130_fd_sc_hd__a22o_1
X_30609_ _35542_/Q _29328_/X _30627_/S VGND VGND VPWR VPWR _30610_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_1046 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34377_ _34633_/CLK _34377_/D VGND VGND VPWR VPWR _34377_/Q sky130_fd_sc_hd__dfxtp_1
X_22391_ _22106_/X _22389_/X _22390_/X _22109_/X VGND VGND VPWR VPWR _22391_/X sky130_fd_sc_hd__a22o_1
XFILLER_136_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31589_ _31589_/A VGND VGND VPWR VPWR _36006_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36116_ _36117_/CLK _36116_/D VGND VGND VPWR VPWR _36116_/Q sky130_fd_sc_hd__dfxtp_1
X_24130_ _32603_/Q _23246_/X _24138_/S VGND VGND VPWR VPWR _24131_/A sky130_fd_sc_hd__mux2_1
X_21342_ _34153_/Q _34089_/Q _34025_/Q _33961_/Q _21340_/X _21341_/X VGND VGND VPWR
+ VPWR _21342_/X sky130_fd_sc_hd__mux4_1
XFILLER_11_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33328_ _33904_/CLK _33328_/D VGND VGND VPWR VPWR _33328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36047_ _36047_/CLK _36047_/D VGND VGND VPWR VPWR _36047_/Q sky130_fd_sc_hd__dfxtp_1
X_24061_ _23005_/X _32572_/Q _24063_/S VGND VGND VPWR VPWR _24062_/A sky130_fd_sc_hd__mux2_1
X_33259_ _36075_/CLK _33259_/D VGND VGND VPWR VPWR _33259_/Q sky130_fd_sc_hd__dfxtp_1
X_21273_ _33895_/Q _33831_/Q _33767_/Q _36071_/Q _21271_/X _21272_/X VGND VGND VPWR
+ VPWR _21273_/X sky130_fd_sc_hd__mux4_1
X_23012_ _23083_/S VGND VGND VPWR VPWR _23040_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_116_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20224_ _20220_/X _20223_/X _20146_/X _20147_/X VGND VGND VPWR VPWR _20241_/B sky130_fd_sc_hd__o211a_1
XFILLER_11_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27820_ _27819_/X _34255_/Q _27826_/S VGND VGND VPWR VPWR _27821_/A sky130_fd_sc_hd__mux2_1
X_20155_ _33096_/Q _32072_/Q _35848_/Q _35784_/Q _20084_/X _20085_/X VGND VGND VPWR
+ VPWR _20155_/X sky130_fd_sc_hd__mux4_1
XFILLER_213_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_246_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20086_ _33094_/Q _32070_/Q _35846_/Q _35782_/Q _20084_/X _20085_/X VGND VGND VPWR
+ VPWR _20086_/X sky130_fd_sc_hd__mux4_1
X_24963_ _24963_/A VGND VGND VPWR VPWR _32970_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27751_ input29/X VGND VGND VPWR VPWR _27751_/X sky130_fd_sc_hd__buf_2
XTAP_4216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26702_ _26702_/A VGND VGND VPWR VPWR _33784_/D sky130_fd_sc_hd__clkbuf_1
X_23914_ _23914_/A VGND VGND VPWR VPWR _32502_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27682_ _27682_/A VGND VGND VPWR VPWR _34210_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24894_ _24892_/X _32948_/Q _24921_/S VGND VGND VPWR VPWR _24895_/A sky130_fd_sc_hd__mux2_1
XFILLER_246_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_246_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26633_ _26633_/A VGND VGND VPWR VPWR _33751_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29421_ _29421_/A VGND VGND VPWR VPWR _34995_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23845_ _23977_/S VGND VGND VPWR VPWR _23864_/S sky130_fd_sc_hd__buf_4
XTAP_3559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29352_ _34973_/Q _29351_/X _29358_/S VGND VGND VPWR VPWR _29353_/A sky130_fd_sc_hd__mux2_1
X_26564_ _24908_/X _33721_/Q _26572_/S VGND VGND VPWR VPWR _26565_/A sky130_fd_sc_hd__mux2_1
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23776_ _22987_/X _32374_/Q _23790_/S VGND VGND VPWR VPWR _23777_/A sky130_fd_sc_hd__mux2_1
X_20988_ _22561_/A VGND VGND VPWR VPWR _20988_/X sky130_fd_sc_hd__clkbuf_8
X_25515_ _25515_/A VGND VGND VPWR VPWR _33224_/D sky130_fd_sc_hd__clkbuf_1
X_28303_ _27726_/X _34481_/Q _28307_/S VGND VGND VPWR VPWR _28304_/A sky130_fd_sc_hd__mux2_1
X_22727_ _22727_/A _22727_/B _22727_/C _22727_/D VGND VGND VPWR VPWR _22728_/A sky130_fd_sc_hd__or4_4
X_29283_ _34944_/Q _27165_/X _29297_/S VGND VGND VPWR VPWR _29284_/A sky130_fd_sc_hd__mux2_1
X_26495_ _24806_/X _33688_/Q _26509_/S VGND VGND VPWR VPWR _26496_/A sky130_fd_sc_hd__mux2_1
XFILLER_242_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28234_ _28234_/A VGND VGND VPWR VPWR _34448_/D sky130_fd_sc_hd__clkbuf_1
X_25446_ _24855_/X _33192_/Q _25448_/S VGND VGND VPWR VPWR _25447_/A sky130_fd_sc_hd__mux2_1
X_22658_ _20601_/X _22656_/X _22657_/X _20607_/X VGND VGND VPWR VPWR _22658_/X sky130_fd_sc_hd__a22o_1
XFILLER_199_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21609_ _34672_/Q _34608_/Q _34544_/Q _34480_/Q _21539_/X _21540_/X VGND VGND VPWR
+ VPWR _21609_/X sky130_fd_sc_hd__mux4_1
X_28165_ _28165_/A VGND VGND VPWR VPWR _34415_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25377_ _33160_/Q _23453_/X _25395_/S VGND VGND VPWR VPWR _25378_/A sky130_fd_sc_hd__mux2_1
X_22589_ _22373_/X _22587_/X _22588_/X _22377_/X VGND VGND VPWR VPWR _22589_/X sky130_fd_sc_hd__a22o_1
X_27116_ _33968_/Q _27115_/X _27125_/S VGND VGND VPWR VPWR _27117_/A sky130_fd_sc_hd__mux2_1
X_24328_ _24328_/A VGND VGND VPWR VPWR _32695_/D sky130_fd_sc_hd__clkbuf_1
X_28096_ _34383_/Q _27211_/X _28100_/S VGND VGND VPWR VPWR _28097_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27047_ input45/X VGND VGND VPWR VPWR _27047_/X sky130_fd_sc_hd__clkbuf_4
X_24259_ _24259_/A VGND VGND VPWR VPWR _32662_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18820_ _34658_/Q _34594_/Q _34530_/Q _34466_/Q _18533_/X _18534_/X VGND VGND VPWR
+ VPWR _18820_/X sky130_fd_sc_hd__mux4_1
XTAP_6130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28998_ _34809_/Q _27143_/X _29006_/S VGND VGND VPWR VPWR _28999_/A sky130_fd_sc_hd__mux2_1
XFILLER_136_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18751_ _18747_/X _18748_/X _18749_/X _18750_/X VGND VGND VPWR VPWR _18751_/X sky130_fd_sc_hd__a22o_1
X_27949_ _27801_/X _34313_/Q _27965_/S VGND VGND VPWR VPWR _27950_/A sky130_fd_sc_hd__mux2_1
XTAP_6185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17702_ _17420_/X _17698_/X _17701_/X _17424_/X VGND VGND VPWR VPWR _17702_/X sky130_fd_sc_hd__a22o_1
XFILLER_188_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_248_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18682_ _18391_/X _18680_/X _18681_/X _18401_/X VGND VGND VPWR VPWR _18682_/X sky130_fd_sc_hd__a22o_1
XTAP_5484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30960_ _35709_/Q input33/X _30960_/S VGND VGND VPWR VPWR _30961_/A sky130_fd_sc_hd__mux2_1
XTAP_5495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29619_ _35073_/Q _29463_/X _29631_/S VGND VGND VPWR VPWR _29620_/A sky130_fd_sc_hd__mux2_1
XTAP_4783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17633_ _17986_/A VGND VGND VPWR VPWR _17633_/X sky130_fd_sc_hd__buf_6
XFILLER_64_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30891_ _35676_/Q input61/X _30897_/S VGND VGND VPWR VPWR _30892_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32630_ _36023_/CLK _32630_/D VGND VGND VPWR VPWR _32630_/Q sky130_fd_sc_hd__dfxtp_1
X_17564_ _17558_/X _17563_/X _17485_/X VGND VGND VPWR VPWR _17588_/A sky130_fd_sc_hd__o21ba_1
XFILLER_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19303_ _20164_/A VGND VGND VPWR VPWR _19303_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_225_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16515_ _16292_/X _16513_/X _16514_/X _16295_/X VGND VGND VPWR VPWR _16515_/X sky130_fd_sc_hd__a22o_1
XFILLER_210_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32561_ _35953_/CLK _32561_/D VGND VGND VPWR VPWR _32561_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17495_ _17489_/X _17492_/X _17493_/X _17494_/X VGND VGND VPWR VPWR _17520_/B sky130_fd_sc_hd__o211a_1
XFILLER_204_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34300_ _36154_/CLK _34300_/D VGND VGND VPWR VPWR _34300_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31512_ _27779_/X _35970_/Q _31522_/S VGND VGND VPWR VPWR _31513_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19234_ _18945_/X _19232_/X _19233_/X _18948_/X VGND VGND VPWR VPWR _19234_/X sky130_fd_sc_hd__a22o_1
X_35280_ _35729_/CLK _35280_/D VGND VGND VPWR VPWR _35280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16446_ _16441_/X _16444_/X _16445_/X VGND VGND VPWR VPWR _16461_/C sky130_fd_sc_hd__o21ba_1
XFILLER_220_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32492_ _35883_/CLK _32492_/D VGND VGND VPWR VPWR _32492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_1330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34231_ _36150_/CLK _34231_/D VGND VGND VPWR VPWR _34231_/Q sky130_fd_sc_hd__dfxtp_1
X_16377_ _34654_/Q _34590_/Q _34526_/Q _34462_/Q _16233_/X _16234_/X VGND VGND VPWR
+ VPWR _16377_/X sky130_fd_sc_hd__mux4_1
X_31443_ _27677_/X _35937_/Q _31459_/S VGND VGND VPWR VPWR _31444_/A sky130_fd_sc_hd__mux2_1
X_19165_ _19161_/X _19164_/X _19087_/X _19088_/X VGND VGND VPWR VPWR _19182_/B sky130_fd_sc_hd__o211a_1
XFILLER_9_962 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18116_ _35472_/Q _35408_/Q _35344_/Q _35280_/Q _17960_/X _17961_/X VGND VGND VPWR
+ VPWR _18116_/X sky130_fd_sc_hd__mux4_1
XFILLER_129_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31374_ _31374_/A VGND VGND VPWR VPWR _35904_/D sky130_fd_sc_hd__clkbuf_1
X_34162_ _35635_/CLK _34162_/D VGND VGND VPWR VPWR _34162_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19096_ _33066_/Q _32042_/Q _35818_/Q _35754_/Q _19025_/X _19026_/X VGND VGND VPWR
+ VPWR _19096_/X sky130_fd_sc_hd__mux4_1
XFILLER_184_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33113_ _34135_/CLK _33113_/D VGND VGND VPWR VPWR _33113_/Q sky130_fd_sc_hd__dfxtp_1
X_30325_ _35408_/Q _29509_/X _30327_/S VGND VGND VPWR VPWR _30326_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18047_ _33166_/Q _36046_/Q _33038_/Q _32974_/Q _17768_/X _17769_/X VGND VGND VPWR
+ VPWR _18047_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34093_ _34093_/CLK _34093_/D VGND VGND VPWR VPWR _34093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33044_ _36052_/CLK _33044_/D VGND VGND VPWR VPWR _33044_/Q sky130_fd_sc_hd__dfxtp_1
X_30256_ _35375_/Q _29407_/X _30264_/S VGND VGND VPWR VPWR _30257_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_1115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30187_ _30187_/A VGND VGND VPWR VPWR _35342_/D sky130_fd_sc_hd__clkbuf_1
X_19998_ _32132_/Q _32324_/Q _32388_/Q _35908_/Q _19933_/X _19721_/X VGND VGND VPWR
+ VPWR _19998_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_1320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18949_ _18945_/X _18946_/X _18947_/X _18948_/X VGND VGND VPWR VPWR _18949_/X sky130_fd_sc_hd__a22o_1
XFILLER_39_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34995_ _35567_/CLK _34995_/D VGND VGND VPWR VPWR _34995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_1326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33946_ _36219_/CLK _33946_/D VGND VGND VPWR VPWR _33946_/Q sky130_fd_sc_hd__dfxtp_1
X_21960_ _21956_/X _21957_/X _21958_/X _21959_/X VGND VGND VPWR VPWR _21960_/X sky130_fd_sc_hd__a22o_1
XFILLER_239_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1066 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20911_ _20907_/X _20910_/X _20704_/X VGND VGND VPWR VPWR _20912_/D sky130_fd_sc_hd__o21ba_1
XFILLER_66_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33877_ _33941_/CLK _33877_/D VGND VGND VPWR VPWR _33877_/Q sky130_fd_sc_hd__dfxtp_1
X_21891_ _21887_/X _21890_/X _21751_/X VGND VGND VPWR VPWR _21901_/C sky130_fd_sc_hd__o21ba_1
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35616_ _35618_/CLK _35616_/D VGND VGND VPWR VPWR _35616_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23630_ _23630_/A VGND VGND VPWR VPWR _32306_/D sky130_fd_sc_hd__clkbuf_1
X_20842_ _20842_/A _20842_/B _20842_/C _20842_/D VGND VGND VPWR VPWR _20843_/A sky130_fd_sc_hd__or4_1
X_32828_ _32895_/CLK _32828_/D VGND VGND VPWR VPWR _32828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23561_ _32275_/Q _23492_/X _23565_/S VGND VGND VPWR VPWR _23562_/A sky130_fd_sc_hd__mux2_1
X_35547_ _35547_/CLK _35547_/D VGND VGND VPWR VPWR _35547_/Q sky130_fd_sc_hd__dfxtp_1
X_20773_ _34904_/Q _34840_/Q _34776_/Q _34712_/Q _20696_/X _20698_/X VGND VGND VPWR
+ VPWR _20773_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_1266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32759_ _32887_/CLK _32759_/D VGND VGND VPWR VPWR _32759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25300_ _25300_/A VGND VGND VPWR VPWR _33123_/D sky130_fd_sc_hd__clkbuf_1
X_22512_ _22512_/A VGND VGND VPWR VPWR _22512_/X sky130_fd_sc_hd__clkbuf_4
X_26280_ _26280_/A VGND VGND VPWR VPWR _33587_/D sky130_fd_sc_hd__clkbuf_1
X_35478_ _35735_/CLK _35478_/D VGND VGND VPWR VPWR _35478_/Q sky130_fd_sc_hd__dfxtp_1
X_23492_ input58/X VGND VGND VPWR VPWR _23492_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_161_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25231_ _25231_/A VGND VGND VPWR VPWR _33091_/D sky130_fd_sc_hd__clkbuf_1
X_22443_ _32136_/Q _32328_/Q _32392_/Q _35912_/Q _22233_/X _22374_/X VGND VGND VPWR
+ VPWR _22443_/X sky130_fd_sc_hd__mux4_1
X_34429_ _36157_/CLK _34429_/D VGND VGND VPWR VPWR _34429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25162_ _25162_/A VGND VGND VPWR VPWR _33058_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22374_ _22374_/A VGND VGND VPWR VPWR _22374_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_164_966 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24113_ _23082_/X _32597_/Q _24113_/S VGND VGND VPWR VPWR _24114_/A sky130_fd_sc_hd__mux2_1
X_21325_ _22535_/A VGND VGND VPWR VPWR _21325_/X sky130_fd_sc_hd__buf_6
XFILLER_202_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25093_ _24939_/X _33027_/Q _25101_/S VGND VGND VPWR VPWR _25094_/A sky130_fd_sc_hd__mux2_1
X_29970_ _29970_/A VGND VGND VPWR VPWR _35239_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28921_ _34773_/Q _27229_/X _28921_/S VGND VGND VPWR VPWR _28922_/A sky130_fd_sc_hd__mux2_1
X_24044_ _24113_/S VGND VGND VPWR VPWR _24063_/S sky130_fd_sc_hd__buf_4
X_21256_ _34662_/Q _34598_/Q _34534_/Q _34470_/Q _21186_/X _21187_/X VGND VGND VPWR
+ VPWR _21256_/X sky130_fd_sc_hd__mux4_1
XFILLER_132_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_47__f_CLK clkbuf_5_23_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_47__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_20207_ _20207_/A VGND VGND VPWR VPWR _20207_/X sky130_fd_sc_hd__buf_4
XFILLER_46_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28852_ _28921_/S VGND VGND VPWR VPWR _28871_/S sky130_fd_sc_hd__buf_4
XFILLER_133_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21187_ _22599_/A VGND VGND VPWR VPWR _21187_/X sky130_fd_sc_hd__buf_4
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27803_ _27803_/A VGND VGND VPWR VPWR _34249_/D sky130_fd_sc_hd__clkbuf_1
X_20138_ _20138_/A VGND VGND VPWR VPWR _20138_/X sky130_fd_sc_hd__buf_2
X_28783_ _28783_/A VGND VGND VPWR VPWR _34708_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25995_ _24868_/X _33452_/Q _26009_/S VGND VGND VPWR VPWR _25996_/A sky130_fd_sc_hd__mux2_1
XTAP_4013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24946_ _24945_/X _32965_/Q _24952_/S VGND VGND VPWR VPWR _24947_/A sky130_fd_sc_hd__mux2_1
X_20069_ _20074_/A VGND VGND VPWR VPWR _20069_/X sky130_fd_sc_hd__clkbuf_4
XTAP_4035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27734_ _27734_/A VGND VGND VPWR VPWR _34227_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27665_ _27664_/X _34205_/Q _27671_/S VGND VGND VPWR VPWR _27666_/A sky130_fd_sc_hd__mux2_1
XFILLER_218_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24877_ input18/X VGND VGND VPWR VPWR _24877_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29404_ input17/X VGND VGND VPWR VPWR _29404_/X sky130_fd_sc_hd__buf_2
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26616_ _24985_/X _33746_/Q _26622_/S VGND VGND VPWR VPWR _26617_/A sky130_fd_sc_hd__mux2_1
X_23828_ _23064_/X _32399_/Q _23832_/S VGND VGND VPWR VPWR _23829_/A sky130_fd_sc_hd__mux2_1
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27596_ _34177_/Q _27168_/X _27608_/S VGND VGND VPWR VPWR _27597_/A sky130_fd_sc_hd__mux2_1
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29335_ _29335_/A VGND VGND VPWR VPWR _34967_/D sky130_fd_sc_hd__clkbuf_1
X_26547_ _24883_/X _33713_/Q _26551_/S VGND VGND VPWR VPWR _26548_/A sky130_fd_sc_hd__mux2_1
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23759_ _22962_/X _32366_/Q _23769_/S VGND VGND VPWR VPWR _23760_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16300_ _17869_/A VGND VGND VPWR VPWR _16300_/X sky130_fd_sc_hd__buf_4
XFILLER_18_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17280_ _17986_/A VGND VGND VPWR VPWR _17280_/X sky130_fd_sc_hd__buf_6
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26478_ _33681_/Q _23484_/X _26478_/S VGND VGND VPWR VPWR _26479_/A sky130_fd_sc_hd__mux2_1
X_29266_ _34936_/Q _27140_/X _29276_/S VGND VGND VPWR VPWR _29267_/A sky130_fd_sc_hd__mux2_1
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_1478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16231_ _16060_/X _16229_/X _16230_/X _16072_/X VGND VGND VPWR VPWR _16231_/X sky130_fd_sc_hd__a22o_1
X_28217_ _27797_/X _34440_/Q _28235_/S VGND VGND VPWR VPWR _28218_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25429_ _25540_/S VGND VGND VPWR VPWR _25448_/S sky130_fd_sc_hd__buf_4
X_29197_ _34903_/Q _27038_/X _29213_/S VGND VGND VPWR VPWR _29198_/A sky130_fd_sc_hd__mux2_1
XFILLER_224_1393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16162_ _16048_/X _16160_/X _16161_/X _16058_/X VGND VGND VPWR VPWR _16162_/X sky130_fd_sc_hd__a22o_1
XFILLER_142_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28148_ _28148_/A VGND VGND VPWR VPWR _34407_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28079_ _34375_/Q _27186_/X _28079_/S VGND VGND VPWR VPWR _28080_/A sky130_fd_sc_hd__mux2_1
X_16093_ _17766_/A VGND VGND VPWR VPWR _16877_/A sky130_fd_sc_hd__buf_8
XFILLER_142_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30110_ _30200_/S VGND VGND VPWR VPWR _30129_/S sky130_fd_sc_hd__buf_6
X_19921_ _19921_/A VGND VGND VPWR VPWR _32449_/D sky130_fd_sc_hd__clkbuf_4
X_31090_ _31090_/A VGND VGND VPWR VPWR _35770_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30041_ _35273_/Q _29488_/X _30057_/S VGND VGND VPWR VPWR _30042_/A sky130_fd_sc_hd__mux2_1
X_19852_ _20205_/A VGND VGND VPWR VPWR _19852_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_155_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_150_CLK clkbuf_6_29__f_CLK/X VGND VGND VPWR VPWR _36181_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_150_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18803_ _20169_/A VGND VGND VPWR VPWR _18803_/X sky130_fd_sc_hd__buf_4
XFILLER_1_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19783_ _33918_/Q _33854_/Q _33790_/Q _36094_/Q _19677_/X _19678_/X VGND VGND VPWR
+ VPWR _19783_/X sky130_fd_sc_hd__mux4_1
X_16995_ _32880_/Q _32816_/Q _32752_/Q _32688_/Q _16993_/X _16994_/X VGND VGND VPWR
+ VPWR _16995_/X sky130_fd_sc_hd__mux4_1
XFILLER_62_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33800_ _36105_/CLK _33800_/D VGND VGND VPWR VPWR _33800_/Q sky130_fd_sc_hd__dfxtp_1
X_18734_ _20146_/A VGND VGND VPWR VPWR _18734_/X sky130_fd_sc_hd__buf_2
X_34780_ _36242_/CLK _34780_/D VGND VGND VPWR VPWR _34780_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31992_ _34405_/CLK _31992_/D VGND VGND VPWR VPWR _31992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33731_ _35843_/CLK _33731_/D VGND VGND VPWR VPWR _33731_/Q sky130_fd_sc_hd__dfxtp_1
X_18665_ _20215_/A VGND VGND VPWR VPWR _18665_/X sky130_fd_sc_hd__clkbuf_4
X_30943_ _30943_/A VGND VGND VPWR VPWR _35700_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_209_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17616_ _34433_/Q _36161_/Q _34305_/Q _34241_/Q _17582_/X _17583_/X VGND VGND VPWR
+ VPWR _17616_/X sky130_fd_sc_hd__mux4_1
X_33662_ _35456_/CLK _33662_/D VGND VGND VPWR VPWR _33662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30874_ _30874_/A VGND VGND VPWR VPWR _35668_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18596_ _18592_/X _18593_/X _18594_/X _18595_/X VGND VGND VPWR VPWR _18596_/X sky130_fd_sc_hd__a22o_1
XTAP_3890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35401_ _35466_/CLK _35401_/D VGND VGND VPWR VPWR _35401_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32613_ _35943_/CLK _32613_/D VGND VGND VPWR VPWR _32613_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17547_ _34943_/Q _34879_/Q _34815_/Q _34751_/Q _17513_/X _17514_/X VGND VGND VPWR
+ VPWR _17547_/X sky130_fd_sc_hd__mux4_1
XFILLER_211_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33593_ _33913_/CLK _33593_/D VGND VGND VPWR VPWR _33593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35332_ _35843_/CLK _35332_/D VGND VGND VPWR VPWR _35332_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32544_ _35938_/CLK _32544_/D VGND VGND VPWR VPWR _32544_/Q sky130_fd_sc_hd__dfxtp_1
X_17478_ _34174_/Q _34110_/Q _34046_/Q _33982_/Q _17446_/X _17447_/X VGND VGND VPWR
+ VPWR _17478_/X sky130_fd_sc_hd__mux4_1
XFILLER_149_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19217_ _34158_/Q _34094_/Q _34030_/Q _33966_/Q _19040_/X _19041_/X VGND VGND VPWR
+ VPWR _19217_/X sky130_fd_sc_hd__mux4_1
X_35263_ _35839_/CLK _35263_/D VGND VGND VPWR VPWR _35263_/Q sky130_fd_sc_hd__dfxtp_1
X_16429_ _33120_/Q _36000_/Q _32992_/Q _32928_/Q _16356_/X _16357_/X VGND VGND VPWR
+ VPWR _16429_/X sky130_fd_sc_hd__mux4_1
XFILLER_242_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32475_ _35994_/CLK _32475_/D VGND VGND VPWR VPWR _32475_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34214_ _34405_/CLK _34214_/D VGND VGND VPWR VPWR _34214_/Q sky130_fd_sc_hd__dfxtp_1
X_31426_ _27652_/X _35929_/Q _31438_/S VGND VGND VPWR VPWR _31427_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19148_ _20207_/A VGND VGND VPWR VPWR _19148_/X sky130_fd_sc_hd__clkbuf_4
X_35194_ _35194_/CLK _35194_/D VGND VGND VPWR VPWR _35194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34145_ _34593_/CLK _34145_/D VGND VGND VPWR VPWR _34145_/Q sky130_fd_sc_hd__dfxtp_1
X_19079_ _20138_/A VGND VGND VPWR VPWR _19079_/X sky130_fd_sc_hd__buf_2
X_31357_ _31357_/A VGND VGND VPWR VPWR _35896_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_246_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21110_ _32866_/Q _32802_/Q _32738_/Q _32674_/Q _20887_/X _20888_/X VGND VGND VPWR
+ VPWR _21110_/X sky130_fd_sc_hd__mux4_1
X_30308_ _30335_/S VGND VGND VPWR VPWR _30327_/S sky130_fd_sc_hd__buf_4
XFILLER_246_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34076_ _36211_/CLK _34076_/D VGND VGND VPWR VPWR _34076_/Q sky130_fd_sc_hd__dfxtp_1
X_22090_ _32126_/Q _32318_/Q _32382_/Q _35902_/Q _21880_/X _22021_/X VGND VGND VPWR
+ VPWR _22090_/X sky130_fd_sc_hd__mux4_1
X_31288_ _31288_/A VGND VGND VPWR VPWR _35863_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_1415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33027_ _35779_/CLK _33027_/D VGND VGND VPWR VPWR _33027_/Q sky130_fd_sc_hd__dfxtp_1
X_21041_ _20892_/X _21037_/X _21040_/X _20895_/X VGND VGND VPWR VPWR _21041_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_141_CLK clkbuf_6_28__f_CLK/X VGND VGND VPWR VPWR _35929_/CLK sky130_fd_sc_hd__clkbuf_16
X_30239_ _35367_/Q _29382_/X _30243_/S VGND VGND VPWR VPWR _30240_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24800_ _24995_/S VGND VGND VPWR VPWR _24828_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_75_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25780_ _25780_/A VGND VGND VPWR VPWR _33350_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22992_ _22992_/A VGND VGND VPWR VPWR _32055_/D sky130_fd_sc_hd__clkbuf_1
X_34978_ _35177_/CLK _34978_/D VGND VGND VPWR VPWR _34978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24731_ _24731_/A VGND VGND VPWR VPWR _32886_/D sky130_fd_sc_hd__clkbuf_1
X_33929_ _36104_/CLK _33929_/D VGND VGND VPWR VPWR _33929_/Q sky130_fd_sc_hd__dfxtp_1
X_21943_ _33146_/Q _36026_/Q _33018_/Q _32954_/Q _21662_/X _21663_/X VGND VGND VPWR
+ VPWR _21943_/X sky130_fd_sc_hd__mux4_1
XFILLER_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27450_ _34108_/Q _27152_/X _27452_/S VGND VGND VPWR VPWR _27451_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24662_ _24794_/S VGND VGND VPWR VPWR _24681_/S sky130_fd_sc_hd__clkbuf_8
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21874_ _21806_/X _21872_/X _21873_/X _21809_/X VGND VGND VPWR VPWR _21874_/X sky130_fd_sc_hd__a22o_1
XFILLER_54_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26401_ _33644_/Q _23299_/X _26415_/S VGND VGND VPWR VPWR _26402_/A sky130_fd_sc_hd__mux2_1
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23613_ _22949_/X _32298_/Q _23631_/S VGND VGND VPWR VPWR _23614_/A sky130_fd_sc_hd__mux2_1
X_27381_ _34075_/Q _27050_/X _27389_/S VGND VGND VPWR VPWR _27382_/A sky130_fd_sc_hd__mux2_1
X_20825_ _20820_/X _20824_/X _20644_/X _20646_/X VGND VGND VPWR VPWR _20842_/B sky130_fd_sc_hd__o211a_1
XFILLER_39_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24593_ _22984_/X _32821_/Q _24609_/S VGND VGND VPWR VPWR _24594_/A sky130_fd_sc_hd__mux2_1
XFILLER_247_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26332_ _24967_/X _33612_/Q _26342_/S VGND VGND VPWR VPWR _26333_/A sky130_fd_sc_hd__mux2_1
X_29120_ _34867_/Q _27124_/X _29120_/S VGND VGND VPWR VPWR _29121_/A sky130_fd_sc_hd__mux2_1
XFILLER_208_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23544_ _23544_/A VGND VGND VPWR VPWR _32266_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20756_ _32088_/Q _32280_/Q _32344_/Q _35864_/Q _20632_/X _22467_/A VGND VGND VPWR
+ VPWR _20756_/X sky130_fd_sc_hd__mux4_1
XFILLER_126_1044 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29051_ _29051_/A VGND VGND VPWR VPWR _34834_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26263_ _24865_/X _33579_/Q _26279_/S VGND VGND VPWR VPWR _26264_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23475_ input52/X VGND VGND VPWR VPWR _23475_/X sky130_fd_sc_hd__buf_4
X_20687_ _22371_/A VGND VGND VPWR VPWR _21756_/A sky130_fd_sc_hd__buf_8
X_28002_ _34338_/Q _27072_/X _28016_/S VGND VGND VPWR VPWR _28003_/A sky130_fd_sc_hd__mux2_1
X_25214_ _25214_/A VGND VGND VPWR VPWR _33083_/D sky130_fd_sc_hd__clkbuf_1
X_22426_ _22111_/X _22424_/X _22425_/X _22116_/X VGND VGND VPWR VPWR _22426_/X sky130_fd_sc_hd__a22o_1
XFILLER_196_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26194_ _26194_/A VGND VGND VPWR VPWR _33546_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25145_ _25145_/A VGND VGND VPWR VPWR _33050_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22357_ _22357_/A VGND VGND VPWR VPWR _36229_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_380_CLK clkbuf_6_42__f_CLK/X VGND VGND VPWR VPWR _33661_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_124_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21308_ _32616_/Q _32552_/Q _32488_/Q _35944_/Q _21170_/X _21307_/X VGND VGND VPWR
+ VPWR _21308_/X sky130_fd_sc_hd__mux4_1
X_29953_ _29953_/A VGND VGND VPWR VPWR _35231_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25076_ _24914_/X _33019_/Q _25080_/S VGND VGND VPWR VPWR _25077_/A sky130_fd_sc_hd__mux2_1
X_22288_ _33668_/Q _33604_/Q _33540_/Q _33476_/Q _22153_/X _22154_/X VGND VGND VPWR
+ VPWR _22288_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28904_ _28904_/A VGND VGND VPWR VPWR _34764_/D sky130_fd_sc_hd__clkbuf_1
X_24027_ _24027_/A VGND VGND VPWR VPWR _32555_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_132_CLK clkbuf_6_23__f_CLK/X VGND VGND VPWR VPWR _34903_/CLK sky130_fd_sc_hd__clkbuf_16
X_21239_ _32102_/Q _32294_/Q _32358_/Q _35878_/Q _21174_/X _20962_/X VGND VGND VPWR
+ VPWR _21239_/X sky130_fd_sc_hd__mux4_1
X_29884_ _29884_/A VGND VGND VPWR VPWR _35198_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28835_ _28835_/A VGND VGND VPWR VPWR _34731_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28766_ _34700_/Q _27202_/X _28776_/S VGND VGND VPWR VPWR _28767_/A sky130_fd_sc_hd__mux2_1
X_16780_ _16773_/X _16778_/X _16779_/X VGND VGND VPWR VPWR _16814_/A sky130_fd_sc_hd__o21ba_1
XFILLER_19_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25978_ _24843_/X _33444_/Q _25988_/S VGND VGND VPWR VPWR _25979_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_1102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27717_ input17/X VGND VGND VPWR VPWR _27717_/X sky130_fd_sc_hd__buf_2
XTAP_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24929_ _24929_/A VGND VGND VPWR VPWR _32959_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28697_ _34667_/Q _27100_/X _28713_/S VGND VGND VPWR VPWR _28698_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_1368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18450_ _20169_/A VGND VGND VPWR VPWR _18450_/X sky130_fd_sc_hd__clkbuf_8
XTAP_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27648_ _27648_/A VGND VGND VPWR VPWR _34199_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17401_ _17158_/X _17399_/X _17400_/X _17163_/X VGND VGND VPWR VPWR _17401_/X sky130_fd_sc_hd__a22o_1
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18381_ _34646_/Q _34582_/Q _34518_/Q _34454_/Q _18379_/X _18380_/X VGND VGND VPWR
+ VPWR _18381_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_199_CLK clkbuf_6_49__f_CLK/X VGND VGND VPWR VPWR _35723_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27579_ _34169_/Q _27143_/X _27587_/S VGND VGND VPWR VPWR _27580_/A sky130_fd_sc_hd__mux2_1
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29318_ _34961_/Q _27217_/X _29318_/S VGND VGND VPWR VPWR _29319_/A sky130_fd_sc_hd__mux2_1
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17332_ _17328_/X _17331_/X _17165_/X VGND VGND VPWR VPWR _17333_/D sky130_fd_sc_hd__o21ba_1
X_30590_ _30590_/A VGND VGND VPWR VPWR _35533_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29249_ _34928_/Q _27115_/X _29255_/S VGND VGND VPWR VPWR _29250_/A sky130_fd_sc_hd__mux2_1
X_17263_ _34423_/Q _36151_/Q _34295_/Q _34231_/Q _17229_/X _17230_/X VGND VGND VPWR
+ VPWR _17263_/X sky130_fd_sc_hd__mux4_1
XFILLER_186_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19002_ _33384_/Q _33320_/Q _33256_/Q _33192_/Q _18721_/X _18722_/X VGND VGND VPWR
+ VPWR _19002_/X sky130_fd_sc_hd__mux4_1
X_16214_ _33882_/Q _33818_/Q _33754_/Q _36058_/Q _16112_/X _16113_/X VGND VGND VPWR
+ VPWR _16214_/X sky130_fd_sc_hd__mux4_1
X_32260_ _34693_/CLK _32260_/D VGND VGND VPWR VPWR _32260_/Q sky130_fd_sc_hd__dfxtp_1
X_17194_ _34933_/Q _34869_/Q _34805_/Q _34741_/Q _17160_/X _17161_/X VGND VGND VPWR
+ VPWR _17194_/X sky130_fd_sc_hd__mux4_1
XFILLER_128_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16145_ _17862_/A VGND VGND VPWR VPWR _16145_/X sky130_fd_sc_hd__buf_4
X_31211_ _31211_/A VGND VGND VPWR VPWR _35827_/D sky130_fd_sc_hd__clkbuf_1
X_32191_ _35684_/CLK _32191_/D VGND VGND VPWR VPWR _32191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_914 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_371_CLK clkbuf_6_43__f_CLK/X VGND VGND VPWR VPWR _34685_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_155_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16076_ _16059_/X _16073_/X _16075_/X VGND VGND VPWR VPWR _16106_/C sky130_fd_sc_hd__o21ba_1
X_31142_ _31142_/A VGND VGND VPWR VPWR _35795_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19904_ _35713_/Q _32223_/Q _35585_/Q _35521_/Q _19617_/X _19618_/X VGND VGND VPWR
+ VPWR _19904_/X sky130_fd_sc_hd__mux4_1
X_31073_ _31073_/A VGND VGND VPWR VPWR _35762_/D sky130_fd_sc_hd__clkbuf_1
X_35950_ _35951_/CLK _35950_/D VGND VGND VPWR VPWR _35950_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_123_CLK clkbuf_6_21__f_CLK/X VGND VGND VPWR VPWR _36235_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_233_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_30__f_CLK clkbuf_5_15_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_30__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_123_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34901_ _36181_/CLK _34901_/D VGND VGND VPWR VPWR _34901_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_233_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30024_ _35265_/Q _29463_/X _30036_/S VGND VGND VPWR VPWR _30025_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19835_ _19831_/X _19834_/X _19793_/X _19794_/X VGND VGND VPWR VPWR _19850_/B sky130_fd_sc_hd__o211a_1
XFILLER_111_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35881_ _35947_/CLK _35881_/D VGND VGND VPWR VPWR _35881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34832_ _34897_/CLK _34832_/D VGND VGND VPWR VPWR _34832_/Q sky130_fd_sc_hd__dfxtp_1
X_19766_ _19656_/X _19764_/X _19765_/X _19659_/X VGND VGND VPWR VPWR _19766_/X sky130_fd_sc_hd__a22o_1
X_16978_ _16805_/X _16976_/X _16977_/X _16810_/X VGND VGND VPWR VPWR _16978_/X sky130_fd_sc_hd__a22o_1
XFILLER_231_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput4 DW[12] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__buf_6
XFILLER_237_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18717_ _18717_/A VGND VGND VPWR VPWR _32415_/D sky130_fd_sc_hd__clkbuf_1
X_34763_ _34957_/CLK _34763_/D VGND VGND VPWR VPWR _34763_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_225_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31975_ _34790_/CLK _31975_/D VGND VGND VPWR VPWR _31975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19697_ _35195_/Q _35131_/Q _35067_/Q _32251_/Q _19663_/X _19664_/X VGND VGND VPWR
+ VPWR _19697_/X sky130_fd_sc_hd__mux4_1
XFILLER_188_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33714_ _35633_/CLK _33714_/D VGND VGND VPWR VPWR _33714_/Q sky130_fd_sc_hd__dfxtp_1
X_18648_ _18440_/X _18646_/X _18647_/X _18445_/X VGND VGND VPWR VPWR _18648_/X sky130_fd_sc_hd__a22o_1
X_30926_ _30926_/A VGND VGND VPWR VPWR _35692_/D sky130_fd_sc_hd__clkbuf_1
X_34694_ _34694_/CLK _34694_/D VGND VGND VPWR VPWR _34694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33645_ _33902_/CLK _33645_/D VGND VGND VPWR VPWR _33645_/Q sky130_fd_sc_hd__dfxtp_1
X_30857_ _35660_/Q input50/X _30867_/S VGND VGND VPWR VPWR _30858_/A sky130_fd_sc_hd__mux2_1
X_18579_ _33372_/Q _33308_/Q _33244_/Q _33180_/Q _18302_/X _18303_/X VGND VGND VPWR
+ VPWR _18579_/X sky130_fd_sc_hd__mux4_1
XFILLER_178_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20610_ _20663_/A VGND VGND VPWR VPWR _22561_/A sky130_fd_sc_hd__buf_12
XFILLER_221_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33576_ _35622_/CLK _33576_/D VGND VGND VPWR VPWR _33576_/Q sky130_fd_sc_hd__dfxtp_1
X_21590_ _33136_/Q _36016_/Q _33008_/Q _32944_/Q _21309_/X _21310_/X VGND VGND VPWR
+ VPWR _21590_/X sky130_fd_sc_hd__mux4_1
X_30788_ _35627_/Q input14/X _30804_/S VGND VGND VPWR VPWR _30789_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_1247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35315_ _35764_/CLK _35315_/D VGND VGND VPWR VPWR _35315_/Q sky130_fd_sc_hd__dfxtp_1
X_20541_ _35220_/Q _35156_/Q _35092_/Q _32276_/Q _18392_/X _18394_/X VGND VGND VPWR
+ VPWR _20541_/X sky130_fd_sc_hd__mux4_1
X_32527_ _35983_/CLK _32527_/D VGND VGND VPWR VPWR _32527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23260_ _23260_/A VGND VGND VPWR VPWR _32159_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35246_ _35438_/CLK _35246_/D VGND VGND VPWR VPWR _35246_/Q sky130_fd_sc_hd__dfxtp_1
X_20472_ _20468_/X _20471_/X _20146_/A _20147_/A VGND VGND VPWR VPWR _20487_/B sky130_fd_sc_hd__o211a_1
X_32458_ _36077_/CLK _32458_/D VGND VGND VPWR VPWR _32458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22211_ _21956_/X _22209_/X _22210_/X _21959_/X VGND VGND VPWR VPWR _22211_/X sky130_fd_sc_hd__a22o_1
XFILLER_145_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31409_ _31409_/A VGND VGND VPWR VPWR _35921_/D sky130_fd_sc_hd__clkbuf_1
X_23191_ _23191_/A VGND VGND VPWR VPWR _32133_/D sky130_fd_sc_hd__clkbuf_1
X_35177_ _35177_/CLK _35177_/D VGND VGND VPWR VPWR _35177_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_362_CLK clkbuf_6_44__f_CLK/X VGND VGND VPWR VPWR _35835_/CLK sky130_fd_sc_hd__clkbuf_16
X_32389_ _32901_/CLK _32389_/D VGND VGND VPWR VPWR _32389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34128_ _34192_/CLK _34128_/D VGND VGND VPWR VPWR _34128_/Q sky130_fd_sc_hd__dfxtp_1
X_22142_ _22138_/X _22141_/X _22104_/X VGND VGND VPWR VPWR _22150_/C sky130_fd_sc_hd__o21ba_1
XFILLER_10_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34059_ _34187_/CLK _34059_/D VGND VGND VPWR VPWR _34059_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_114_CLK clkbuf_6_20__f_CLK/X VGND VGND VPWR VPWR _35609_/CLK sky130_fd_sc_hd__clkbuf_16
X_26950_ _33902_/Q _23305_/X _26960_/S VGND VGND VPWR VPWR _26951_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22073_ _21758_/X _22071_/X _22072_/X _21763_/X VGND VGND VPWR VPWR _22073_/X sky130_fd_sc_hd__a22o_1
XTAP_6729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25901_ _25901_/A VGND VGND VPWR VPWR _33407_/D sky130_fd_sc_hd__clkbuf_1
X_21024_ _33888_/Q _33824_/Q _33760_/Q _36064_/Q _20918_/X _20919_/X VGND VGND VPWR
+ VPWR _21024_/X sky130_fd_sc_hd__mux4_1
XFILLER_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26881_ _26881_/A VGND VGND VPWR VPWR _33869_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28620_ _28620_/A VGND VGND VPWR VPWR _34631_/D sky130_fd_sc_hd__clkbuf_1
X_25832_ _24827_/X _33375_/Q _25832_/S VGND VGND VPWR VPWR _25833_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28551_ _28551_/A VGND VGND VPWR VPWR _34598_/D sky130_fd_sc_hd__clkbuf_1
X_25763_ _24923_/X _33342_/Q _25781_/S VGND VGND VPWR VPWR _25764_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22975_ _22974_/X _32050_/Q _22978_/S VGND VGND VPWR VPWR _22976_/A sky130_fd_sc_hd__mux2_1
X_27502_ _34133_/Q _27229_/X _27502_/S VGND VGND VPWR VPWR _27503_/A sky130_fd_sc_hd__mux2_1
X_24714_ _24714_/A VGND VGND VPWR VPWR _32878_/D sky130_fd_sc_hd__clkbuf_1
X_21926_ _34681_/Q _34617_/Q _34553_/Q _34489_/Q _21892_/X _21893_/X VGND VGND VPWR
+ VPWR _21926_/X sky130_fd_sc_hd__mux4_1
X_28482_ _27791_/X _34566_/Q _28484_/S VGND VGND VPWR VPWR _28483_/A sky130_fd_sc_hd__mux2_1
X_25694_ _25694_/A VGND VGND VPWR VPWR _33309_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24645_ _23061_/X _32846_/Q _24651_/S VGND VGND VPWR VPWR _24646_/A sky130_fd_sc_hd__mux2_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27433_ _27502_/S VGND VGND VPWR VPWR _27452_/S sky130_fd_sc_hd__buf_4
XFILLER_188_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21857_ _33079_/Q _32055_/Q _35831_/Q _35767_/Q _21678_/X _21679_/X VGND VGND VPWR
+ VPWR _21857_/X sky130_fd_sc_hd__mux4_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20808_ _20808_/A _20808_/B _20808_/C _20808_/D VGND VGND VPWR VPWR _20809_/A sky130_fd_sc_hd__or4_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27364_ _27364_/A VGND VGND VPWR VPWR _34067_/D sky130_fd_sc_hd__clkbuf_1
X_24576_ _22959_/X _32813_/Q _24588_/S VGND VGND VPWR VPWR _24577_/A sky130_fd_sc_hd__mux2_1
X_21788_ _21603_/X _21786_/X _21787_/X _21606_/X VGND VGND VPWR VPWR _21788_/X sky130_fd_sc_hd__a22o_1
XFILLER_93_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29103_ _29103_/A VGND VGND VPWR VPWR _34858_/D sky130_fd_sc_hd__clkbuf_1
X_26315_ _24942_/X _33604_/Q _26321_/S VGND VGND VPWR VPWR _26316_/A sky130_fd_sc_hd__mux2_1
X_23527_ _23527_/A VGND VGND VPWR VPWR _32258_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20739_ _20739_/A VGND VGND VPWR VPWR _36183_/D sky130_fd_sc_hd__clkbuf_2
X_27295_ _27295_/A VGND VGND VPWR VPWR _34034_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29034_ _34826_/Q _27196_/X _29048_/S VGND VGND VPWR VPWR _29035_/A sky130_fd_sc_hd__mux2_1
XFILLER_221_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26246_ _24840_/X _33571_/Q _26258_/S VGND VGND VPWR VPWR _26247_/A sky130_fd_sc_hd__mux2_1
X_23458_ _32231_/Q _23387_/X _23515_/S VGND VGND VPWR VPWR _23459_/A sky130_fd_sc_hd__mux2_1
XFILLER_221_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22409_ _22365_/X _22407_/X _22408_/X _22371_/X VGND VGND VPWR VPWR _22409_/X sky130_fd_sc_hd__a22o_1
X_26177_ _26177_/A VGND VGND VPWR VPWR _33538_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23389_ _32208_/Q _23387_/X _23418_/S VGND VGND VPWR VPWR _23390_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_1134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_353_CLK clkbuf_6_46__f_CLK/X VGND VGND VPWR VPWR _35451_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_137_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25128_ _24991_/X _33044_/Q _25130_/S VGND VGND VPWR VPWR _25129_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29936_ _35223_/Q _29333_/X _29952_/S VGND VGND VPWR VPWR _29937_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_105_CLK clkbuf_leaf_99_CLK/A VGND VGND VPWR VPWR _35547_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_151_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17950_ _32651_/Q _32587_/Q _32523_/Q _35979_/Q _17629_/X _17766_/X VGND VGND VPWR
+ VPWR _17950_/X sky130_fd_sc_hd__mux4_1
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25059_ _24889_/X _33011_/Q _25059_/S VGND VGND VPWR VPWR _25060_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16901_ _17960_/A VGND VGND VPWR VPWR _16901_/X sky130_fd_sc_hd__buf_4
XFILLER_78_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17881_ _17877_/X _17880_/X _17838_/X VGND VGND VPWR VPWR _17903_/A sky130_fd_sc_hd__o21ba_2
X_29867_ _29867_/A VGND VGND VPWR VPWR _35190_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19620_ _35641_/Q _35001_/Q _34361_/Q _33721_/Q _19444_/X _19445_/X VGND VGND VPWR
+ VPWR _19620_/X sky130_fd_sc_hd__mux4_1
X_16832_ _16645_/X _16830_/X _16831_/X _16648_/X VGND VGND VPWR VPWR _16832_/X sky130_fd_sc_hd__a22o_1
X_28818_ _28818_/A VGND VGND VPWR VPWR _34723_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29798_ _29930_/S VGND VGND VPWR VPWR _29817_/S sky130_fd_sc_hd__buf_6
XFILLER_8_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19551_ _35703_/Q _32212_/Q _35575_/Q _35511_/Q _19264_/X _19265_/X VGND VGND VPWR
+ VPWR _19551_/X sky130_fd_sc_hd__mux4_1
XFILLER_207_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28749_ _34692_/Q _27177_/X _28755_/S VGND VGND VPWR VPWR _28750_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16763_ _35177_/Q _35113_/Q _35049_/Q _32169_/Q _16657_/X _16658_/X VGND VGND VPWR
+ VPWR _16763_/X sky130_fd_sc_hd__mux4_1
XFILLER_247_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18502_ _35161_/Q _35097_/Q _35033_/Q _32153_/Q _18383_/X _18385_/X VGND VGND VPWR
+ VPWR _18502_/X sky130_fd_sc_hd__mux4_1
XFILLER_207_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_975 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31760_ _31760_/A VGND VGND VPWR VPWR _36087_/D sky130_fd_sc_hd__clkbuf_1
X_19482_ _19478_/X _19481_/X _19440_/X _19441_/X VGND VGND VPWR VPWR _19497_/B sky130_fd_sc_hd__o211a_1
XFILLER_185_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16694_ _34919_/Q _34855_/Q _34791_/Q _34727_/Q _16454_/X _16455_/X VGND VGND VPWR
+ VPWR _16694_/X sky130_fd_sc_hd__mux4_1
XFILLER_34_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18433_ _18378_/X _18431_/X _18432_/X _18388_/X VGND VGND VPWR VPWR _18433_/X sky130_fd_sc_hd__a22o_1
X_30711_ _35591_/Q _29481_/X _30711_/S VGND VGND VPWR VPWR _30712_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31691_ _31691_/A VGND VGND VPWR VPWR _36054_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33430_ _35861_/CLK _33430_/D VGND VGND VPWR VPWR _33430_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18364_ _20151_/A VGND VGND VPWR VPWR _18364_/X sky130_fd_sc_hd__buf_4
XFILLER_203_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30642_ _35558_/Q _29379_/X _30648_/S VGND VGND VPWR VPWR _30643_/A sky130_fd_sc_hd__mux2_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17315_ _17067_/X _17313_/X _17314_/X _17071_/X VGND VGND VPWR VPWR _17315_/X sky130_fd_sc_hd__a22o_1
X_33361_ _36106_/CLK _33361_/D VGND VGND VPWR VPWR _33361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18295_ _20100_/A VGND VGND VPWR VPWR _18295_/X sky130_fd_sc_hd__clkbuf_4
X_30573_ _30573_/A VGND VGND VPWR VPWR _35525_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_222_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35100_ _36219_/CLK _35100_/D VGND VGND VPWR VPWR _35100_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32312_ _32889_/CLK _32312_/D VGND VGND VPWR VPWR _32312_/Q sky130_fd_sc_hd__dfxtp_1
X_36080_ _36080_/CLK _36080_/D VGND VGND VPWR VPWR _36080_/Q sky130_fd_sc_hd__dfxtp_1
X_17246_ _17059_/X _17244_/X _17245_/X _17065_/X VGND VGND VPWR VPWR _17246_/X sky130_fd_sc_hd__a22o_1
X_33292_ _33425_/CLK _33292_/D VGND VGND VPWR VPWR _33292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35031_ _35799_/CLK _35031_/D VGND VGND VPWR VPWR _35031_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32243_ _35731_/CLK _32243_/D VGND VGND VPWR VPWR _32243_/Q sky130_fd_sc_hd__dfxtp_1
X_17177_ _33141_/Q _36021_/Q _33013_/Q _32949_/Q _17062_/X _17063_/X VGND VGND VPWR
+ VPWR _17177_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_344_CLK clkbuf_6_45__f_CLK/X VGND VGND VPWR VPWR _35964_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_116_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16128_ _33047_/Q _32023_/Q _35799_/Q _35735_/Q _16067_/X _16069_/X VGND VGND VPWR
+ VPWR _16128_/X sky130_fd_sc_hd__mux4_1
XFILLER_157_1324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32174_ _36142_/CLK _32174_/D VGND VGND VPWR VPWR _32174_/Q sky130_fd_sc_hd__dfxtp_1
X_31125_ _35787_/Q input49/X _31137_/S VGND VGND VPWR VPWR _31126_/A sky130_fd_sc_hd__mux2_1
X_16059_ _16048_/X _16051_/X _16056_/X _16058_/X VGND VGND VPWR VPWR _16059_/X sky130_fd_sc_hd__a22o_1
XFILLER_88_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35933_ _35998_/CLK _35933_/D VGND VGND VPWR VPWR _35933_/Q sky130_fd_sc_hd__dfxtp_1
X_31056_ _35754_/Q input13/X _31074_/S VGND VGND VPWR VPWR _31057_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19818_ _20171_/A VGND VGND VPWR VPWR _19818_/X sky130_fd_sc_hd__buf_2
X_30007_ _35257_/Q _29438_/X _30015_/S VGND VGND VPWR VPWR _30008_/A sky130_fd_sc_hd__mux2_1
XFILLER_57_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35864_ _35990_/CLK _35864_/D VGND VGND VPWR VPWR _35864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34815_ _34815_/CLK _34815_/D VGND VGND VPWR VPWR _34815_/Q sky130_fd_sc_hd__dfxtp_1
X_19749_ _19499_/X _19745_/X _19748_/X _19504_/X VGND VGND VPWR VPWR _19749_/X sky130_fd_sc_hd__a22o_1
X_35795_ _35859_/CLK _35795_/D VGND VGND VPWR VPWR _35795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22760_ _34194_/Q _34130_/Q _34066_/Q _34002_/Q _20649_/X _20650_/X VGND VGND VPWR
+ VPWR _22760_/X sky130_fd_sc_hd__mux4_1
X_34746_ _36153_/CLK _34746_/D VGND VGND VPWR VPWR _34746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31958_ _34148_/CLK _31958_/D VGND VGND VPWR VPWR _31958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21711_ _35443_/Q _35379_/Q _35315_/Q _35251_/Q _21501_/X _21502_/X VGND VGND VPWR
+ VPWR _21711_/X sky130_fd_sc_hd__mux4_1
XFILLER_213_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30909_ _30909_/A VGND VGND VPWR VPWR _35684_/D sky130_fd_sc_hd__clkbuf_1
X_22691_ _35215_/Q _35151_/Q _35087_/Q _32271_/Q _20692_/X _20694_/X VGND VGND VPWR
+ VPWR _22691_/X sky130_fd_sc_hd__mux4_1
XFILLER_25_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34677_ _35126_/CLK _34677_/D VGND VGND VPWR VPWR _34677_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31889_ _31889_/A VGND VGND VPWR VPWR _36148_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24430_ _22943_/X _32744_/Q _24432_/S VGND VGND VPWR VPWR _24431_/A sky130_fd_sc_hd__mux2_1
XFILLER_244_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33628_ _36211_/CLK _33628_/D VGND VGND VPWR VPWR _33628_/Q sky130_fd_sc_hd__dfxtp_1
X_21642_ _21638_/X _21641_/X _21398_/X VGND VGND VPWR VPWR _21650_/C sky130_fd_sc_hd__o21ba_1
XFILLER_75_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_240_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24361_ _24361_/A VGND VGND VPWR VPWR _32711_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33559_ _35995_/CLK _33559_/D VGND VGND VPWR VPWR _33559_/Q sky130_fd_sc_hd__dfxtp_1
X_21573_ _34671_/Q _34607_/Q _34543_/Q _34479_/Q _21539_/X _21540_/X VGND VGND VPWR
+ VPWR _21573_/X sky130_fd_sc_hd__mux4_1
X_26100_ _24824_/X _33502_/Q _26102_/S VGND VGND VPWR VPWR _26101_/A sky130_fd_sc_hd__mux2_1
X_23312_ _30877_/A _29662_/B VGND VGND VPWR VPWR _23499_/S sky130_fd_sc_hd__nor2_8
X_20524_ _18330_/X _20522_/X _20523_/X _18341_/X VGND VGND VPWR VPWR _20524_/X sky130_fd_sc_hd__a22o_1
X_27080_ _27080_/A VGND VGND VPWR VPWR _33956_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24292_ _24292_/A VGND VGND VPWR VPWR _32678_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26031_ _26031_/A VGND VGND VPWR VPWR _33469_/D sky130_fd_sc_hd__clkbuf_1
X_23243_ input45/X VGND VGND VPWR VPWR _23243_/X sky130_fd_sc_hd__buf_4
X_35229_ _35677_/CLK _35229_/D VGND VGND VPWR VPWR _35229_/Q sky130_fd_sc_hd__dfxtp_1
X_20455_ _20164_/X _20453_/X _20454_/X _20169_/X VGND VGND VPWR VPWR _20455_/X sky130_fd_sc_hd__a22o_1
XFILLER_181_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_335_CLK clkbuf_6_44__f_CLK/X VGND VGND VPWR VPWR _35961_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_105_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23174_ _23174_/A VGND VGND VPWR VPWR _32125_/D sky130_fd_sc_hd__clkbuf_1
X_20386_ _35471_/Q _35407_/Q _35343_/Q _35279_/Q _20260_/X _20261_/X VGND VGND VPWR
+ VPWR _20386_/X sky130_fd_sc_hd__mux4_1
XFILLER_106_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22125_ _33407_/Q _33343_/Q _33279_/Q _33215_/Q _22080_/X _22081_/X VGND VGND VPWR
+ VPWR _22125_/X sky130_fd_sc_hd__mux4_1
XFILLER_122_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27982_ _27982_/A VGND VGND VPWR VPWR _34328_/D sky130_fd_sc_hd__clkbuf_1
Xoutput160 _36197_/Q VGND VGND VPWR VPWR D2[15] sky130_fd_sc_hd__buf_2
XTAP_6526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput171 _36207_/Q VGND VGND VPWR VPWR D2[25] sky130_fd_sc_hd__buf_2
XFILLER_248_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput182 _36217_/Q VGND VGND VPWR VPWR D2[35] sky130_fd_sc_hd__buf_2
X_29721_ _29721_/A VGND VGND VPWR VPWR _35121_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput193 _36227_/Q VGND VGND VPWR VPWR D2[45] sky130_fd_sc_hd__buf_2
XFILLER_173_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26933_ _33894_/Q _23280_/X _26939_/S VGND VGND VPWR VPWR _26934_/A sky130_fd_sc_hd__mux2_1
X_22056_ _22012_/X _22054_/X _22055_/X _22018_/X VGND VGND VPWR VPWR _22056_/X sky130_fd_sc_hd__a22o_1
XTAP_6559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1075 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21007_ _20897_/X _21005_/X _21006_/X _20900_/X VGND VGND VPWR VPWR _21007_/X sky130_fd_sc_hd__a22o_1
X_29652_ _35089_/Q _29512_/X _29652_/S VGND VGND VPWR VPWR _29653_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26864_ _26864_/A VGND VGND VPWR VPWR _33861_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28603_ _27770_/X _34623_/Q _28619_/S VGND VGND VPWR VPWR _28604_/A sky130_fd_sc_hd__mux2_1
X_25815_ _25815_/A VGND VGND VPWR VPWR _33366_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29583_ _35056_/Q _29410_/X _29589_/S VGND VGND VPWR VPWR _29584_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26795_ _26795_/A VGND VGND VPWR VPWR _33828_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28534_ _28534_/A VGND VGND VPWR VPWR _34590_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25746_ _24899_/X _33334_/Q _25760_/S VGND VGND VPWR VPWR _25747_/A sky130_fd_sc_hd__mux2_1
X_22958_ _22958_/A VGND VGND VPWR VPWR _32044_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21909_ _21905_/X _21908_/X _21732_/X VGND VGND VPWR VPWR _21933_/A sky130_fd_sc_hd__o21ba_1
XFILLER_245_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28465_ _28513_/S VGND VGND VPWR VPWR _28484_/S sky130_fd_sc_hd__buf_4
X_22889_ _22879_/X _32022_/Q _22916_/S VGND VGND VPWR VPWR _22890_/A sky130_fd_sc_hd__mux2_1
X_25677_ _31823_/A _26352_/B VGND VGND VPWR VPWR _25810_/S sky130_fd_sc_hd__nand2_8
X_27416_ _27416_/A VGND VGND VPWR VPWR _34091_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24628_ _23036_/X _32838_/Q _24630_/S VGND VGND VPWR VPWR _24629_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28396_ _27664_/X _34525_/Q _28400_/S VGND VGND VPWR VPWR _28397_/A sky130_fd_sc_hd__mux2_1
XFILLER_223_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27347_ _34059_/Q _27199_/X _27359_/S VGND VGND VPWR VPWR _27348_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24559_ _22934_/X _32805_/Q _24567_/S VGND VGND VPWR VPWR _24560_/A sky130_fd_sc_hd__mux2_1
XFILLER_212_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17100_ _17096_/X _17099_/X _16779_/X VGND VGND VPWR VPWR _17122_/A sky130_fd_sc_hd__o21ba_1
XFILLER_7_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18080_ _32911_/Q _32847_/Q _32783_/Q _32719_/Q _15984_/X _15987_/X VGND VGND VPWR
+ VPWR _18080_/X sky130_fd_sc_hd__mux4_1
XFILLER_168_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27278_ _34026_/Q _27096_/X _27296_/S VGND VGND VPWR VPWR _27279_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29017_ _34818_/Q _27171_/X _29027_/S VGND VGND VPWR VPWR _29018_/A sky130_fd_sc_hd__mux2_1
X_17031_ _16706_/X _17029_/X _17030_/X _16712_/X VGND VGND VPWR VPWR _17031_/X sky130_fd_sc_hd__a22o_1
X_26229_ _24815_/X _33563_/Q _26237_/S VGND VGND VPWR VPWR _26230_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_326_CLK clkbuf_6_39__f_CLK/X VGND VGND VPWR VPWR _32887_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_194_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18982_ _18978_/X _18981_/X _18734_/X _18735_/X VGND VGND VPWR VPWR _18997_/B sky130_fd_sc_hd__o211a_1
XFILLER_112_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29919_ _29919_/A VGND VGND VPWR VPWR _35215_/D sky130_fd_sc_hd__clkbuf_1
X_17933_ _35210_/Q _35146_/Q _35082_/Q _32266_/Q _17716_/X _17717_/X VGND VGND VPWR
+ VPWR _17933_/X sky130_fd_sc_hd__mux4_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32930_ _36002_/CLK _32930_/D VGND VGND VPWR VPWR _32930_/Q sky130_fd_sc_hd__dfxtp_1
X_17864_ _17864_/A VGND VGND VPWR VPWR _17864_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_38_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19603_ _33657_/Q _33593_/Q _33529_/Q _33465_/Q _19500_/X _19501_/X VGND VGND VPWR
+ VPWR _19603_/X sky130_fd_sc_hd__mux4_1
XFILLER_113_1249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16815_ _16815_/A VGND VGND VPWR VPWR _31978_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32861_ _35870_/CLK _32861_/D VGND VGND VPWR VPWR _32861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17795_ _17791_/X _17794_/X _17518_/X VGND VGND VPWR VPWR _17796_/D sky130_fd_sc_hd__o21ba_1
XFILLER_226_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34600_ _35365_/CLK _34600_/D VGND VGND VPWR VPWR _34600_/Q sky130_fd_sc_hd__dfxtp_1
X_31812_ _31812_/A VGND VGND VPWR VPWR _36112_/D sky130_fd_sc_hd__clkbuf_1
X_19534_ _19528_/X _19533_/X _19465_/X VGND VGND VPWR VPWR _19535_/D sky130_fd_sc_hd__o21ba_1
X_16746_ _16500_/X _16744_/X _16745_/X _16503_/X VGND VGND VPWR VPWR _16746_/X sky130_fd_sc_hd__a22o_1
X_35580_ _35708_/CLK _35580_/D VGND VGND VPWR VPWR _35580_/Q sky130_fd_sc_hd__dfxtp_1
X_32792_ _33941_/CLK _32792_/D VGND VGND VPWR VPWR _32792_/Q sky130_fd_sc_hd__dfxtp_1
X_34531_ _36209_/CLK _34531_/D VGND VGND VPWR VPWR _34531_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31743_ _31743_/A VGND VGND VPWR VPWR _36079_/D sky130_fd_sc_hd__clkbuf_1
X_19465_ _20171_/A VGND VGND VPWR VPWR _19465_/X sky130_fd_sc_hd__buf_2
XFILLER_222_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16677_ _33127_/Q _36007_/Q _32999_/Q _32935_/Q _16356_/X _16357_/X VGND VGND VPWR
+ VPWR _16677_/X sky130_fd_sc_hd__mux4_1
X_18416_ _18410_/X _18415_/X _18315_/X VGND VGND VPWR VPWR _18438_/A sky130_fd_sc_hd__o21ba_1
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34462_ _36229_/CLK _34462_/D VGND VGND VPWR VPWR _34462_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31674_ _27819_/X _36047_/Q _31678_/S VGND VGND VPWR VPWR _31675_/A sky130_fd_sc_hd__mux2_1
X_19396_ _19146_/X _19392_/X _19395_/X _19151_/X VGND VGND VPWR VPWR _19396_/X sky130_fd_sc_hd__a22o_1
XFILLER_107_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36201_ _36207_/CLK _36201_/D VGND VGND VPWR VPWR _36201_/Q sky130_fd_sc_hd__dfxtp_1
X_33413_ _33415_/CLK _33413_/D VGND VGND VPWR VPWR _33413_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18347_ _18328_/X _18342_/X _18344_/X _18346_/X VGND VGND VPWR VPWR _18406_/B sky130_fd_sc_hd__o211a_1
X_30625_ _35550_/Q _29354_/X _30627_/S VGND VGND VPWR VPWR _30626_/A sky130_fd_sc_hd__mux2_1
X_34393_ _36121_/CLK _34393_/D VGND VGND VPWR VPWR _34393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36132_ _36136_/CLK _36132_/D VGND VGND VPWR VPWR _36132_/Q sky130_fd_sc_hd__dfxtp_1
X_33344_ _33921_/CLK _33344_/D VGND VGND VPWR VPWR _33344_/Q sky130_fd_sc_hd__dfxtp_1
X_18278_ _18278_/A VGND VGND VPWR VPWR _32021_/D sky130_fd_sc_hd__clkbuf_1
X_30556_ _30556_/A VGND VGND VPWR VPWR _35517_/D sky130_fd_sc_hd__clkbuf_1
X_36063_ _36128_/CLK _36063_/D VGND VGND VPWR VPWR _36063_/Q sky130_fd_sc_hd__dfxtp_1
Xinput40 DW[45] VGND VGND VPWR VPWR input40/X sky130_fd_sc_hd__buf_6
X_17229_ _17935_/A VGND VGND VPWR VPWR _17229_/X sky130_fd_sc_hd__buf_8
Xclkbuf_leaf_317_CLK clkbuf_6_37__f_CLK/X VGND VGND VPWR VPWR _32909_/CLK sky130_fd_sc_hd__clkbuf_16
X_33275_ _33531_/CLK _33275_/D VGND VGND VPWR VPWR _33275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30487_ _30487_/A VGND VGND VPWR VPWR _35484_/D sky130_fd_sc_hd__clkbuf_1
Xinput51 DW[55] VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__buf_12
Xinput62 DW[7] VGND VGND VPWR VPWR input62/X sky130_fd_sc_hd__buf_8
Xinput73 R2[2] VGND VGND VPWR VPWR input73/X sky130_fd_sc_hd__buf_4
X_35014_ _35525_/CLK _35014_/D VGND VGND VPWR VPWR _35014_/Q sky130_fd_sc_hd__dfxtp_1
Xinput84 RW[1] VGND VGND VPWR VPWR input84/X sky130_fd_sc_hd__clkbuf_4
X_20240_ _20234_/X _20239_/X _20171_/X VGND VGND VPWR VPWR _20241_/D sky130_fd_sc_hd__o21ba_1
X_32226_ _35716_/CLK _32226_/D VGND VGND VPWR VPWR _32226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20171_ _20171_/A VGND VGND VPWR VPWR _20171_/X sky130_fd_sc_hd__buf_2
X_32157_ _36223_/CLK _32157_/D VGND VGND VPWR VPWR _32157_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31108_ _35779_/Q input40/X _31116_/S VGND VGND VPWR VPWR _31109_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32088_ _32856_/CLK _32088_/D VGND VGND VPWR VPWR _32088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35916_ _35916_/CLK _35916_/D VGND VGND VPWR VPWR _35916_/Q sky130_fd_sc_hd__dfxtp_1
X_23930_ _23011_/X _32510_/Q _23948_/S VGND VGND VPWR VPWR _23931_/A sky130_fd_sc_hd__mux2_1
X_31039_ _35746_/Q input4/X _31053_/S VGND VGND VPWR VPWR _31040_/A sky130_fd_sc_hd__mux2_1
XFILLER_218_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_845 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23861_ _23861_/A VGND VGND VPWR VPWR _32477_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35847_ _35847_/CLK _35847_/D VGND VGND VPWR VPWR _35847_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22812_ _20648_/X _22810_/X _22811_/X _20658_/X VGND VGND VPWR VPWR _22812_/X sky130_fd_sc_hd__a22o_1
X_25600_ _24883_/X _33265_/Q _25604_/S VGND VGND VPWR VPWR _25601_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26580_ _26580_/A VGND VGND VPWR VPWR _33728_/D sky130_fd_sc_hd__clkbuf_1
X_23792_ _23840_/S VGND VGND VPWR VPWR _23811_/S sky130_fd_sc_hd__buf_4
XFILLER_37_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35778_ _35841_/CLK _35778_/D VGND VGND VPWR VPWR _35778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25531_ _25531_/A VGND VGND VPWR VPWR _33232_/D sky130_fd_sc_hd__clkbuf_1
X_22743_ _35729_/Q _32240_/Q _35601_/Q _35537_/Q _20593_/X _20595_/X VGND VGND VPWR
+ VPWR _22743_/X sky130_fd_sc_hd__mux4_1
XFILLER_168_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34729_ _34915_/CLK _34729_/D VGND VGND VPWR VPWR _34729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28250_ _28250_/A VGND VGND VPWR VPWR _34455_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25462_ _25462_/A VGND VGND VPWR VPWR _33199_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_240_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22674_ _22512_/X _22672_/X _22673_/X _22515_/X VGND VGND VPWR VPWR _22674_/X sky130_fd_sc_hd__a22o_1
XFILLER_13_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27201_ _27201_/A VGND VGND VPWR VPWR _33995_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24413_ _24524_/S VGND VGND VPWR VPWR _24432_/S sky130_fd_sc_hd__buf_4
XFILLER_16_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21625_ _22451_/A VGND VGND VPWR VPWR _21625_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25393_ _33168_/Q _23481_/X _25395_/S VGND VGND VPWR VPWR _25394_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28181_ _27745_/X _34423_/Q _28193_/S VGND VGND VPWR VPWR _28182_/A sky130_fd_sc_hd__mux2_1
X_24344_ _23015_/X _32703_/Q _24360_/S VGND VGND VPWR VPWR _24345_/A sky130_fd_sc_hd__mux2_1
X_27132_ _33973_/Q _27131_/X _27156_/S VGND VGND VPWR VPWR _27133_/A sky130_fd_sc_hd__mux2_1
XFILLER_205_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21556_ _21552_/X _21555_/X _21379_/X VGND VGND VPWR VPWR _21580_/A sky130_fd_sc_hd__o21ba_1
XFILLER_142_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20507_ _33107_/Q _32083_/Q _35859_/Q _35795_/Q _18379_/X _18380_/X VGND VGND VPWR
+ VPWR _20507_/X sky130_fd_sc_hd__mux4_1
X_27063_ _33951_/Q _27062_/X _27063_/S VGND VGND VPWR VPWR _27064_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_308_CLK clkbuf_6_50__f_CLK/X VGND VGND VPWR VPWR _36038_/CLK sky130_fd_sc_hd__clkbuf_16
X_24275_ _24275_/A VGND VGND VPWR VPWR _32670_/D sky130_fd_sc_hd__clkbuf_1
X_21487_ _33389_/Q _33325_/Q _33261_/Q _33197_/Q _21374_/X _21375_/X VGND VGND VPWR
+ VPWR _21487_/X sky130_fd_sc_hd__mux4_1
XFILLER_14_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26014_ _24896_/X _33461_/Q _26030_/S VGND VGND VPWR VPWR _26015_/A sky130_fd_sc_hd__mux2_1
X_23226_ input88/X input86/X input87/X VGND VGND VPWR VPWR _23227_/A sky130_fd_sc_hd__or3b_1
XFILLER_180_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20438_ _19453_/A _20436_/X _20437_/X _19456_/A VGND VGND VPWR VPWR _20438_/X sky130_fd_sc_hd__a22o_1
XTAP_7002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23157_ _22984_/X _32117_/Q _23173_/S VGND VGND VPWR VPWR _23158_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20369_ _33679_/Q _33615_/Q _33551_/Q _33487_/Q _20206_/X _20207_/X VGND VGND VPWR
+ VPWR _20369_/X sky130_fd_sc_hd__mux4_1
XTAP_6301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22108_ _35198_/Q _35134_/Q _35070_/Q _32254_/Q _21963_/X _21964_/X VGND VGND VPWR
+ VPWR _22108_/X sky130_fd_sc_hd__mux4_1
XFILLER_161_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27965_ _27825_/X _34321_/Q _27965_/S VGND VGND VPWR VPWR _27966_/A sky130_fd_sc_hd__mux2_1
XTAP_6345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23088_ _25132_/A input83/X input89/X _27232_/B VGND VGND VPWR VPWR _23089_/A sky130_fd_sc_hd__and4bb_1
XTAP_6356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29704_ _29704_/A VGND VGND VPWR VPWR _35113_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26916_ _33886_/Q _23255_/X _26918_/S VGND VGND VPWR VPWR _26917_/A sky130_fd_sc_hd__mux2_1
X_22039_ _34428_/Q _36156_/Q _34300_/Q _34236_/Q _21829_/X _21830_/X VGND VGND VPWR
+ VPWR _22039_/X sky130_fd_sc_hd__mux4_1
XTAP_6389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27896_ _27723_/X _34288_/Q _27902_/S VGND VGND VPWR VPWR _27897_/A sky130_fd_sc_hd__mux2_1
XFILLER_236_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29635_ _29635_/A VGND VGND VPWR VPWR _35080_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26847_ _26847_/A VGND VGND VPWR VPWR _33853_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16600_ _33381_/Q _33317_/Q _33253_/Q _33189_/Q _16421_/X _16422_/X VGND VGND VPWR
+ VPWR _16600_/X sky130_fd_sc_hd__mux4_1
XTAP_4987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17580_ _35200_/Q _35136_/Q _35072_/Q _32256_/Q _17363_/X _17364_/X VGND VGND VPWR
+ VPWR _17580_/X sky130_fd_sc_hd__mux4_1
X_29566_ _35048_/Q _29385_/X _29568_/S VGND VGND VPWR VPWR _29567_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26778_ _26778_/A VGND VGND VPWR VPWR _33820_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28517_ _27639_/X _34582_/Q _28535_/S VGND VGND VPWR VPWR _28518_/A sky130_fd_sc_hd__mux2_1
X_16531_ _33635_/Q _33571_/Q _33507_/Q _33443_/Q _16494_/X _16495_/X VGND VGND VPWR
+ VPWR _16531_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25729_ _24874_/X _33326_/Q _25739_/S VGND VGND VPWR VPWR _25730_/A sky130_fd_sc_hd__mux2_1
X_29497_ input50/X VGND VGND VPWR VPWR _29497_/X sky130_fd_sc_hd__buf_2
XFILLER_147_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19250_ _33647_/Q _33583_/Q _33519_/Q _33455_/Q _19147_/X _19148_/X VGND VGND VPWR
+ VPWR _19250_/X sky130_fd_sc_hd__mux4_1
X_16462_ _16462_/A VGND VGND VPWR VPWR _31968_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28448_ _28448_/A VGND VGND VPWR VPWR _34549_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18201_ _17158_/A _18199_/X _18200_/X _17163_/A VGND VGND VPWR VPWR _18201_/X sky130_fd_sc_hd__a22o_1
XPHY_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19181_ _19175_/X _19180_/X _19112_/X VGND VGND VPWR VPWR _19182_/D sky130_fd_sc_hd__o21ba_1
XPHY_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28379_ _28379_/A VGND VGND VPWR VPWR _34517_/D sky130_fd_sc_hd__clkbuf_1
X_16393_ _16147_/X _16391_/X _16392_/X _16150_/X VGND VGND VPWR VPWR _16393_/X sky130_fd_sc_hd__a22o_1
XPHY_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18132_ _33425_/Q _33361_/Q _33297_/Q _33233_/Q _17833_/X _17834_/X VGND VGND VPWR
+ VPWR _18132_/X sky130_fd_sc_hd__mux4_2
XFILLER_200_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30410_ _35448_/Q _29435_/X _30420_/S VGND VGND VPWR VPWR _30411_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31390_ _27797_/X _35912_/Q _31408_/S VGND VGND VPWR VPWR _31391_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18063_ _34446_/Q _36174_/Q _34318_/Q _34254_/Q _17935_/X _17936_/X VGND VGND VPWR
+ VPWR _18063_/X sky130_fd_sc_hd__mux4_1
X_30341_ _35415_/Q _29333_/X _30357_/S VGND VGND VPWR VPWR _30342_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17014_ _34416_/Q _36144_/Q _34288_/Q _34224_/Q _16876_/X _16877_/X VGND VGND VPWR
+ VPWR _17014_/X sky130_fd_sc_hd__mux4_1
XFILLER_176_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33060_ _35812_/CLK _33060_/D VGND VGND VPWR VPWR _33060_/Q sky130_fd_sc_hd__dfxtp_1
X_30272_ _30272_/A VGND VGND VPWR VPWR _35382_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_217_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32011_ _36202_/CLK _32011_/D VGND VGND VPWR VPWR _32011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18965_ _18965_/A _18965_/B _18965_/C _18965_/D VGND VGND VPWR VPWR _18966_/A sky130_fd_sc_hd__or4_2
XFILLER_234_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17916_ _17912_/X _17913_/X _17914_/X _17915_/X VGND VGND VPWR VPWR _17916_/X sky130_fd_sc_hd__a22o_1
XFILLER_67_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33962_ _35627_/CLK _33962_/D VGND VGND VPWR VPWR _33962_/Q sky130_fd_sc_hd__dfxtp_1
X_18896_ _18896_/A VGND VGND VPWR VPWR _32420_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32913_ _32913_/CLK _32913_/D VGND VGND VPWR VPWR _32913_/Q sky130_fd_sc_hd__dfxtp_1
X_35701_ _35701_/CLK _35701_/D VGND VGND VPWR VPWR _35701_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17847_ _17847_/A VGND VGND VPWR VPWR _17847_/X sky130_fd_sc_hd__clkbuf_4
X_33893_ _35622_/CLK _33893_/D VGND VGND VPWR VPWR _33893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32844_ _32909_/CLK _32844_/D VGND VGND VPWR VPWR _32844_/Q sky130_fd_sc_hd__dfxtp_1
X_35632_ _35632_/CLK _35632_/D VGND VGND VPWR VPWR _35632_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17778_ _17773_/X _17775_/X _17776_/X _17777_/X VGND VGND VPWR VPWR _17778_/X sky130_fd_sc_hd__a22o_1
XFILLER_78_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19517_ _19367_/X _19515_/X _19516_/X _19371_/X VGND VGND VPWR VPWR _19517_/X sky130_fd_sc_hd__a22o_1
XFILLER_240_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35563_ _35691_/CLK _35563_/D VGND VGND VPWR VPWR _35563_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16729_ _16723_/X _16728_/X _16445_/X VGND VGND VPWR VPWR _16737_/C sky130_fd_sc_hd__o21ba_1
XFILLER_228_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32775_ _32905_/CLK _32775_/D VGND VGND VPWR VPWR _32775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34514_ _36115_/CLK _34514_/D VGND VGND VPWR VPWR _34514_/Q sky130_fd_sc_hd__dfxtp_1
X_31726_ _31726_/A VGND VGND VPWR VPWR _36071_/D sky130_fd_sc_hd__clkbuf_1
X_19448_ _35444_/Q _35380_/Q _35316_/Q _35252_/Q _19201_/X _19202_/X VGND VGND VPWR
+ VPWR _19448_/X sky130_fd_sc_hd__mux4_1
XFILLER_23_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35494_ _35559_/CLK _35494_/D VGND VGND VPWR VPWR _35494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34445_ _34956_/CLK _34445_/D VGND VGND VPWR VPWR _34445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31657_ _27794_/X _36039_/Q _31657_/S VGND VGND VPWR VPWR _31658_/A sky130_fd_sc_hd__mux2_1
X_19379_ _20236_/A VGND VGND VPWR VPWR _19379_/X sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_94_CLK clkbuf_leaf_96_CLK/A VGND VGND VPWR VPWR _36205_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_50_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21410_ _21763_/A VGND VGND VPWR VPWR _21410_/X sky130_fd_sc_hd__buf_2
XFILLER_202_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30608_ _30740_/S VGND VGND VPWR VPWR _30627_/S sky130_fd_sc_hd__buf_6
XFILLER_37_1194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34376_ _34633_/CLK _34376_/D VGND VGND VPWR VPWR _34376_/Q sky130_fd_sc_hd__dfxtp_1
X_22390_ _35206_/Q _35142_/Q _35078_/Q _32262_/Q _22316_/X _22317_/X VGND VGND VPWR
+ VPWR _22390_/X sky130_fd_sc_hd__mux4_1
XFILLER_202_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31588_ _27692_/X _36006_/Q _31594_/S VGND VGND VPWR VPWR _31589_/A sky130_fd_sc_hd__mux2_1
XFILLER_176_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36115_ _36115_/CLK _36115_/D VGND VGND VPWR VPWR _36115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21341_ _22561_/A VGND VGND VPWR VPWR _21341_/X sky130_fd_sc_hd__buf_4
X_33327_ _36080_/CLK _33327_/D VGND VGND VPWR VPWR _33327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30539_ _35509_/Q _29426_/X _30555_/S VGND VGND VPWR VPWR _30540_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36046_ _36047_/CLK _36046_/D VGND VGND VPWR VPWR _36046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24060_ _24060_/A VGND VGND VPWR VPWR _32571_/D sky130_fd_sc_hd__clkbuf_1
X_21272_ _22451_/A VGND VGND VPWR VPWR _21272_/X sky130_fd_sc_hd__buf_4
X_33258_ _36075_/CLK _33258_/D VGND VGND VPWR VPWR _33258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23011_ input35/X VGND VGND VPWR VPWR _23011_/X sky130_fd_sc_hd__buf_2
XFILLER_11_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20223_ _20073_/X _20221_/X _20222_/X _20077_/X VGND VGND VPWR VPWR _20223_/X sky130_fd_sc_hd__a22o_1
X_32209_ _35124_/CLK _32209_/D VGND VGND VPWR VPWR _32209_/Q sky130_fd_sc_hd__dfxtp_1
X_33189_ _36070_/CLK _33189_/D VGND VGND VPWR VPWR _33189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20154_ _35464_/Q _35400_/Q _35336_/Q _35272_/Q _19907_/X _19908_/X VGND VGND VPWR
+ VPWR _20154_/X sky130_fd_sc_hd__mux4_1
XFILLER_98_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27750_ _27750_/A VGND VGND VPWR VPWR _34232_/D sky130_fd_sc_hd__clkbuf_1
X_20085_ _20236_/A VGND VGND VPWR VPWR _20085_/X sky130_fd_sc_hd__clkbuf_4
X_24962_ _24961_/X _32970_/Q _24983_/S VGND VGND VPWR VPWR _24963_/A sky130_fd_sc_hd__mux2_1
XTAP_4206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_246_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26701_ _33784_/Q _23402_/X _26711_/S VGND VGND VPWR VPWR _26702_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_942 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23913_ _22987_/X _32502_/Q _23927_/S VGND VGND VPWR VPWR _23914_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27681_ _27680_/X _34210_/Q _27702_/S VGND VGND VPWR VPWR _27682_/A sky130_fd_sc_hd__mux2_1
XTAP_3516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24893_ _24995_/S VGND VGND VPWR VPWR _24921_/S sky130_fd_sc_hd__buf_4
XTAP_3527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29420_ _34995_/Q _29419_/X _29420_/S VGND VGND VPWR VPWR _29421_/A sky130_fd_sc_hd__mux2_1
X_26632_ _33751_/Q _23234_/X _26648_/S VGND VGND VPWR VPWR _26633_/A sky130_fd_sc_hd__mux2_1
XTAP_3538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23844_ _31418_/A _28380_/A VGND VGND VPWR VPWR _23977_/S sky130_fd_sc_hd__nand2_8
XTAP_3549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29351_ input62/X VGND VGND VPWR VPWR _29351_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26563_ _26563_/A VGND VGND VPWR VPWR _33720_/D sky130_fd_sc_hd__clkbuf_1
X_23775_ _23775_/A VGND VGND VPWR VPWR _32373_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20987_ _22560_/A VGND VGND VPWR VPWR _20987_/X sky130_fd_sc_hd__buf_6
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28302_ _28302_/A VGND VGND VPWR VPWR _34480_/D sky130_fd_sc_hd__clkbuf_1
X_25514_ _24954_/X _33224_/Q _25532_/S VGND VGND VPWR VPWR _25515_/A sky130_fd_sc_hd__mux2_1
XFILLER_198_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22726_ _22722_/X _22725_/X _22471_/X VGND VGND VPWR VPWR _22727_/D sky130_fd_sc_hd__o21ba_1
X_29282_ _29282_/A VGND VGND VPWR VPWR _34943_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26494_ _26494_/A VGND VGND VPWR VPWR _33687_/D sky130_fd_sc_hd__clkbuf_1
X_28233_ _27822_/X _34448_/Q _28235_/S VGND VGND VPWR VPWR _28234_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_22 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22657_ _33102_/Q _32078_/Q _35854_/Q _35790_/Q _22384_/X _22385_/X VGND VGND VPWR
+ VPWR _22657_/X sky130_fd_sc_hd__mux4_1
X_25445_ _25445_/A VGND VGND VPWR VPWR _33191_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_213_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_85_CLK clkbuf_leaf_88_CLK/A VGND VGND VPWR VPWR _33119_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_201_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21608_ _21602_/X _21607_/X _21398_/X VGND VGND VPWR VPWR _21618_/C sky130_fd_sc_hd__o21ba_1
XFILLER_167_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28164_ _27720_/X _34415_/Q _28172_/S VGND VGND VPWR VPWR _28165_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25376_ _25403_/S VGND VGND VPWR VPWR _25395_/S sky130_fd_sc_hd__buf_4
X_22588_ _32908_/Q _32844_/Q _32780_/Q _32716_/Q _22299_/X _22300_/X VGND VGND VPWR
+ VPWR _22588_/X sky130_fd_sc_hd__mux4_1
XFILLER_142_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27115_ input19/X VGND VGND VPWR VPWR _27115_/X sky130_fd_sc_hd__buf_2
XFILLER_182_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21539_ _22598_/A VGND VGND VPWR VPWR _21539_/X sky130_fd_sc_hd__buf_6
XFILLER_103_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24327_ _22990_/X _32695_/Q _24339_/S VGND VGND VPWR VPWR _24328_/A sky130_fd_sc_hd__mux2_1
X_28095_ _28095_/A VGND VGND VPWR VPWR _34382_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24258_ _22879_/X _32662_/Q _24276_/S VGND VGND VPWR VPWR _24259_/A sky130_fd_sc_hd__mux2_1
X_27046_ _27046_/A VGND VGND VPWR VPWR _33945_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23209_ _23061_/X _32142_/Q _23215_/S VGND VGND VPWR VPWR _23210_/A sky130_fd_sc_hd__mux2_1
XFILLER_175_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24189_ _32631_/Q _23399_/X _24201_/S VGND VGND VPWR VPWR _24190_/A sky130_fd_sc_hd__mux2_1
XFILLER_175_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28997_ _28997_/A VGND VGND VPWR VPWR _34808_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18750_ _19456_/A VGND VGND VPWR VPWR _18750_/X sky130_fd_sc_hd__buf_4
X_27948_ _27948_/A VGND VGND VPWR VPWR _34312_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17701_ _32900_/Q _32836_/Q _32772_/Q _32708_/Q _17699_/X _17700_/X VGND VGND VPWR
+ VPWR _17701_/X sky130_fd_sc_hd__mux4_1
XFILLER_209_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18681_ _34910_/Q _34846_/Q _34782_/Q _34718_/Q _18396_/X _18398_/X VGND VGND VPWR
+ VPWR _18681_/X sky130_fd_sc_hd__mux4_1
XFILLER_237_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27879_ _27698_/X _34280_/Q _27881_/S VGND VGND VPWR VPWR _27880_/A sky130_fd_sc_hd__mux2_1
XFILLER_236_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29618_ _29618_/A VGND VGND VPWR VPWR _35072_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17632_ _17412_/X _17630_/X _17631_/X _17418_/X VGND VGND VPWR VPWR _17632_/X sky130_fd_sc_hd__a22o_1
XFILLER_48_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30890_ _30890_/A VGND VGND VPWR VPWR _35675_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17563_ _17559_/X _17560_/X _17561_/X _17562_/X VGND VGND VPWR VPWR _17563_/X sky130_fd_sc_hd__a22o_1
XFILLER_1_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29549_ _29660_/S VGND VGND VPWR VPWR _29568_/S sky130_fd_sc_hd__buf_6
XFILLER_91_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_1442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19302_ _19298_/X _19299_/X _19300_/X _19301_/X VGND VGND VPWR VPWR _19302_/X sky130_fd_sc_hd__a22o_1
XFILLER_210_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16514_ _35618_/Q _34978_/Q _34338_/Q _33698_/Q _16438_/X _16439_/X VGND VGND VPWR
+ VPWR _16514_/X sky130_fd_sc_hd__mux4_1
XFILLER_95_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32560_ _35952_/CLK _32560_/D VGND VGND VPWR VPWR _32560_/Q sky130_fd_sc_hd__dfxtp_1
X_17494_ _17847_/A VGND VGND VPWR VPWR _17494_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_147_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31511_ _31511_/A VGND VGND VPWR VPWR _35969_/D sky130_fd_sc_hd__clkbuf_1
X_19233_ _35630_/Q _34990_/Q _34350_/Q _33710_/Q _19091_/X _19092_/X VGND VGND VPWR
+ VPWR _19233_/X sky130_fd_sc_hd__mux4_1
X_16445_ _17857_/A VGND VGND VPWR VPWR _16445_/X sky130_fd_sc_hd__buf_2
XFILLER_204_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32491_ _35947_/CLK _32491_/D VGND VGND VPWR VPWR _32491_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_76_CLK clkbuf_leaf_77_CLK/A VGND VGND VPWR VPWR _35997_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_158_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34230_ _35126_/CLK _34230_/D VGND VGND VPWR VPWR _34230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_1052 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31442_ _31442_/A VGND VGND VPWR VPWR _35936_/D sky130_fd_sc_hd__clkbuf_1
X_19164_ _19014_/X _19162_/X _19163_/X _19018_/X VGND VGND VPWR VPWR _19164_/X sky130_fd_sc_hd__a22o_1
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16376_ _16370_/X _16375_/X _16075_/X VGND VGND VPWR VPWR _16384_/C sky130_fd_sc_hd__o21ba_1
XFILLER_129_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18115_ _15981_/X _18113_/X _18114_/X _15991_/X VGND VGND VPWR VPWR _18115_/X sky130_fd_sc_hd__a22o_1
XFILLER_9_974 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34161_ _35635_/CLK _34161_/D VGND VGND VPWR VPWR _34161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31373_ _27773_/X _35904_/Q _31387_/S VGND VGND VPWR VPWR _31374_/A sky130_fd_sc_hd__mux2_1
X_19095_ _35434_/Q _35370_/Q _35306_/Q _35242_/Q _18848_/X _18849_/X VGND VGND VPWR
+ VPWR _19095_/X sky130_fd_sc_hd__mux4_1
XFILLER_157_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33112_ _35992_/CLK _33112_/D VGND VGND VPWR VPWR _33112_/Q sky130_fd_sc_hd__dfxtp_1
X_30324_ _30324_/A VGND VGND VPWR VPWR _35407_/D sky130_fd_sc_hd__clkbuf_1
X_18046_ _32654_/Q _32590_/Q _32526_/Q _35982_/Q _17982_/X _17766_/X VGND VGND VPWR
+ VPWR _18046_/X sky130_fd_sc_hd__mux4_1
X_34092_ _34093_/CLK _34092_/D VGND VGND VPWR VPWR _34092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33043_ _35859_/CLK _33043_/D VGND VGND VPWR VPWR _33043_/Q sky130_fd_sc_hd__dfxtp_1
X_30255_ _30255_/A VGND VGND VPWR VPWR _35374_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30186_ _35342_/Q _29503_/X _30192_/S VGND VGND VPWR VPWR _30187_/A sky130_fd_sc_hd__mux2_1
X_19997_ _19712_/X _19995_/X _19996_/X _19718_/X VGND VGND VPWR VPWR _19997_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_1108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18948_ _20162_/A VGND VGND VPWR VPWR _18948_/X sky130_fd_sc_hd__clkbuf_4
X_34994_ _35764_/CLK _34994_/D VGND VGND VPWR VPWR _34994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33945_ _36219_/CLK _33945_/D VGND VGND VPWR VPWR _33945_/Q sky130_fd_sc_hd__dfxtp_1
X_18879_ _35684_/Q _32191_/Q _35556_/Q _35492_/Q _18558_/X _18559_/X VGND VGND VPWR
+ VPWR _18879_/X sky130_fd_sc_hd__mux4_1
XFILLER_132_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1078 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20910_ _20691_/X _20908_/X _20909_/X _20701_/X VGND VGND VPWR VPWR _20910_/X sky130_fd_sc_hd__a22o_1
X_33876_ _33941_/CLK _33876_/D VGND VGND VPWR VPWR _33876_/Q sky130_fd_sc_hd__dfxtp_1
X_21890_ _21603_/X _21888_/X _21889_/X _21606_/X VGND VGND VPWR VPWR _21890_/X sky130_fd_sc_hd__a22o_1
XFILLER_81_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20841_ _20837_/X _20840_/X _20704_/X VGND VGND VPWR VPWR _20842_/D sky130_fd_sc_hd__o21ba_1
X_35615_ _35615_/CLK _35615_/D VGND VGND VPWR VPWR _35615_/Q sky130_fd_sc_hd__dfxtp_1
X_32827_ _32891_/CLK _32827_/D VGND VGND VPWR VPWR _32827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23560_ _23560_/A VGND VGND VPWR VPWR _32274_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20772_ _34392_/Q _36120_/Q _34264_/Q _34200_/Q _20770_/X _20771_/X VGND VGND VPWR
+ VPWR _20772_/X sky130_fd_sc_hd__mux4_1
XFILLER_223_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35546_ _35609_/CLK _35546_/D VGND VGND VPWR VPWR _35546_/Q sky130_fd_sc_hd__dfxtp_1
X_32758_ _32887_/CLK _32758_/D VGND VGND VPWR VPWR _32758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22511_ _22505_/X _22508_/X _22509_/X _22510_/X VGND VGND VPWR VPWR _22511_/X sky130_fd_sc_hd__a22o_1
XFILLER_39_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31709_ _31709_/A VGND VGND VPWR VPWR _36063_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35477_ _36055_/CLK _35477_/D VGND VGND VPWR VPWR _35477_/Q sky130_fd_sc_hd__dfxtp_1
X_23491_ _23491_/A VGND VGND VPWR VPWR _32242_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_67_CLK clkbuf_leaf_73_CLK/A VGND VGND VPWR VPWR _35989_/CLK sky130_fd_sc_hd__clkbuf_16
X_32689_ _35953_/CLK _32689_/D VGND VGND VPWR VPWR _32689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_241_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25230_ _33091_/Q _23438_/X _25238_/S VGND VGND VPWR VPWR _25231_/A sky130_fd_sc_hd__mux2_1
X_22442_ _22365_/X _22440_/X _22441_/X _22371_/X VGND VGND VPWR VPWR _22442_/X sky130_fd_sc_hd__a22o_1
X_34428_ _36157_/CLK _34428_/D VGND VGND VPWR VPWR _34428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25161_ _33058_/Q _23268_/X _25175_/S VGND VGND VPWR VPWR _25162_/A sky130_fd_sc_hd__mux2_1
XFILLER_136_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22373_ _22373_/A VGND VGND VPWR VPWR _22373_/X sky130_fd_sc_hd__clkbuf_4
X_34359_ _35768_/CLK _34359_/D VGND VGND VPWR VPWR _34359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24112_ _24112_/A VGND VGND VPWR VPWR _32596_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21324_ _35432_/Q _35368_/Q _35304_/Q _35240_/Q _21148_/X _21149_/X VGND VGND VPWR
+ VPWR _21324_/X sky130_fd_sc_hd__mux4_1
X_25092_ _25092_/A VGND VGND VPWR VPWR _33026_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28920_ _28920_/A VGND VGND VPWR VPWR _34772_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24043_ _24043_/A VGND VGND VPWR VPWR _32563_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21255_ _21249_/X _21254_/X _21045_/X VGND VGND VPWR VPWR _21265_/C sky130_fd_sc_hd__o21ba_1
X_36029_ _36029_/CLK _36029_/D VGND VGND VPWR VPWR _36029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20206_ _20206_/A VGND VGND VPWR VPWR _20206_/X sky130_fd_sc_hd__buf_6
X_28851_ _28851_/A VGND VGND VPWR VPWR _34739_/D sky130_fd_sc_hd__clkbuf_1
X_21186_ _22598_/A VGND VGND VPWR VPWR _21186_/X sky130_fd_sc_hd__buf_6
XFILLER_89_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27802_ _27801_/X _34249_/Q _27826_/S VGND VGND VPWR VPWR _27803_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20137_ _19859_/X _20135_/X _20136_/X _19862_/X VGND VGND VPWR VPWR _20137_/X sky130_fd_sc_hd__a22o_1
X_28782_ _34708_/Q _27226_/X _28784_/S VGND VGND VPWR VPWR _28783_/A sky130_fd_sc_hd__mux2_1
X_25994_ _25994_/A VGND VGND VPWR VPWR _33451_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27733_ _27732_/X _34227_/Q _27733_/S VGND VGND VPWR VPWR _27734_/A sky130_fd_sc_hd__mux2_1
XFILLER_219_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24945_ input42/X VGND VGND VPWR VPWR _24945_/X sky130_fd_sc_hd__buf_4
X_20068_ _20286_/A VGND VGND VPWR VPWR _20068_/X sky130_fd_sc_hd__buf_4
XTAP_4036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27664_ input62/X VGND VGND VPWR VPWR _27664_/X sky130_fd_sc_hd__buf_4
XFILLER_73_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24876_ _24876_/A VGND VGND VPWR VPWR _32942_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29403_ _29403_/A VGND VGND VPWR VPWR _34989_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26615_ _26615_/A VGND VGND VPWR VPWR _33745_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23827_ _23827_/A VGND VGND VPWR VPWR _32398_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27595_ _27595_/A VGND VGND VPWR VPWR _34176_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29334_ _34967_/Q _29333_/X _29358_/S VGND VGND VPWR VPWR _29335_/A sky130_fd_sc_hd__mux2_1
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26546_ _26546_/A VGND VGND VPWR VPWR _33712_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23758_ _23758_/A VGND VGND VPWR VPWR _32365_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22709_ _32144_/Q _32336_/Q _32400_/Q _35920_/Q _22586_/X _21611_/A VGND VGND VPWR
+ VPWR _22709_/X sky130_fd_sc_hd__mux4_1
X_29265_ _29265_/A VGND VGND VPWR VPWR _34935_/D sky130_fd_sc_hd__clkbuf_1
X_26477_ _26477_/A VGND VGND VPWR VPWR _33680_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23689_ _23689_/A VGND VGND VPWR VPWR _32334_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_58_CLK clkbuf_leaf_61_CLK/A VGND VGND VPWR VPWR _35946_/CLK sky130_fd_sc_hd__clkbuf_16
X_28216_ _28243_/S VGND VGND VPWR VPWR _28235_/S sky130_fd_sc_hd__buf_4
X_16230_ _33050_/Q _32026_/Q _35802_/Q _35738_/Q _16067_/X _16069_/X VGND VGND VPWR
+ VPWR _16230_/X sky130_fd_sc_hd__mux4_1
XFILLER_220_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25428_ _25428_/A VGND VGND VPWR VPWR _33183_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29196_ _29196_/A VGND VGND VPWR VPWR _34902_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_761 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16161_ _35608_/Q _34968_/Q _34328_/Q _33688_/Q _16053_/X _16055_/X VGND VGND VPWR
+ VPWR _16161_/X sky130_fd_sc_hd__mux4_1
X_28147_ _27695_/X _34407_/Q _28151_/S VGND VGND VPWR VPWR _28148_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25359_ _25359_/A VGND VGND VPWR VPWR _33151_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16092_ _17716_/A VGND VGND VPWR VPWR _16092_/X sky130_fd_sc_hd__clkbuf_8
X_28078_ _28078_/A VGND VGND VPWR VPWR _34374_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27029_ _33940_/Q _23495_/X _27031_/S VGND VGND VPWR VPWR _27030_/A sky130_fd_sc_hd__mux2_1
X_19920_ _19920_/A _19920_/B _19920_/C _19920_/D VGND VGND VPWR VPWR _19921_/A sky130_fd_sc_hd__or4_4
XFILLER_108_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30040_ _30040_/A VGND VGND VPWR VPWR _35272_/D sky130_fd_sc_hd__clkbuf_1
X_19851_ _19851_/A VGND VGND VPWR VPWR _32447_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_122_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18802_ _33890_/Q _33826_/Q _33762_/Q _36066_/Q _18618_/X _18619_/X VGND VGND VPWR
+ VPWR _18802_/X sky130_fd_sc_hd__mux4_1
X_19782_ _33406_/Q _33342_/Q _33278_/Q _33214_/Q _19780_/X _19781_/X VGND VGND VPWR
+ VPWR _19782_/X sky130_fd_sc_hd__mux4_1
XFILLER_122_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16994_ _17834_/A VGND VGND VPWR VPWR _16994_/X sky130_fd_sc_hd__clkbuf_4
X_18733_ _18661_/X _18731_/X _18732_/X _18665_/X VGND VGND VPWR VPWR _18733_/X sky130_fd_sc_hd__a22o_1
XTAP_5260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31991_ _34405_/CLK _31991_/D VGND VGND VPWR VPWR _31991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33730_ _35458_/CLK _33730_/D VGND VGND VPWR VPWR _33730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18664_ _32862_/Q _32798_/Q _32734_/Q _32670_/Q _18587_/X _18588_/X VGND VGND VPWR
+ VPWR _18664_/X sky130_fd_sc_hd__mux4_1
X_30942_ _35700_/Q input24/X _30960_/S VGND VGND VPWR VPWR _30943_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17615_ _17506_/X _17613_/X _17614_/X _17509_/X VGND VGND VPWR VPWR _17615_/X sky130_fd_sc_hd__a22o_1
XTAP_4592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_990 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33661_ _33661_/CLK _33661_/D VGND VGND VPWR VPWR _33661_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30873_ _35668_/Q input59/X _30875_/S VGND VGND VPWR VPWR _30874_/A sky130_fd_sc_hd__mux2_1
X_18595_ _20162_/A VGND VGND VPWR VPWR _18595_/X sky130_fd_sc_hd__buf_4
XTAP_3880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35400_ _35466_/CLK _35400_/D VGND VGND VPWR VPWR _35400_/Q sky130_fd_sc_hd__dfxtp_1
X_32612_ _36007_/CLK _32612_/D VGND VGND VPWR VPWR _32612_/Q sky130_fd_sc_hd__dfxtp_1
X_17546_ _34431_/Q _36159_/Q _34303_/Q _34239_/Q _17229_/X _17230_/X VGND VGND VPWR
+ VPWR _17546_/X sky130_fd_sc_hd__mux4_1
XFILLER_45_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33592_ _35641_/CLK _33592_/D VGND VGND VPWR VPWR _33592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_233_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35331_ _35651_/CLK _35331_/D VGND VGND VPWR VPWR _35331_/Q sky130_fd_sc_hd__dfxtp_1
X_32543_ _35998_/CLK _32543_/D VGND VGND VPWR VPWR _32543_/Q sky130_fd_sc_hd__dfxtp_1
X_17477_ _33662_/Q _33598_/Q _33534_/Q _33470_/Q _17200_/X _17201_/X VGND VGND VPWR
+ VPWR _17477_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_49_CLK clkbuf_leaf_49_CLK/A VGND VGND VPWR VPWR _36011_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_20_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_1450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19216_ _33646_/Q _33582_/Q _33518_/Q _33454_/Q _19147_/X _19148_/X VGND VGND VPWR
+ VPWR _19216_/X sky130_fd_sc_hd__mux4_1
XFILLER_32_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_6_53__f_CLK clkbuf_5_26_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_53__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_16428_ _32608_/Q _32544_/Q _32480_/Q _35936_/Q _16217_/X _16354_/X VGND VGND VPWR
+ VPWR _16428_/X sky130_fd_sc_hd__mux4_1
X_35262_ _35453_/CLK _35262_/D VGND VGND VPWR VPWR _35262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32474_ _36055_/CLK _32474_/D VGND VGND VPWR VPWR _32474_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_912 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34213_ _34405_/CLK _34213_/D VGND VGND VPWR VPWR _34213_/Q sky130_fd_sc_hd__dfxtp_1
X_31425_ _31425_/A VGND VGND VPWR VPWR _35928_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19147_ _20206_/A VGND VGND VPWR VPWR _19147_/X sky130_fd_sc_hd__buf_4
X_16359_ _17910_/A VGND VGND VPWR VPWR _16359_/X sky130_fd_sc_hd__clkbuf_4
X_35193_ _35193_/CLK _35193_/D VGND VGND VPWR VPWR _35193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34144_ _34594_/CLK _34144_/D VGND VGND VPWR VPWR _34144_/Q sky130_fd_sc_hd__dfxtp_1
X_19078_ _18800_/X _19076_/X _19077_/X _18803_/X VGND VGND VPWR VPWR _19078_/X sky130_fd_sc_hd__a22o_1
X_31356_ _27748_/X _35896_/Q _31366_/S VGND VGND VPWR VPWR _31357_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18029_ _18025_/X _18028_/X _17857_/X VGND VGND VPWR VPWR _18037_/C sky130_fd_sc_hd__o21ba_1
X_30307_ _30307_/A VGND VGND VPWR VPWR _35399_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34075_ _36212_/CLK _34075_/D VGND VGND VPWR VPWR _34075_/Q sky130_fd_sc_hd__dfxtp_1
X_31287_ _27646_/X _35863_/Q _31303_/S VGND VGND VPWR VPWR _31288_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33026_ _36034_/CLK _33026_/D VGND VGND VPWR VPWR _33026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21040_ _35616_/Q _34976_/Q _34336_/Q _33696_/Q _21038_/X _21039_/X VGND VGND VPWR
+ VPWR _21040_/X sky130_fd_sc_hd__mux4_1
X_30238_ _30238_/A VGND VGND VPWR VPWR _35366_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30169_ _35334_/Q _29478_/X _30171_/S VGND VGND VPWR VPWR _30170_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34977_ _35618_/CLK _34977_/D VGND VGND VPWR VPWR _34977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22991_ _22990_/X _32055_/Q _23009_/S VGND VGND VPWR VPWR _22992_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24730_ _22987_/X _32886_/Q _24744_/S VGND VGND VPWR VPWR _24731_/A sky130_fd_sc_hd__mux2_1
X_33928_ _36104_/CLK _33928_/D VGND VGND VPWR VPWR _33928_/Q sky130_fd_sc_hd__dfxtp_1
X_21942_ _32634_/Q _32570_/Q _32506_/Q _35962_/Q _21876_/X _21660_/X VGND VGND VPWR
+ VPWR _21942_/X sky130_fd_sc_hd__mux4_1
XFILLER_131_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24661_ _28110_/A _31553_/B VGND VGND VPWR VPWR _24794_/S sky130_fd_sc_hd__nand2_8
XFILLER_15_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21873_ _33912_/Q _33848_/Q _33784_/Q _36088_/Q _21624_/X _21625_/X VGND VGND VPWR
+ VPWR _21873_/X sky130_fd_sc_hd__mux4_1
X_33859_ _36100_/CLK _33859_/D VGND VGND VPWR VPWR _33859_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26400_ _26400_/A VGND VGND VPWR VPWR _33643_/D sky130_fd_sc_hd__clkbuf_1
X_20824_ _20630_/X _20822_/X _20823_/X _20641_/X VGND VGND VPWR VPWR _20824_/X sky130_fd_sc_hd__a22o_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23612_ _23702_/S VGND VGND VPWR VPWR _23631_/S sky130_fd_sc_hd__buf_4
X_27380_ _27380_/A VGND VGND VPWR VPWR _34074_/D sky130_fd_sc_hd__clkbuf_1
X_24592_ _24592_/A VGND VGND VPWR VPWR _32820_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26331_ _26331_/A VGND VGND VPWR VPWR _33611_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_223_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20755_ _20618_/X _20753_/X _20754_/X _20627_/X VGND VGND VPWR VPWR _20755_/X sky130_fd_sc_hd__a22o_1
X_23543_ _32266_/Q _23463_/X _23557_/S VGND VGND VPWR VPWR _23544_/A sky130_fd_sc_hd__mux2_1
X_35529_ _35658_/CLK _35529_/D VGND VGND VPWR VPWR _35529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29050_ _34834_/Q _27220_/X _29056_/S VGND VGND VPWR VPWR _29051_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23474_ _23474_/A VGND VGND VPWR VPWR _32236_/D sky130_fd_sc_hd__clkbuf_1
X_26262_ _26262_/A VGND VGND VPWR VPWR _33578_/D sky130_fd_sc_hd__clkbuf_1
X_20686_ _35158_/Q _35094_/Q _35030_/Q _32150_/Q _20683_/X _20685_/X VGND VGND VPWR
+ VPWR _20686_/X sky130_fd_sc_hd__mux4_1
XFILLER_195_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28001_ _28001_/A VGND VGND VPWR VPWR _34337_/D sky130_fd_sc_hd__clkbuf_1
X_22425_ _34951_/Q _34887_/Q _34823_/Q _34759_/Q _22113_/X _22114_/X VGND VGND VPWR
+ VPWR _22425_/X sky130_fd_sc_hd__mux4_1
XFILLER_183_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25213_ _33083_/Q _23411_/X _25217_/S VGND VGND VPWR VPWR _25214_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26193_ _24961_/X _33546_/Q _26207_/S VGND VGND VPWR VPWR _26194_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22356_ _22356_/A _22356_/B _22356_/C _22356_/D VGND VGND VPWR VPWR _22357_/A sky130_fd_sc_hd__or4_4
X_25144_ _33050_/Q _23243_/X _25154_/S VGND VGND VPWR VPWR _25145_/A sky130_fd_sc_hd__mux2_1
XFILLER_237_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21307_ _22366_/A VGND VGND VPWR VPWR _21307_/X sky130_fd_sc_hd__clkbuf_4
X_29952_ _35231_/Q _29357_/X _29952_/S VGND VGND VPWR VPWR _29953_/A sky130_fd_sc_hd__mux2_1
X_25075_ _25075_/A VGND VGND VPWR VPWR _33018_/D sky130_fd_sc_hd__clkbuf_1
X_22287_ _22287_/A VGND VGND VPWR VPWR _36227_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_959 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28903_ _34764_/Q _27202_/X _28913_/S VGND VGND VPWR VPWR _28904_/A sky130_fd_sc_hd__mux2_1
X_24026_ _22953_/X _32555_/Q _24042_/S VGND VGND VPWR VPWR _24027_/A sky130_fd_sc_hd__mux2_1
X_21238_ _20953_/X _21236_/X _21237_/X _20959_/X VGND VGND VPWR VPWR _21238_/X sky130_fd_sc_hd__a22o_1
X_29883_ _35198_/Q _29453_/X _29901_/S VGND VGND VPWR VPWR _29884_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28834_ _34731_/Q _27100_/X _28850_/S VGND VGND VPWR VPWR _28835_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21169_ _21165_/X _21168_/X _21026_/X VGND VGND VPWR VPWR _21195_/A sky130_fd_sc_hd__o21ba_1
XFILLER_133_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28765_ _28765_/A VGND VGND VPWR VPWR _34699_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25977_ _25977_/A VGND VGND VPWR VPWR _33443_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_995 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27716_ _27716_/A VGND VGND VPWR VPWR _34221_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24928_ _24927_/X _32959_/Q _24952_/S VGND VGND VPWR VPWR _24929_/A sky130_fd_sc_hd__mux2_1
XTAP_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28696_ _28696_/A VGND VGND VPWR VPWR _34666_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_248_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27647_ _27646_/X _34199_/Q _27671_/S VGND VGND VPWR VPWR _27648_/A sky130_fd_sc_hd__mux2_1
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24859_ _24858_/X _32937_/Q _24859_/S VGND VGND VPWR VPWR _24860_/A sky130_fd_sc_hd__mux2_1
XTAP_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17400_ _34939_/Q _34875_/Q _34811_/Q _34747_/Q _17160_/X _17161_/X VGND VGND VPWR
+ VPWR _17400_/X sky130_fd_sc_hd__mux4_1
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18380_ _20236_/A VGND VGND VPWR VPWR _18380_/X sky130_fd_sc_hd__buf_6
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27578_ _27578_/A VGND VGND VPWR VPWR _34168_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29317_ _29317_/A VGND VGND VPWR VPWR _34960_/D sky130_fd_sc_hd__clkbuf_1
X_17331_ _17158_/X _17329_/X _17330_/X _17163_/X VGND VGND VPWR VPWR _17331_/X sky130_fd_sc_hd__a22o_1
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26529_ _26529_/A VGND VGND VPWR VPWR _33704_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29248_ _29248_/A VGND VGND VPWR VPWR _34927_/D sky130_fd_sc_hd__clkbuf_1
X_17262_ _17153_/X _17260_/X _17261_/X _17156_/X VGND VGND VPWR VPWR _17262_/X sky130_fd_sc_hd__a22o_1
XFILLER_105_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19001_ _18793_/X _18999_/X _19000_/X _18798_/X VGND VGND VPWR VPWR _19001_/X sky130_fd_sc_hd__a22o_1
XFILLER_197_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16213_ _33370_/Q _33306_/Q _33242_/Q _33178_/Q _16002_/X _16003_/X VGND VGND VPWR
+ VPWR _16213_/X sky130_fd_sc_hd__mux4_1
XFILLER_122_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29179_ _34895_/Q _27211_/X _29183_/S VGND VGND VPWR VPWR _29180_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17193_ _34421_/Q _36149_/Q _34293_/Q _34229_/Q _16876_/X _16877_/X VGND VGND VPWR
+ VPWR _17193_/X sky130_fd_sc_hd__mux4_1
XFILLER_155_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31210_ _27732_/X _35827_/Q _31210_/S VGND VGND VPWR VPWR _31211_/A sky130_fd_sc_hd__mux2_1
X_16144_ _34136_/Q _34072_/Q _34008_/Q _33944_/Q _16009_/X _16011_/X VGND VGND VPWR
+ VPWR _16144_/X sky130_fd_sc_hd__mux4_1
XFILLER_60_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32190_ _35684_/CLK _32190_/D VGND VGND VPWR VPWR _32190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31141_ _35795_/Q input58/X _31145_/S VGND VGND VPWR VPWR _31142_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16075_ _17857_/A VGND VGND VPWR VPWR _16075_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19903_ _19899_/X _19902_/X _19793_/X _19794_/X VGND VGND VPWR VPWR _19920_/B sky130_fd_sc_hd__o211a_1
XFILLER_29_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31072_ _35762_/Q input21/X _31074_/S VGND VGND VPWR VPWR _31073_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34900_ _34964_/CLK _34900_/D VGND VGND VPWR VPWR _34900_/Q sky130_fd_sc_hd__dfxtp_1
X_30023_ _30023_/A VGND VGND VPWR VPWR _35264_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19834_ _19720_/X _19832_/X _19833_/X _19724_/X VGND VGND VPWR VPWR _19834_/X sky130_fd_sc_hd__a22o_1
XFILLER_233_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35880_ _35947_/CLK _35880_/D VGND VGND VPWR VPWR _35880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_867 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34831_ _34961_/CLK _34831_/D VGND VGND VPWR VPWR _34831_/Q sky130_fd_sc_hd__dfxtp_1
X_16977_ _34927_/Q _34863_/Q _34799_/Q _34735_/Q _16807_/X _16808_/X VGND VGND VPWR
+ VPWR _16977_/X sky130_fd_sc_hd__mux4_1
X_19765_ _33085_/Q _32061_/Q _35837_/Q _35773_/Q _19731_/X _19732_/X VGND VGND VPWR
+ VPWR _19765_/X sky130_fd_sc_hd__mux4_1
Xinput5 DW[13] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__buf_8
X_18716_ _18716_/A _18716_/B _18716_/C _18716_/D VGND VGND VPWR VPWR _18717_/A sky130_fd_sc_hd__or4_4
XFILLER_37_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34762_ _34957_/CLK _34762_/D VGND VGND VPWR VPWR _34762_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31974_ _34085_/CLK _31974_/D VGND VGND VPWR VPWR _31974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19696_ _34683_/Q _34619_/Q _34555_/Q _34491_/Q _19592_/X _19593_/X VGND VGND VPWR
+ VPWR _19696_/X sky130_fd_sc_hd__mux4_1
XFILLER_37_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18647_ _34142_/Q _34078_/Q _34014_/Q _33950_/Q _18309_/X _18311_/X VGND VGND VPWR
+ VPWR _18647_/X sky130_fd_sc_hd__mux4_1
XFILLER_36_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33713_ _35633_/CLK _33713_/D VGND VGND VPWR VPWR _33713_/Q sky130_fd_sc_hd__dfxtp_1
X_30925_ _35692_/Q input15/X _30939_/S VGND VGND VPWR VPWR _30926_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34693_ _34693_/CLK _34693_/D VGND VGND VPWR VPWR _34693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_818 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30856_ _30856_/A VGND VGND VPWR VPWR _35659_/D sky130_fd_sc_hd__clkbuf_1
X_18578_ _18440_/X _18576_/X _18577_/X _18445_/X VGND VGND VPWR VPWR _18578_/X sky130_fd_sc_hd__a22o_1
X_33644_ _34093_/CLK _33644_/D VGND VGND VPWR VPWR _33644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_212_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17529_ _32639_/Q _32575_/Q _32511_/Q _35967_/Q _17276_/X _17413_/X VGND VGND VPWR
+ VPWR _17529_/X sky130_fd_sc_hd__mux4_1
X_33575_ _36073_/CLK _33575_/D VGND VGND VPWR VPWR _33575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30787_ _30787_/A VGND VGND VPWR VPWR _35626_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20540_ _34708_/Q _34644_/Q _34580_/Q _34516_/Q _20298_/X _20299_/X VGND VGND VPWR
+ VPWR _20540_/X sky130_fd_sc_hd__mux4_1
X_32526_ _35982_/CLK _32526_/D VGND VGND VPWR VPWR _32526_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35314_ _35828_/CLK _35314_/D VGND VGND VPWR VPWR _35314_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_242_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20471_ _19458_/A _20469_/X _20470_/X _19463_/A VGND VGND VPWR VPWR _20471_/X sky130_fd_sc_hd__a22o_1
X_32457_ _36076_/CLK _32457_/D VGND VGND VPWR VPWR _32457_/Q sky130_fd_sc_hd__dfxtp_1
X_35245_ _35566_/CLK _35245_/D VGND VGND VPWR VPWR _35245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22210_ _33089_/Q _32065_/Q _35841_/Q _35777_/Q _22031_/X _22032_/X VGND VGND VPWR
+ VPWR _22210_/X sky130_fd_sc_hd__mux4_1
X_31408_ _27825_/X _35921_/Q _31408_/S VGND VGND VPWR VPWR _31409_/A sky130_fd_sc_hd__mux2_1
X_23190_ _23033_/X _32133_/Q _23194_/S VGND VGND VPWR VPWR _23191_/A sky130_fd_sc_hd__mux2_1
X_35176_ _35176_/CLK _35176_/D VGND VGND VPWR VPWR _35176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32388_ _35973_/CLK _32388_/D VGND VGND VPWR VPWR _32388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34127_ _34192_/CLK _34127_/D VGND VGND VPWR VPWR _34127_/Q sky130_fd_sc_hd__dfxtp_1
X_22141_ _21956_/X _22139_/X _22140_/X _21959_/X VGND VGND VPWR VPWR _22141_/X sky130_fd_sc_hd__a22o_1
X_31339_ _27723_/X _35888_/Q _31345_/S VGND VGND VPWR VPWR _31340_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34058_ _34187_/CLK _34058_/D VGND VGND VPWR VPWR _34058_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22072_ _34941_/Q _34877_/Q _34813_/Q _34749_/Q _21760_/X _21761_/X VGND VGND VPWR
+ VPWR _22072_/X sky130_fd_sc_hd__mux4_1
XTAP_6719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25900_ _24927_/X _33407_/Q _25916_/S VGND VGND VPWR VPWR _25901_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21023_ _33376_/Q _33312_/Q _33248_/Q _33184_/Q _21021_/X _21022_/X VGND VGND VPWR
+ VPWR _21023_/X sky130_fd_sc_hd__mux4_1
XFILLER_47_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33009_ _36016_/CLK _33009_/D VGND VGND VPWR VPWR _33009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26880_ _33869_/Q _23472_/X _26888_/S VGND VGND VPWR VPWR _26881_/A sky130_fd_sc_hd__mux2_1
X_25831_ _25831_/A VGND VGND VPWR VPWR _33374_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28550_ _27692_/X _34598_/Q _28556_/S VGND VGND VPWR VPWR _28551_/A sky130_fd_sc_hd__mux2_1
X_25762_ _25810_/S VGND VGND VPWR VPWR _25781_/S sky130_fd_sc_hd__buf_4
XFILLER_216_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22974_ input21/X VGND VGND VPWR VPWR _22974_/X sky130_fd_sc_hd__buf_2
XFILLER_210_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27501_ _27501_/A VGND VGND VPWR VPWR _34132_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24713_ _22962_/X _32878_/Q _24723_/S VGND VGND VPWR VPWR _24714_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28481_ _28481_/A VGND VGND VPWR VPWR _34565_/D sky130_fd_sc_hd__clkbuf_1
X_21925_ _21921_/X _21924_/X _21751_/X VGND VGND VPWR VPWR _21933_/C sky130_fd_sc_hd__o21ba_1
X_25693_ _24821_/X _33309_/Q _25697_/S VGND VGND VPWR VPWR _25694_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27432_ _27432_/A VGND VGND VPWR VPWR _34099_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24644_ _24644_/A VGND VGND VPWR VPWR _32845_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21856_ _35447_/Q _35383_/Q _35319_/Q _35255_/Q _21854_/X _21855_/X VGND VGND VPWR
+ VPWR _21856_/X sky130_fd_sc_hd__mux4_1
XFILLER_215_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27363_ _34067_/Q _27223_/X _27367_/S VGND VGND VPWR VPWR _27364_/A sky130_fd_sc_hd__mux2_1
X_20807_ _20803_/X _20806_/X _20704_/X VGND VGND VPWR VPWR _20808_/D sky130_fd_sc_hd__o21ba_1
XFILLER_168_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24575_ _24575_/A VGND VGND VPWR VPWR _32812_/D sky130_fd_sc_hd__clkbuf_1
X_21787_ _33077_/Q _32053_/Q _35829_/Q _35765_/Q _21678_/X _21679_/X VGND VGND VPWR
+ VPWR _21787_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29102_ _34858_/Q _27096_/X _29120_/S VGND VGND VPWR VPWR _29103_/A sky130_fd_sc_hd__mux2_1
X_26314_ _26314_/A VGND VGND VPWR VPWR _33603_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_212_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23526_ _32258_/Q _23435_/X _23536_/S VGND VGND VPWR VPWR _23527_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20738_ _20738_/A _20738_/B _20738_/C _20738_/D VGND VGND VPWR VPWR _20739_/A sky130_fd_sc_hd__or4_2
X_27294_ _34034_/Q _27121_/X _27296_/S VGND VGND VPWR VPWR _27295_/A sky130_fd_sc_hd__mux2_1
XFILLER_243_1099 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29033_ _29033_/A VGND VGND VPWR VPWR _34825_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26245_ _26245_/A VGND VGND VPWR VPWR _33570_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20669_ _22536_/A VGND VGND VPWR VPWR _20669_/X sky130_fd_sc_hd__buf_4
X_23457_ _23565_/S VGND VGND VPWR VPWR _23515_/S sky130_fd_sc_hd__buf_4
XFILLER_171_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22408_ _33159_/Q _36039_/Q _33031_/Q _32967_/Q _22368_/X _22369_/X VGND VGND VPWR
+ VPWR _22408_/X sky130_fd_sc_hd__mux4_1
X_26176_ _24936_/X _33538_/Q _26186_/S VGND VGND VPWR VPWR _26177_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23388_ _23499_/S VGND VGND VPWR VPWR _23418_/S sky130_fd_sc_hd__buf_8
XFILLER_87_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25127_ _25127_/A VGND VGND VPWR VPWR _33043_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22339_ _32901_/Q _32837_/Q _32773_/Q _32709_/Q _22299_/X _22300_/X VGND VGND VPWR
+ VPWR _22339_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29935_ _29935_/A VGND VGND VPWR VPWR _35222_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25058_ _25058_/A VGND VGND VPWR VPWR _33010_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16900_ _16645_/X _16898_/X _16899_/X _16648_/X VGND VGND VPWR VPWR _16900_/X sky130_fd_sc_hd__a22o_1
X_24009_ _22928_/X _32547_/Q _24021_/S VGND VGND VPWR VPWR _24010_/A sky130_fd_sc_hd__mux2_1
X_17880_ _17559_/X _17878_/X _17879_/X _17562_/X VGND VGND VPWR VPWR _17880_/X sky130_fd_sc_hd__a22o_1
X_29866_ _35190_/Q _29429_/X _29880_/S VGND VGND VPWR VPWR _29867_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16831_ _35627_/Q _34987_/Q _34347_/Q _33707_/Q _16791_/X _16792_/X VGND VGND VPWR
+ VPWR _16831_/X sky130_fd_sc_hd__mux4_1
X_28817_ _34723_/Q _27075_/X _28829_/S VGND VGND VPWR VPWR _28818_/A sky130_fd_sc_hd__mux2_1
X_29797_ _29797_/A _30877_/B VGND VGND VPWR VPWR _29930_/S sky130_fd_sc_hd__nor2_8
XFILLER_78_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19550_ _19546_/X _19549_/X _19440_/X _19441_/X VGND VGND VPWR VPWR _19567_/B sky130_fd_sc_hd__o211a_1
XFILLER_247_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28748_ _28748_/A VGND VGND VPWR VPWR _34691_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16762_ _34665_/Q _34601_/Q _34537_/Q _34473_/Q _16586_/X _16587_/X VGND VGND VPWR
+ VPWR _16762_/X sky130_fd_sc_hd__mux4_1
XFILLER_76_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18501_ _34649_/Q _34585_/Q _34521_/Q _34457_/Q _18379_/X _18380_/X VGND VGND VPWR
+ VPWR _18501_/X sky130_fd_sc_hd__mux4_1
X_19481_ _19367_/X _19479_/X _19480_/X _19371_/X VGND VGND VPWR VPWR _19481_/X sky130_fd_sc_hd__a22o_1
XFILLER_111_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16693_ _34407_/Q _36135_/Q _34279_/Q _34215_/Q _16523_/X _16524_/X VGND VGND VPWR
+ VPWR _16693_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28679_ _28679_/A VGND VGND VPWR VPWR _34658_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18432_ _35159_/Q _35095_/Q _35031_/Q _32151_/Q _18383_/X _18385_/X VGND VGND VPWR
+ VPWR _18432_/X sky130_fd_sc_hd__mux4_1
X_30710_ _30710_/A VGND VGND VPWR VPWR _35590_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31690_ _36054_/Q input1/X _31708_/S VGND VGND VPWR VPWR _31691_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_1218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18363_ _18363_/A VGND VGND VPWR VPWR _20151_/A sky130_fd_sc_hd__buf_12
X_30641_ _30641_/A VGND VGND VPWR VPWR _35557_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17314_ _32889_/Q _32825_/Q _32761_/Q _32697_/Q _16993_/X _16994_/X VGND VGND VPWR
+ VPWR _17314_/X sky130_fd_sc_hd__mux4_1
X_33360_ _34186_/CLK _33360_/D VGND VGND VPWR VPWR _33360_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18294_ _18363_/A VGND VGND VPWR VPWR _20100_/A sky130_fd_sc_hd__buf_12
XFILLER_186_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30572_ _35525_/Q _29475_/X _30576_/S VGND VGND VPWR VPWR _30573_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32311_ _35895_/CLK _32311_/D VGND VGND VPWR VPWR _32311_/Q sky130_fd_sc_hd__dfxtp_1
X_17245_ _33143_/Q _36023_/Q _33015_/Q _32951_/Q _17062_/X _17063_/X VGND VGND VPWR
+ VPWR _17245_/X sky130_fd_sc_hd__mux4_1
X_33291_ _34186_/CLK _33291_/D VGND VGND VPWR VPWR _33291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35030_ _36118_/CLK _35030_/D VGND VGND VPWR VPWR _35030_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32242_ _36149_/CLK _32242_/D VGND VGND VPWR VPWR _32242_/Q sky130_fd_sc_hd__dfxtp_1
X_17176_ _32629_/Q _32565_/Q _32501_/Q _35957_/Q _16923_/X _17060_/X VGND VGND VPWR
+ VPWR _17176_/X sky130_fd_sc_hd__mux4_1
XFILLER_128_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16127_ _35415_/Q _35351_/Q _35287_/Q _35223_/Q _16062_/X _16064_/X VGND VGND VPWR
+ VPWR _16127_/X sky130_fd_sc_hd__mux4_1
XFILLER_116_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32173_ _35181_/CLK _32173_/D VGND VGND VPWR VPWR _32173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31124_ _31124_/A VGND VGND VPWR VPWR _35786_/D sky130_fd_sc_hd__clkbuf_1
X_16058_ _17862_/A VGND VGND VPWR VPWR _16058_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35932_ _35998_/CLK _35932_/D VGND VGND VPWR VPWR _35932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31055_ _31145_/S VGND VGND VPWR VPWR _31074_/S sky130_fd_sc_hd__buf_4
X_30006_ _30006_/A VGND VGND VPWR VPWR _35256_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_229_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19817_ _19811_/X _19812_/X _19815_/X _19816_/X VGND VGND VPWR VPWR _19817_/X sky130_fd_sc_hd__a22o_1
X_35863_ _35863_/CLK _35863_/D VGND VGND VPWR VPWR _35863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34814_ _36161_/CLK _34814_/D VGND VGND VPWR VPWR _34814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19748_ _34173_/Q _34109_/Q _34045_/Q _33981_/Q _19746_/X _19747_/X VGND VGND VPWR
+ VPWR _19748_/X sky130_fd_sc_hd__mux4_1
X_35794_ _35858_/CLK _35794_/D VGND VGND VPWR VPWR _35794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34745_ _36152_/CLK _34745_/D VGND VGND VPWR VPWR _34745_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31957_ _31957_/A VGND VGND VPWR VPWR _36181_/D sky130_fd_sc_hd__clkbuf_1
X_19679_ _33915_/Q _33851_/Q _33787_/Q _36091_/Q _19677_/X _19678_/X VGND VGND VPWR
+ VPWR _19679_/X sky130_fd_sc_hd__mux4_1
XFILLER_53_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_280_CLK clkbuf_6_59__f_CLK/X VGND VGND VPWR VPWR _35648_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_25_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21710_ _21598_/X _21708_/X _21709_/X _21601_/X VGND VGND VPWR VPWR _21710_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22690_ _34703_/Q _34639_/Q _34575_/Q _34511_/Q _22598_/X _22599_/X VGND VGND VPWR
+ VPWR _22690_/X sky130_fd_sc_hd__mux4_1
XFILLER_168_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30908_ _35684_/Q input6/X _30918_/S VGND VGND VPWR VPWR _30909_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34676_ _35829_/CLK _34676_/D VGND VGND VPWR VPWR _34676_/Q sky130_fd_sc_hd__dfxtp_1
X_31888_ _23387_/X _36148_/Q _31906_/S VGND VGND VPWR VPWR _31889_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21641_ _21603_/X _21639_/X _21640_/X _21606_/X VGND VGND VPWR VPWR _21641_/X sky130_fd_sc_hd__a22o_1
X_33627_ _36211_/CLK _33627_/D VGND VGND VPWR VPWR _33627_/Q sky130_fd_sc_hd__dfxtp_1
X_30839_ _30839_/A VGND VGND VPWR VPWR _35651_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24360_ _23039_/X _32711_/Q _24360_/S VGND VGND VPWR VPWR _24361_/A sky130_fd_sc_hd__mux2_1
X_21572_ _21568_/X _21571_/X _21398_/X VGND VGND VPWR VPWR _21580_/C sky130_fd_sc_hd__o21ba_1
X_33558_ _35861_/CLK _33558_/D VGND VGND VPWR VPWR _33558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20523_ _33940_/Q _33876_/Q _33812_/Q _36116_/Q _18362_/X _18364_/X VGND VGND VPWR
+ VPWR _20523_/X sky130_fd_sc_hd__mux4_1
X_23311_ _23311_/A VGND VGND VPWR VPWR _29662_/B sky130_fd_sc_hd__buf_6
XFILLER_36_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24291_ _22937_/X _32678_/Q _24297_/S VGND VGND VPWR VPWR _24292_/A sky130_fd_sc_hd__mux2_1
X_32509_ _35965_/CLK _32509_/D VGND VGND VPWR VPWR _32509_/Q sky130_fd_sc_hd__dfxtp_1
X_33489_ _34441_/CLK _33489_/D VGND VGND VPWR VPWR _33489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26030_ _24920_/X _33469_/Q _26030_/S VGND VGND VPWR VPWR _26031_/A sky130_fd_sc_hd__mux2_1
X_20454_ _34961_/Q _34897_/Q _34833_/Q _34769_/Q _20166_/X _20167_/X VGND VGND VPWR
+ VPWR _20454_/X sky130_fd_sc_hd__mux4_1
X_23242_ _23242_/A VGND VGND VPWR VPWR _32153_/D sky130_fd_sc_hd__clkbuf_1
X_35228_ _35613_/CLK _35228_/D VGND VGND VPWR VPWR _35228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23173_ _23008_/X _32125_/Q _23173_/S VGND VGND VPWR VPWR _23174_/A sky130_fd_sc_hd__mux2_1
X_35159_ _36118_/CLK _35159_/D VGND VGND VPWR VPWR _35159_/Q sky130_fd_sc_hd__dfxtp_1
X_20385_ _18281_/X _20383_/X _20384_/X _18291_/X VGND VGND VPWR VPWR _20385_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22124_ _21799_/X _22122_/X _22123_/X _21804_/X VGND VGND VPWR VPWR _22124_/X sky130_fd_sc_hd__a22o_1
XTAP_6505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27981_ _34328_/Q _27041_/X _27995_/S VGND VGND VPWR VPWR _27982_/A sky130_fd_sc_hd__mux2_1
Xoutput150 _31964_/Q VGND VGND VPWR VPWR D1[6] sky130_fd_sc_hd__buf_2
XTAP_6516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput161 _36198_/Q VGND VGND VPWR VPWR D2[16] sky130_fd_sc_hd__buf_2
XFILLER_133_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput172 _36208_/Q VGND VGND VPWR VPWR D2[26] sky130_fd_sc_hd__buf_2
X_29720_ _35121_/Q _29413_/X _29724_/S VGND VGND VPWR VPWR _29721_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput183 _36218_/Q VGND VGND VPWR VPWR D2[36] sky130_fd_sc_hd__buf_2
X_26932_ _26932_/A VGND VGND VPWR VPWR _33893_/D sky130_fd_sc_hd__clkbuf_1
X_22055_ _33149_/Q _36029_/Q _33021_/Q _32957_/Q _22015_/X _22016_/X VGND VGND VPWR
+ VPWR _22055_/X sky130_fd_sc_hd__mux4_1
XTAP_6549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput194 _36228_/Q VGND VGND VPWR VPWR D2[46] sky130_fd_sc_hd__buf_2
XTAP_5815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21006_ _33055_/Q _32031_/Q _35807_/Q _35743_/Q _20972_/X _20973_/X VGND VGND VPWR
+ VPWR _21006_/X sky130_fd_sc_hd__mux4_1
XFILLER_47_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29651_ _29651_/A VGND VGND VPWR VPWR _35088_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26863_ _33861_/Q _23444_/X _26867_/S VGND VGND VPWR VPWR _26864_/A sky130_fd_sc_hd__mux2_1
XTAP_5848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28602_ _28602_/A VGND VGND VPWR VPWR _34622_/D sky130_fd_sc_hd__clkbuf_1
X_25814_ _24796_/X _33366_/Q _25832_/S VGND VGND VPWR VPWR _25815_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29582_ _29582_/A VGND VGND VPWR VPWR _35055_/D sky130_fd_sc_hd__clkbuf_1
X_26794_ _33828_/Q _23274_/X _26804_/S VGND VGND VPWR VPWR _26795_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28533_ _27667_/X _34590_/Q _28535_/S VGND VGND VPWR VPWR _28534_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_1464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25745_ _25745_/A VGND VGND VPWR VPWR _33333_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22957_ _22956_/X _32044_/Q _22978_/S VGND VGND VPWR VPWR _22958_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_271_CLK clkbuf_6_57__f_CLK/X VGND VGND VPWR VPWR _35655_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_16_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_244_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21908_ _21806_/X _21906_/X _21907_/X _21809_/X VGND VGND VPWR VPWR _21908_/X sky130_fd_sc_hd__a22o_1
X_28464_ _28464_/A VGND VGND VPWR VPWR _34557_/D sky130_fd_sc_hd__clkbuf_1
X_25676_ _25676_/A VGND VGND VPWR VPWR _33301_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22888_ _23083_/S VGND VGND VPWR VPWR _22916_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_15_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27415_ _34091_/Q _27100_/X _27431_/S VGND VGND VPWR VPWR _27416_/A sky130_fd_sc_hd__mux2_1
XFILLER_231_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24627_ _24627_/A VGND VGND VPWR VPWR _32837_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28395_ _28395_/A VGND VGND VPWR VPWR _34524_/D sky130_fd_sc_hd__clkbuf_1
X_21839_ _21799_/X _21837_/X _21838_/X _21804_/X VGND VGND VPWR VPWR _21839_/X sky130_fd_sc_hd__a22o_1
XFILLER_197_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27346_ _27346_/A VGND VGND VPWR VPWR _34058_/D sky130_fd_sc_hd__clkbuf_1
X_24558_ _24558_/A VGND VGND VPWR VPWR _32804_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_1186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23509_ _32250_/Q _23408_/X _23515_/S VGND VGND VPWR VPWR _23510_/A sky130_fd_sc_hd__mux2_1
X_27277_ _27367_/S VGND VGND VPWR VPWR _27296_/S sky130_fd_sc_hd__buf_4
XFILLER_12_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24489_ _23030_/X _32772_/Q _24495_/S VGND VGND VPWR VPWR _24490_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29016_ _29016_/A VGND VGND VPWR VPWR _34817_/D sky130_fd_sc_hd__clkbuf_1
X_17030_ _33137_/Q _36017_/Q _33009_/Q _32945_/Q _16709_/X _16710_/X VGND VGND VPWR
+ VPWR _17030_/X sky130_fd_sc_hd__mux4_1
X_26228_ _26228_/A VGND VGND VPWR VPWR _33562_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26159_ _24911_/X _33530_/Q _26165_/S VGND VGND VPWR VPWR _26160_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18981_ _18661_/X _18979_/X _18980_/X _18665_/X VGND VGND VPWR VPWR _18981_/X sky130_fd_sc_hd__a22o_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17932_ _34698_/Q _34634_/Q _34570_/Q _34506_/Q _17645_/X _17646_/X VGND VGND VPWR
+ VPWR _17932_/X sky130_fd_sc_hd__mux4_1
X_29918_ _35215_/Q _29506_/X _29922_/S VGND VGND VPWR VPWR _29919_/A sky130_fd_sc_hd__mux2_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17863_ _17859_/X _17860_/X _17861_/X _17862_/X VGND VGND VPWR VPWR _17863_/X sky130_fd_sc_hd__a22o_1
XFILLER_23_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_984 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29849_ _35182_/Q _29404_/X _29859_/S VGND VGND VPWR VPWR _29850_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19602_ _19602_/A VGND VGND VPWR VPWR _32440_/D sky130_fd_sc_hd__buf_2
XFILLER_38_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16814_ _16814_/A _16814_/B _16814_/C _16814_/D VGND VGND VPWR VPWR _16815_/A sky130_fd_sc_hd__or4_4
X_17794_ _17511_/X _17792_/X _17793_/X _17516_/X VGND VGND VPWR VPWR _17794_/X sky130_fd_sc_hd__a22o_1
X_32860_ _36053_/CLK _32860_/D VGND VGND VPWR VPWR _32860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31811_ _36112_/Q input54/X _31813_/S VGND VGND VPWR VPWR _31812_/A sky130_fd_sc_hd__mux2_1
XFILLER_207_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16745_ _33897_/Q _33833_/Q _33769_/Q _36073_/Q _16671_/X _16672_/X VGND VGND VPWR
+ VPWR _16745_/X sky130_fd_sc_hd__mux4_1
X_19533_ _19458_/X _19531_/X _19532_/X _19463_/X VGND VGND VPWR VPWR _19533_/X sky130_fd_sc_hd__a22o_1
X_32791_ _32856_/CLK _32791_/D VGND VGND VPWR VPWR _32791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_235_874 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_262_CLK clkbuf_6_62__f_CLK/X VGND VGND VPWR VPWR _33415_/CLK sky130_fd_sc_hd__clkbuf_16
X_31742_ _36079_/Q input18/X _31750_/S VGND VGND VPWR VPWR _31743_/A sky130_fd_sc_hd__mux2_1
X_19464_ _19458_/X _19459_/X _19462_/X _19463_/X VGND VGND VPWR VPWR _19464_/X sky130_fd_sc_hd__a22o_1
X_34530_ _36209_/CLK _34530_/D VGND VGND VPWR VPWR _34530_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16676_ _32615_/Q _32551_/Q _32487_/Q _35943_/Q _16570_/X _16354_/X VGND VGND VPWR
+ VPWR _16676_/X sky130_fd_sc_hd__mux4_1
XFILLER_228_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18415_ _18301_/X _18411_/X _18414_/X _18307_/X VGND VGND VPWR VPWR _18415_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34461_ _36229_/CLK _34461_/D VGND VGND VPWR VPWR _34461_/Q sky130_fd_sc_hd__dfxtp_1
X_31673_ _31673_/A VGND VGND VPWR VPWR _36046_/D sky130_fd_sc_hd__clkbuf_1
X_19395_ _34163_/Q _34099_/Q _34035_/Q _33971_/Q _19393_/X _19394_/X VGND VGND VPWR
+ VPWR _19395_/X sky130_fd_sc_hd__mux4_1
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_938 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36200_ _36202_/CLK _36200_/D VGND VGND VPWR VPWR _36200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_1392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33412_ _33415_/CLK _33412_/D VGND VGND VPWR VPWR _33412_/Q sky130_fd_sc_hd__dfxtp_1
X_30624_ _30624_/A VGND VGND VPWR VPWR _35549_/D sky130_fd_sc_hd__clkbuf_1
X_18346_ _20147_/A VGND VGND VPWR VPWR _18346_/X sky130_fd_sc_hd__buf_4
X_34392_ _34904_/CLK _34392_/D VGND VGND VPWR VPWR _34392_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33343_ _36096_/CLK _33343_/D VGND VGND VPWR VPWR _33343_/Q sky130_fd_sc_hd__dfxtp_1
X_36131_ _36210_/CLK _36131_/D VGND VGND VPWR VPWR _36131_/Q sky130_fd_sc_hd__dfxtp_1
X_18277_ _18277_/A _18277_/B _18277_/C _18277_/D VGND VGND VPWR VPWR _18278_/A sky130_fd_sc_hd__or4_4
X_30555_ _35517_/Q _29450_/X _30555_/S VGND VGND VPWR VPWR _30556_/A sky130_fd_sc_hd__mux2_1
X_17228_ _17153_/X _17226_/X _17227_/X _17156_/X VGND VGND VPWR VPWR _17228_/X sky130_fd_sc_hd__a22o_1
X_36062_ _36207_/CLK _36062_/D VGND VGND VPWR VPWR _36062_/Q sky130_fd_sc_hd__dfxtp_1
X_33274_ _33914_/CLK _33274_/D VGND VGND VPWR VPWR _33274_/Q sky130_fd_sc_hd__dfxtp_1
Xinput30 DW[36] VGND VGND VPWR VPWR input30/X sky130_fd_sc_hd__buf_4
XFILLER_162_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30486_ _35484_/Q _29348_/X _30492_/S VGND VGND VPWR VPWR _30487_/A sky130_fd_sc_hd__mux2_1
Xinput41 DW[46] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__buf_6
XFILLER_116_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput52 DW[56] VGND VGND VPWR VPWR input52/X sky130_fd_sc_hd__clkbuf_16
Xinput63 DW[8] VGND VGND VPWR VPWR input63/X sky130_fd_sc_hd__buf_8
XFILLER_200_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35013_ _35525_/CLK _35013_/D VGND VGND VPWR VPWR _35013_/Q sky130_fd_sc_hd__dfxtp_1
X_32225_ _35715_/CLK _32225_/D VGND VGND VPWR VPWR _32225_/Q sky130_fd_sc_hd__dfxtp_1
Xinput74 R2[3] VGND VGND VPWR VPWR input74/X sky130_fd_sc_hd__buf_4
XFILLER_200_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17159_ _34420_/Q _36148_/Q _34292_/Q _34228_/Q _16876_/X _16877_/X VGND VGND VPWR
+ VPWR _17159_/X sky130_fd_sc_hd__mux4_1
Xinput85 RW[2] VGND VGND VPWR VPWR input85/X sky130_fd_sc_hd__clkbuf_4
XFILLER_7_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20170_ _20164_/X _20165_/X _20168_/X _20169_/X VGND VGND VPWR VPWR _20170_/X sky130_fd_sc_hd__a22o_1
X_32156_ _36223_/CLK _32156_/D VGND VGND VPWR VPWR _32156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31107_ _31107_/A VGND VGND VPWR VPWR _35778_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32087_ _35865_/CLK _32087_/D VGND VGND VPWR VPWR _32087_/Q sky130_fd_sc_hd__dfxtp_1
X_35915_ _35980_/CLK _35915_/D VGND VGND VPWR VPWR _35915_/Q sky130_fd_sc_hd__dfxtp_1
X_31038_ _31038_/A VGND VGND VPWR VPWR _35745_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_233_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35846_ _35847_/CLK _35846_/D VGND VGND VPWR VPWR _35846_/Q sky130_fd_sc_hd__dfxtp_1
X_23860_ _22909_/X _32477_/Q _23864_/S VGND VGND VPWR VPWR _23861_/A sky130_fd_sc_hd__mux2_1
XTAP_3709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_6_0__f_CLK clkbuf_5_0_0_CLK/X VGND VGND VPWR VPWR clkbuf_leaf_2_CLK/A sky130_fd_sc_hd__clkbuf_16
XFILLER_85_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22811_ _35219_/Q _35155_/Q _35091_/Q _32275_/Q _20692_/X _20694_/X VGND VGND VPWR
+ VPWR _22811_/X sky130_fd_sc_hd__mux4_1
X_35777_ _35777_/CLK _35777_/D VGND VGND VPWR VPWR _35777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23791_ _23791_/A VGND VGND VPWR VPWR _32381_/D sky130_fd_sc_hd__clkbuf_1
X_32989_ _35805_/CLK _32989_/D VGND VGND VPWR VPWR _32989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_253_CLK clkbuf_6_63__f_CLK/X VGND VGND VPWR VPWR _34179_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_16_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25530_ _24979_/X _33232_/Q _25532_/S VGND VGND VPWR VPWR _25531_/A sky130_fd_sc_hd__mux2_1
X_22742_ _22738_/X _22741_/X _22446_/X _22447_/X VGND VGND VPWR VPWR _22757_/B sky130_fd_sc_hd__o211a_2
X_34728_ _34920_/CLK _34728_/D VGND VGND VPWR VPWR _34728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25461_ _24877_/X _33199_/Q _25469_/S VGND VGND VPWR VPWR _25462_/A sky130_fd_sc_hd__mux2_1
X_22673_ _33935_/Q _33871_/Q _33807_/Q _36111_/Q _20662_/X _20664_/X VGND VGND VPWR
+ VPWR _22673_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34659_ _36197_/CLK _34659_/D VGND VGND VPWR VPWR _34659_/Q sky130_fd_sc_hd__dfxtp_1
X_27200_ _33995_/Q _27199_/X _27218_/S VGND VGND VPWR VPWR _27201_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24412_ _24412_/A VGND VGND VPWR VPWR _32735_/D sky130_fd_sc_hd__clkbuf_1
X_21624_ _22450_/A VGND VGND VPWR VPWR _21624_/X sky130_fd_sc_hd__buf_4
X_28180_ _28180_/A VGND VGND VPWR VPWR _34422_/D sky130_fd_sc_hd__clkbuf_1
X_25392_ _25392_/A VGND VGND VPWR VPWR _33167_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27131_ input25/X VGND VGND VPWR VPWR _27131_/X sky130_fd_sc_hd__buf_2
XFILLER_138_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24343_ _24343_/A VGND VGND VPWR VPWR _32702_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21555_ _21453_/X _21553_/X _21554_/X _21456_/X VGND VGND VPWR VPWR _21555_/X sky130_fd_sc_hd__a22o_1
XFILLER_193_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20506_ _35475_/Q _35411_/Q _35347_/Q _35283_/Q _20260_/X _20261_/X VGND VGND VPWR
+ VPWR _20506_/X sky130_fd_sc_hd__mux4_1
XFILLER_166_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27062_ input64/X VGND VGND VPWR VPWR _27062_/X sky130_fd_sc_hd__buf_4
XFILLER_148_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24274_ _22912_/X _32670_/Q _24276_/S VGND VGND VPWR VPWR _24275_/A sky130_fd_sc_hd__mux2_1
X_21486_ _21446_/X _21484_/X _21485_/X _21451_/X VGND VGND VPWR VPWR _21486_/X sky130_fd_sc_hd__a22o_1
XFILLER_181_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26013_ _26013_/A VGND VGND VPWR VPWR _33460_/D sky130_fd_sc_hd__clkbuf_1
X_23225_ input1/X VGND VGND VPWR VPWR _23225_/X sky130_fd_sc_hd__buf_4
XFILLER_165_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20437_ _33169_/Q _36049_/Q _33041_/Q _32977_/Q _18332_/X _19461_/A VGND VGND VPWR
+ VPWR _20437_/X sky130_fd_sc_hd__mux4_1
XFILLER_10_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20368_ _20368_/A VGND VGND VPWR VPWR _32462_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_161_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23156_ _23156_/A VGND VGND VPWR VPWR _32116_/D sky130_fd_sc_hd__clkbuf_1
XTAP_7036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22107_ _34686_/Q _34622_/Q _34558_/Q _34494_/Q _21892_/X _21893_/X VGND VGND VPWR
+ VPWR _22107_/X sky130_fd_sc_hd__mux4_1
XTAP_7069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27964_ _27964_/A VGND VGND VPWR VPWR _34320_/D sky130_fd_sc_hd__clkbuf_1
X_23087_ input85/X VGND VGND VPWR VPWR _27232_/B sky130_fd_sc_hd__buf_2
XFILLER_121_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20299_ _20299_/A VGND VGND VPWR VPWR _20299_/X sky130_fd_sc_hd__buf_4
XFILLER_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26915_ _26915_/A VGND VGND VPWR VPWR _33885_/D sky130_fd_sc_hd__clkbuf_1
X_29703_ _35113_/Q _29388_/X _29703_/S VGND VGND VPWR VPWR _29704_/A sky130_fd_sc_hd__mux2_1
X_22038_ _21753_/X _22036_/X _22037_/X _21756_/X VGND VGND VPWR VPWR _22038_/X sky130_fd_sc_hd__a22o_1
XTAP_6379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27895_ _27895_/A VGND VGND VPWR VPWR _34287_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_216_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_1127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_492_CLK clkbuf_6_3__f_CLK/X VGND VGND VPWR VPWR _35367_/CLK sky130_fd_sc_hd__clkbuf_16
X_29634_ _35080_/Q _29484_/X _29652_/S VGND VGND VPWR VPWR _29635_/A sky130_fd_sc_hd__mux2_1
XTAP_5678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26846_ _33853_/Q _23417_/X _26846_/S VGND VGND VPWR VPWR _26847_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_1330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_559 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29565_ _29565_/A VGND VGND VPWR VPWR _35047_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26777_ _33820_/Q _23249_/X _26783_/S VGND VGND VPWR VPWR _26778_/A sky130_fd_sc_hd__mux2_1
X_23989_ _23989_/A VGND VGND VPWR VPWR _32537_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_244_CLK clkbuf_6_61__f_CLK/X VGND VGND VPWR VPWR _36106_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_232_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28516_ _28648_/S VGND VGND VPWR VPWR _28535_/S sky130_fd_sc_hd__clkbuf_8
X_16530_ _16530_/A VGND VGND VPWR VPWR _31970_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25728_ _25728_/A VGND VGND VPWR VPWR _33325_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29496_ _29496_/A VGND VGND VPWR VPWR _35019_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28447_ _27739_/X _34549_/Q _28463_/S VGND VGND VPWR VPWR _28448_/A sky130_fd_sc_hd__mux2_1
X_16461_ _16461_/A _16461_/B _16461_/C _16461_/D VGND VGND VPWR VPWR _16462_/A sky130_fd_sc_hd__or4_4
X_25659_ _24970_/X _33293_/Q _25667_/S VGND VGND VPWR VPWR _25660_/A sky130_fd_sc_hd__mux2_1
XFILLER_189_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18200_ _32915_/Q _32851_/Q _32787_/Q _32723_/Q _15984_/X _15987_/X VGND VGND VPWR
+ VPWR _18200_/X sky130_fd_sc_hd__mux4_1
XFILLER_223_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19180_ _19105_/X _19178_/X _19179_/X _19110_/X VGND VGND VPWR VPWR _19180_/X sky130_fd_sc_hd__a22o_1
XPHY_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28378_ _27837_/X _34517_/Q _28378_/S VGND VGND VPWR VPWR _28379_/A sky130_fd_sc_hd__mux2_1
X_16392_ _33887_/Q _33823_/Q _33759_/Q _36063_/Q _16318_/X _16319_/X VGND VGND VPWR
+ VPWR _16392_/X sky130_fd_sc_hd__mux4_1
XPHY_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18131_ _17905_/X _18129_/X _18130_/X _17910_/X VGND VGND VPWR VPWR _18131_/X sky130_fd_sc_hd__a22o_1
XPHY_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27329_ _27329_/A VGND VGND VPWR VPWR _34050_/D sky130_fd_sc_hd__clkbuf_1
XPHY_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30340_ _30340_/A VGND VGND VPWR VPWR _35414_/D sky130_fd_sc_hd__clkbuf_1
X_18062_ _17859_/X _18060_/X _18061_/X _17862_/X VGND VGND VPWR VPWR _18062_/X sky130_fd_sc_hd__a22o_1
XFILLER_106_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17013_ _16800_/X _17009_/X _17012_/X _16803_/X VGND VGND VPWR VPWR _17013_/X sky130_fd_sc_hd__a22o_1
XFILLER_7_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30271_ _35382_/Q _29429_/X _30285_/S VGND VGND VPWR VPWR _30272_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32010_ _36202_/CLK _32010_/D VGND VGND VPWR VPWR _32010_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18964_ _18960_/X _18963_/X _18759_/X VGND VGND VPWR VPWR _18965_/D sky130_fd_sc_hd__o21ba_1
X_17915_ _17915_/A VGND VGND VPWR VPWR _17915_/X sky130_fd_sc_hd__buf_4
XFILLER_140_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33961_ _34153_/CLK _33961_/D VGND VGND VPWR VPWR _33961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_234_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18895_ _18895_/A _18895_/B _18895_/C _18895_/D VGND VGND VPWR VPWR _18896_/A sky130_fd_sc_hd__or4_2
XTAP_6880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35700_ _35701_/CLK _35700_/D VGND VGND VPWR VPWR _35700_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_483_CLK _35560_/CLK VGND VGND VPWR VPWR _33895_/CLK sky130_fd_sc_hd__clkbuf_16
X_32912_ _32913_/CLK _32912_/D VGND VGND VPWR VPWR _32912_/Q sky130_fd_sc_hd__dfxtp_1
X_17846_ _17846_/A VGND VGND VPWR VPWR _17846_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_66_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33892_ _36070_/CLK _33892_/D VGND VGND VPWR VPWR _33892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35631_ _35632_/CLK _35631_/D VGND VGND VPWR VPWR _35631_/Q sky130_fd_sc_hd__dfxtp_1
X_32843_ _32907_/CLK _32843_/D VGND VGND VPWR VPWR _32843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17777_ _17777_/A VGND VGND VPWR VPWR _17777_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_19_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_235_CLK clkbuf_6_54__f_CLK/X VGND VGND VPWR VPWR _36167_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19516_ _32886_/Q _32822_/Q _32758_/Q _32694_/Q _19293_/X _19294_/X VGND VGND VPWR
+ VPWR _19516_/X sky130_fd_sc_hd__mux4_1
XFILLER_235_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35562_ _35691_/CLK _35562_/D VGND VGND VPWR VPWR _35562_/Q sky130_fd_sc_hd__dfxtp_1
X_16728_ _16650_/X _16724_/X _16727_/X _16653_/X VGND VGND VPWR VPWR _16728_/X sky130_fd_sc_hd__a22o_1
X_32774_ _32905_/CLK _32774_/D VGND VGND VPWR VPWR _32774_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34513_ _34705_/CLK _34513_/D VGND VGND VPWR VPWR _34513_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31725_ _36071_/Q input9/X _31729_/S VGND VGND VPWR VPWR _31726_/A sky130_fd_sc_hd__mux2_1
X_19447_ _19298_/X _19443_/X _19446_/X _19301_/X VGND VGND VPWR VPWR _19447_/X sky130_fd_sc_hd__a22o_1
X_16659_ _35174_/Q _35110_/Q _35046_/Q _32166_/Q _16657_/X _16658_/X VGND VGND VPWR
+ VPWR _16659_/X sky130_fd_sc_hd__mux4_1
XFILLER_224_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35493_ _35685_/CLK _35493_/D VGND VGND VPWR VPWR _35493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34444_ _36173_/CLK _34444_/D VGND VGND VPWR VPWR _34444_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31656_ _31656_/A VGND VGND VPWR VPWR _36038_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19378_ _20235_/A VGND VGND VPWR VPWR _19378_/X sky130_fd_sc_hd__buf_6
XFILLER_37_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30607_ _30877_/A _30607_/B VGND VGND VPWR VPWR _30740_/S sky130_fd_sc_hd__nor2_8
XFILLER_147_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18329_ _20073_/A VGND VGND VPWR VPWR _20212_/A sky130_fd_sc_hd__buf_12
X_34375_ _35717_/CLK _34375_/D VGND VGND VPWR VPWR _34375_/Q sky130_fd_sc_hd__dfxtp_1
X_31587_ _31587_/A VGND VGND VPWR VPWR _36005_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36114_ _36114_/CLK _36114_/D VGND VGND VPWR VPWR _36114_/Q sky130_fd_sc_hd__dfxtp_1
X_21340_ _22560_/A VGND VGND VPWR VPWR _21340_/X sky130_fd_sc_hd__buf_4
X_33326_ _36079_/CLK _33326_/D VGND VGND VPWR VPWR _33326_/Q sky130_fd_sc_hd__dfxtp_1
X_30538_ _30538_/A VGND VGND VPWR VPWR _35508_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36045_ _36045_/CLK _36045_/D VGND VGND VPWR VPWR _36045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21271_ _22450_/A VGND VGND VPWR VPWR _21271_/X sky130_fd_sc_hd__buf_4
XFILLER_190_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30469_ _30469_/A VGND VGND VPWR VPWR _35476_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33257_ _35622_/CLK _33257_/D VGND VGND VPWR VPWR _33257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20222_ _32906_/Q _32842_/Q _32778_/Q _32714_/Q _19999_/X _20000_/X VGND VGND VPWR
+ VPWR _20222_/X sky130_fd_sc_hd__mux4_1
X_23010_ _23010_/A VGND VGND VPWR VPWR _32061_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32208_ _35699_/CLK _32208_/D VGND VGND VPWR VPWR _32208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_235_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33188_ _33828_/CLK _33188_/D VGND VGND VPWR VPWR _33188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20153_ _20004_/X _20149_/X _20152_/X _20007_/X VGND VGND VPWR VPWR _20153_/X sky130_fd_sc_hd__a22o_1
X_32139_ _35980_/CLK _32139_/D VGND VGND VPWR VPWR _32139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24961_ input48/X VGND VGND VPWR VPWR _24961_/X sky130_fd_sc_hd__buf_4
X_20084_ _20235_/A VGND VGND VPWR VPWR _20084_/X sky130_fd_sc_hd__buf_6
XFILLER_58_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_474_CLK clkbuf_6_10__f_CLK/X VGND VGND VPWR VPWR _34991_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26700_ _26700_/A VGND VGND VPWR VPWR _33783_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23912_ _23912_/A VGND VGND VPWR VPWR _32501_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_213_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27680_ input4/X VGND VGND VPWR VPWR _27680_/X sky130_fd_sc_hd__buf_4
XFILLER_217_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24892_ input24/X VGND VGND VPWR VPWR _24892_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_57_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26631_ _26631_/A VGND VGND VPWR VPWR _33750_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_1160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23843_ _23843_/A VGND VGND VPWR VPWR _28380_/A sky130_fd_sc_hd__buf_6
XTAP_3539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35829_ _35829_/CLK _35829_/D VGND VGND VPWR VPWR _35829_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_226_CLK clkbuf_6_53__f_CLK/X VGND VGND VPWR VPWR _34440_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_246_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_226_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29350_ _29350_/A VGND VGND VPWR VPWR _34972_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26562_ _24905_/X _33720_/Q _26572_/S VGND VGND VPWR VPWR _26563_/A sky130_fd_sc_hd__mux2_1
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23774_ _22984_/X _32373_/Q _23790_/S VGND VGND VPWR VPWR _23775_/A sky130_fd_sc_hd__mux2_1
XFILLER_232_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20986_ _33631_/Q _33567_/Q _33503_/Q _33439_/Q _20741_/X _20742_/X VGND VGND VPWR
+ VPWR _20986_/X sky130_fd_sc_hd__mux4_1
X_28301_ _27723_/X _34480_/Q _28307_/S VGND VGND VPWR VPWR _28302_/A sky130_fd_sc_hd__mux2_1
X_25513_ _25540_/S VGND VGND VPWR VPWR _25532_/S sky130_fd_sc_hd__buf_4
X_22725_ _22464_/X _22723_/X _22724_/X _22469_/X VGND VGND VPWR VPWR _22725_/X sky130_fd_sc_hd__a22o_1
X_29281_ _34943_/Q _27162_/X _29297_/S VGND VGND VPWR VPWR _29282_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26493_ _24803_/X _33687_/Q _26509_/S VGND VGND VPWR VPWR _26494_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28232_ _28232_/A VGND VGND VPWR VPWR _34447_/D sky130_fd_sc_hd__clkbuf_1
X_25444_ _24852_/X _33191_/Q _25448_/S VGND VGND VPWR VPWR _25445_/A sky130_fd_sc_hd__mux2_1
XFILLER_198_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22656_ _35470_/Q _35406_/Q _35342_/Q _35278_/Q _22560_/X _22561_/X VGND VGND VPWR
+ VPWR _22656_/X sky130_fd_sc_hd__mux4_1
XFILLER_159_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28163_ _28163_/A VGND VGND VPWR VPWR _34414_/D sky130_fd_sc_hd__clkbuf_1
X_21607_ _21603_/X _21604_/X _21605_/X _21606_/X VGND VGND VPWR VPWR _21607_/X sky130_fd_sc_hd__a22o_1
X_25375_ _25375_/A VGND VGND VPWR VPWR _33159_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22587_ _32140_/Q _32332_/Q _32396_/Q _35916_/Q _22586_/X _22374_/X VGND VGND VPWR
+ VPWR _22587_/X sky130_fd_sc_hd__mux4_1
XFILLER_22_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27114_ _27114_/A VGND VGND VPWR VPWR _33967_/D sky130_fd_sc_hd__clkbuf_1
X_24326_ _24326_/A VGND VGND VPWR VPWR _32694_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28094_ _34382_/Q _27208_/X _28100_/S VGND VGND VPWR VPWR _28095_/A sky130_fd_sc_hd__mux2_1
X_21538_ _21534_/X _21537_/X _21398_/X VGND VGND VPWR VPWR _21548_/C sky130_fd_sc_hd__o21ba_1
XFILLER_194_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27045_ _33945_/Q _27044_/X _27063_/S VGND VGND VPWR VPWR _27046_/A sky130_fd_sc_hd__mux2_1
XFILLER_175_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24257_ _24389_/S VGND VGND VPWR VPWR _24276_/S sky130_fd_sc_hd__clkbuf_8
X_21469_ _35436_/Q _35372_/Q _35308_/Q _35244_/Q _21148_/X _21149_/X VGND VGND VPWR
+ VPWR _21469_/X sky130_fd_sc_hd__mux4_1
XFILLER_182_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23208_ _23208_/A VGND VGND VPWR VPWR _32141_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_1030 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24188_ _24188_/A VGND VGND VPWR VPWR _32630_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23139_ _23139_/A VGND VGND VPWR VPWR _32108_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28996_ _34808_/Q _27140_/X _29006_/S VGND VGND VPWR VPWR _28997_/A sky130_fd_sc_hd__mux2_1
XTAP_6143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27947_ _27797_/X _34312_/Q _27965_/S VGND VGND VPWR VPWR _27948_/A sky130_fd_sc_hd__mux2_1
XTAP_6165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17700_ _17834_/A VGND VGND VPWR VPWR _17700_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_465_CLK clkbuf_6_11__f_CLK/X VGND VGND VPWR VPWR _34924_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_236_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18680_ _34398_/Q _36126_/Q _34270_/Q _34206_/Q _18470_/X _18471_/X VGND VGND VPWR
+ VPWR _18680_/X sky130_fd_sc_hd__mux4_1
XTAP_4730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27878_ _27878_/A VGND VGND VPWR VPWR _34279_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29617_ _35072_/Q _29460_/X _29631_/S VGND VGND VPWR VPWR _29618_/A sky130_fd_sc_hd__mux2_1
XTAP_4763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17631_ _33154_/Q _36034_/Q _33026_/Q _32962_/Q _17415_/X _17416_/X VGND VGND VPWR
+ VPWR _17631_/X sky130_fd_sc_hd__mux4_1
XFILLER_91_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26829_ _26829_/A VGND VGND VPWR VPWR _33844_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_247_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_217_CLK clkbuf_6_52__f_CLK/X VGND VGND VPWR VPWR _35212_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17562_ _17915_/A VGND VGND VPWR VPWR _17562_/X sky130_fd_sc_hd__buf_4
XFILLER_217_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29548_ _29548_/A VGND VGND VPWR VPWR _35039_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_223_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19301_ _20162_/A VGND VGND VPWR VPWR _19301_/X sky130_fd_sc_hd__clkbuf_4
X_16513_ _35682_/Q _32189_/Q _35554_/Q _35490_/Q _16258_/X _16259_/X VGND VGND VPWR
+ VPWR _16513_/X sky130_fd_sc_hd__mux4_1
XFILLER_216_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17493_ _17846_/A VGND VGND VPWR VPWR _17493_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_17_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29479_ _35014_/Q _29478_/X _29482_/S VGND VGND VPWR VPWR _29480_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31510_ _27776_/X _35969_/Q _31522_/S VGND VGND VPWR VPWR _31511_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19232_ _35694_/Q _32202_/Q _35566_/Q _35502_/Q _18911_/X _18912_/X VGND VGND VPWR
+ VPWR _19232_/X sky130_fd_sc_hd__mux4_1
X_16444_ _16297_/X _16442_/X _16443_/X _16300_/X VGND VGND VPWR VPWR _16444_/X sky130_fd_sc_hd__a22o_1
XFILLER_177_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32490_ _36010_/CLK _32490_/D VGND VGND VPWR VPWR _32490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_779 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31441_ _27673_/X _35936_/Q _31459_/S VGND VGND VPWR VPWR _31442_/A sky130_fd_sc_hd__mux2_1
X_19163_ _32876_/Q _32812_/Q _32748_/Q _32684_/Q _18940_/X _18941_/X VGND VGND VPWR
+ VPWR _19163_/X sky130_fd_sc_hd__mux4_1
XFILLER_9_920 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_943 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16375_ _16297_/X _16371_/X _16374_/X _16300_/X VGND VGND VPWR VPWR _16375_/X sky130_fd_sc_hd__a22o_1
XFILLER_157_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18114_ _35664_/Q _35024_/Q _34384_/Q _33744_/Q _17850_/X _17851_/X VGND VGND VPWR
+ VPWR _18114_/X sky130_fd_sc_hd__mux4_1
XFILLER_160_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34160_ _35632_/CLK _34160_/D VGND VGND VPWR VPWR _34160_/Q sky130_fd_sc_hd__dfxtp_1
X_31372_ _31372_/A VGND VGND VPWR VPWR _35903_/D sky130_fd_sc_hd__clkbuf_1
X_19094_ _18945_/X _19090_/X _19093_/X _18948_/X VGND VGND VPWR VPWR _19094_/X sky130_fd_sc_hd__a22o_1
XFILLER_219_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_986 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18045_ _18041_/X _18044_/X _17838_/X VGND VGND VPWR VPWR _18067_/A sky130_fd_sc_hd__o21ba_2
X_33111_ _35993_/CLK _33111_/D VGND VGND VPWR VPWR _33111_/Q sky130_fd_sc_hd__dfxtp_1
X_30323_ _35407_/Q _29506_/X _30327_/S VGND VGND VPWR VPWR _30324_/A sky130_fd_sc_hd__mux2_1
X_34091_ _34091_/CLK _34091_/D VGND VGND VPWR VPWR _34091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33042_ _35858_/CLK _33042_/D VGND VGND VPWR VPWR _33042_/Q sky130_fd_sc_hd__dfxtp_1
X_30254_ _35374_/Q _29404_/X _30264_/S VGND VGND VPWR VPWR _30255_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30185_ _30185_/A VGND VGND VPWR VPWR _35341_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19996_ _33156_/Q _36036_/Q _33028_/Q _32964_/Q _19715_/X _19716_/X VGND VGND VPWR
+ VPWR _19996_/X sky130_fd_sc_hd__mux4_1
XFILLER_99_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18947_ _35622_/Q _34982_/Q _34342_/Q _33702_/Q _18738_/X _18739_/X VGND VGND VPWR
+ VPWR _18947_/X sky130_fd_sc_hd__mux4_1
XFILLER_45_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_6_13__f_CLK clkbuf_5_6_0_CLK/X VGND VGND VPWR VPWR clkbuf_leaf_57_CLK/A sky130_fd_sc_hd__clkbuf_16
X_34993_ _35567_/CLK _34993_/D VGND VGND VPWR VPWR _34993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_1344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_456_CLK clkbuf_6_14__f_CLK/X VGND VGND VPWR VPWR _36010_/CLK sky130_fd_sc_hd__clkbuf_16
X_33944_ _35610_/CLK _33944_/D VGND VGND VPWR VPWR _33944_/Q sky130_fd_sc_hd__dfxtp_1
X_18878_ _18873_/X _18877_/X _18734_/X _18735_/X VGND VGND VPWR VPWR _18895_/B sky130_fd_sc_hd__o211a_1
XFILLER_95_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17829_ _17829_/A VGND VGND VPWR VPWR _32007_/D sky130_fd_sc_hd__buf_4
XFILLER_54_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33875_ _33875_/CLK _33875_/D VGND VGND VPWR VPWR _33875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_212_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_208_CLK clkbuf_6_54__f_CLK/X VGND VGND VPWR VPWR _34633_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_54_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35614_ _35615_/CLK _35614_/D VGND VGND VPWR VPWR _35614_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_242_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20840_ _20691_/X _20838_/X _20839_/X _20701_/X VGND VGND VPWR VPWR _20840_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32826_ _32890_/CLK _32826_/D VGND VGND VPWR VPWR _32826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35545_ _35609_/CLK _35545_/D VGND VGND VPWR VPWR _35545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20771_ _21477_/A VGND VGND VPWR VPWR _20771_/X sky130_fd_sc_hd__buf_6
X_32757_ _32885_/CLK _32757_/D VGND VGND VPWR VPWR _32757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_1418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22510_ _22510_/A VGND VGND VPWR VPWR _22510_/X sky130_fd_sc_hd__buf_4
XFILLER_168_718 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31708_ _36063_/Q input64/X _31708_/S VGND VGND VPWR VPWR _31709_/A sky130_fd_sc_hd__mux2_1
X_35476_ _35860_/CLK _35476_/D VGND VGND VPWR VPWR _35476_/Q sky130_fd_sc_hd__dfxtp_1
X_23490_ _32242_/Q _23393_/X _23515_/S VGND VGND VPWR VPWR _23491_/A sky130_fd_sc_hd__mux2_1
X_32688_ _32879_/CLK _32688_/D VGND VGND VPWR VPWR _32688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22441_ _33160_/Q _36040_/Q _33032_/Q _32968_/Q _22368_/X _22369_/X VGND VGND VPWR
+ VPWR _22441_/X sky130_fd_sc_hd__mux4_1
X_34427_ _36157_/CLK _34427_/D VGND VGND VPWR VPWR _34427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31639_ _27766_/X _36030_/Q _31657_/S VGND VGND VPWR VPWR _31640_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25160_ _25160_/A VGND VGND VPWR VPWR _33057_/D sky130_fd_sc_hd__clkbuf_1
X_22372_ _22365_/X _22367_/X _22370_/X _22371_/X VGND VGND VPWR VPWR _22372_/X sky130_fd_sc_hd__a22o_1
X_34358_ _35830_/CLK _34358_/D VGND VGND VPWR VPWR _34358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24111_ _23079_/X _32596_/Q _24113_/S VGND VGND VPWR VPWR _24112_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33309_ _36060_/CLK _33309_/D VGND VGND VPWR VPWR _33309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21323_ _21245_/X _21321_/X _21322_/X _21248_/X VGND VGND VPWR VPWR _21323_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25091_ _24936_/X _33026_/Q _25101_/S VGND VGND VPWR VPWR _25092_/A sky130_fd_sc_hd__mux2_1
X_34289_ _36144_/CLK _34289_/D VGND VGND VPWR VPWR _34289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_873 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21254_ _21250_/X _21251_/X _21252_/X _21253_/X VGND VGND VPWR VPWR _21254_/X sky130_fd_sc_hd__a22o_1
X_24042_ _22977_/X _32563_/Q _24042_/S VGND VGND VPWR VPWR _24043_/A sky130_fd_sc_hd__mux2_1
X_36028_ _36029_/CLK _36028_/D VGND VGND VPWR VPWR _36028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20205_ _20205_/A VGND VGND VPWR VPWR _20205_/X sky130_fd_sc_hd__buf_4
XFILLER_176_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28850_ _34739_/Q _27124_/X _28850_/S VGND VGND VPWR VPWR _28851_/A sky130_fd_sc_hd__mux2_1
X_21185_ _21181_/X _21184_/X _21045_/X VGND VGND VPWR VPWR _21195_/C sky130_fd_sc_hd__o21ba_1
XFILLER_143_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20136_ _33928_/Q _33864_/Q _33800_/Q _36104_/Q _20030_/X _20031_/X VGND VGND VPWR
+ VPWR _20136_/X sky130_fd_sc_hd__mux4_1
X_27801_ input47/X VGND VGND VPWR VPWR _27801_/X sky130_fd_sc_hd__clkbuf_4
X_28781_ _28781_/A VGND VGND VPWR VPWR _34707_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25993_ _24865_/X _33451_/Q _26009_/S VGND VGND VPWR VPWR _25994_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_447_CLK clkbuf_leaf_61_CLK/A VGND VGND VPWR VPWR _35949_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_225_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27732_ input22/X VGND VGND VPWR VPWR _27732_/X sky130_fd_sc_hd__buf_2
XFILLER_86_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24944_ _24944_/A VGND VGND VPWR VPWR _32964_/D sky130_fd_sc_hd__clkbuf_1
X_20067_ _32646_/Q _32582_/Q _32518_/Q _35974_/Q _19929_/X _20066_/X VGND VGND VPWR
+ VPWR _20067_/X sky130_fd_sc_hd__mux4_1
XTAP_4015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_906 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27663_ _27663_/A VGND VGND VPWR VPWR _34204_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24875_ _24874_/X _32942_/Q _24890_/S VGND VGND VPWR VPWR _24876_/A sky130_fd_sc_hd__mux2_1
XTAP_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26614_ _24982_/X _33745_/Q _26614_/S VGND VGND VPWR VPWR _26615_/A sky130_fd_sc_hd__mux2_1
X_29402_ _34989_/Q _29401_/X _29420_/S VGND VGND VPWR VPWR _29403_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23826_ _23061_/X _32398_/Q _23832_/S VGND VGND VPWR VPWR _23827_/A sky130_fd_sc_hd__mux2_1
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27594_ _34176_/Q _27165_/X _27608_/S VGND VGND VPWR VPWR _27595_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29333_ input12/X VGND VGND VPWR VPWR _29333_/X sky130_fd_sc_hd__buf_2
X_26545_ _24880_/X _33712_/Q _26551_/S VGND VGND VPWR VPWR _26546_/A sky130_fd_sc_hd__mux2_1
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23757_ _22959_/X _32365_/Q _23769_/S VGND VGND VPWR VPWR _23758_/A sky130_fd_sc_hd__mux2_1
XFILLER_202_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20969_ _35614_/Q _34974_/Q _34334_/Q _33694_/Q _20653_/X _20655_/X VGND VGND VPWR
+ VPWR _20969_/X sky130_fd_sc_hd__mux4_1
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22708_ _21753_/A _22706_/X _22707_/X _21756_/A VGND VGND VPWR VPWR _22708_/X sky130_fd_sc_hd__a22o_1
X_29264_ _34935_/Q _27137_/X _29276_/S VGND VGND VPWR VPWR _29265_/A sky130_fd_sc_hd__mux2_1
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26476_ _33680_/Q _23481_/X _26478_/S VGND VGND VPWR VPWR _26477_/A sky130_fd_sc_hd__mux2_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23688_ _23061_/X _32334_/Q _23694_/S VGND VGND VPWR VPWR _23689_/A sky130_fd_sc_hd__mux2_1
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28215_ _28215_/A VGND VGND VPWR VPWR _34439_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25427_ _24827_/X _33183_/Q _25427_/S VGND VGND VPWR VPWR _25428_/A sky130_fd_sc_hd__mux2_1
X_29195_ _34902_/Q _27033_/X _29213_/S VGND VGND VPWR VPWR _29196_/A sky130_fd_sc_hd__mux2_1
X_22639_ _33678_/Q _33614_/Q _33550_/Q _33486_/Q _22506_/X _22507_/X VGND VGND VPWR
+ VPWR _22639_/X sky130_fd_sc_hd__mux4_1
XFILLER_201_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16160_ _35672_/Q _32178_/Q _35544_/Q _35480_/Q _16049_/X _16050_/X VGND VGND VPWR
+ VPWR _16160_/X sky130_fd_sc_hd__mux4_1
XFILLER_167_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28146_ _28146_/A VGND VGND VPWR VPWR _34406_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25358_ _33151_/Q _23426_/X _25374_/S VGND VGND VPWR VPWR _25359_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24309_ _24309_/A VGND VGND VPWR VPWR _32686_/D sky130_fd_sc_hd__clkbuf_1
X_16091_ _17158_/A VGND VGND VPWR VPWR _16091_/X sky130_fd_sc_hd__clkbuf_4
X_28077_ _34374_/Q _27183_/X _28079_/S VGND VGND VPWR VPWR _28078_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25289_ _25289_/A VGND VGND VPWR VPWR _33118_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_1136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27028_ _27028_/A VGND VGND VPWR VPWR _33939_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_1450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19850_ _19850_/A _19850_/B _19850_/C _19850_/D VGND VGND VPWR VPWR _19851_/A sky130_fd_sc_hd__or4_4
XFILLER_64_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18801_ _33378_/Q _33314_/Q _33250_/Q _33186_/Q _18721_/X _18722_/X VGND VGND VPWR
+ VPWR _18801_/X sky130_fd_sc_hd__mux4_1
X_19781_ _20134_/A VGND VGND VPWR VPWR _19781_/X sky130_fd_sc_hd__buf_4
X_28979_ _34800_/Q _27115_/X _28985_/S VGND VGND VPWR VPWR _28980_/A sky130_fd_sc_hd__mux2_1
X_16993_ _17833_/A VGND VGND VPWR VPWR _16993_/X sky130_fd_sc_hd__buf_4
XFILLER_0_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_438_CLK clkbuf_6_36__f_CLK/X VGND VGND VPWR VPWR _36016_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_231_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18732_ _32864_/Q _32800_/Q _32736_/Q _32672_/Q _18587_/X _18588_/X VGND VGND VPWR
+ VPWR _18732_/X sky130_fd_sc_hd__mux4_1
XFILLER_209_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31990_ _34914_/CLK _31990_/D VGND VGND VPWR VPWR _31990_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_974 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18663_ _32094_/Q _32286_/Q _32350_/Q _35870_/Q _18521_/X _18662_/X VGND VGND VPWR
+ VPWR _18663_/X sky130_fd_sc_hd__mux4_1
X_30941_ _31010_/S VGND VGND VPWR VPWR _30960_/S sky130_fd_sc_hd__buf_6
XFILLER_188_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17614_ _35201_/Q _35137_/Q _35073_/Q _32257_/Q _17363_/X _17364_/X VGND VGND VPWR
+ VPWR _17614_/X sky130_fd_sc_hd__mux4_1
XTAP_4593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33660_ _33661_/CLK _33660_/D VGND VGND VPWR VPWR _33660_/Q sky130_fd_sc_hd__dfxtp_1
X_30872_ _30872_/A VGND VGND VPWR VPWR _35667_/D sky130_fd_sc_hd__clkbuf_1
X_18594_ _35612_/Q _34972_/Q _34332_/Q _33692_/Q _18353_/X _18355_/X VGND VGND VPWR
+ VPWR _18594_/X sky130_fd_sc_hd__mux4_1
XFILLER_52_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32611_ _35938_/CLK _32611_/D VGND VGND VPWR VPWR _32611_/Q sky130_fd_sc_hd__dfxtp_1
X_17545_ _17506_/X _17543_/X _17544_/X _17509_/X VGND VGND VPWR VPWR _17545_/X sky130_fd_sc_hd__a22o_1
X_33591_ _33850_/CLK _33591_/D VGND VGND VPWR VPWR _33591_/Q sky130_fd_sc_hd__dfxtp_1
X_35330_ _35458_/CLK _35330_/D VGND VGND VPWR VPWR _35330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32542_ _35998_/CLK _32542_/D VGND VGND VPWR VPWR _32542_/Q sky130_fd_sc_hd__dfxtp_1
X_17476_ _17476_/A VGND VGND VPWR VPWR _31997_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19215_ _19215_/A VGND VGND VPWR VPWR _32429_/D sky130_fd_sc_hd__clkbuf_1
X_16427_ _16420_/X _16425_/X _16426_/X VGND VGND VPWR VPWR _16461_/A sky130_fd_sc_hd__o21ba_1
X_35261_ _36029_/CLK _35261_/D VGND VGND VPWR VPWR _35261_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_242_1462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32473_ _35929_/CLK _32473_/D VGND VGND VPWR VPWR _32473_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34212_ _34405_/CLK _34212_/D VGND VGND VPWR VPWR _34212_/Q sky130_fd_sc_hd__dfxtp_1
X_31424_ _27649_/X _35928_/Q _31438_/S VGND VGND VPWR VPWR _31425_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16358_ _33118_/Q _35998_/Q _32990_/Q _32926_/Q _16356_/X _16357_/X VGND VGND VPWR
+ VPWR _16358_/X sky130_fd_sc_hd__mux4_1
XFILLER_125_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19146_ _20205_/A VGND VGND VPWR VPWR _19146_/X sky130_fd_sc_hd__clkbuf_4
X_35192_ _35192_/CLK _35192_/D VGND VGND VPWR VPWR _35192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34143_ _36188_/CLK _34143_/D VGND VGND VPWR VPWR _34143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31355_ _31355_/A VGND VGND VPWR VPWR _35895_/D sky130_fd_sc_hd__clkbuf_1
X_16289_ _32860_/Q _32796_/Q _32732_/Q _32668_/Q _16287_/X _16288_/X VGND VGND VPWR
+ VPWR _16289_/X sky130_fd_sc_hd__mux4_1
X_19077_ _33898_/Q _33834_/Q _33770_/Q _36074_/Q _18971_/X _18972_/X VGND VGND VPWR
+ VPWR _19077_/X sky130_fd_sc_hd__mux4_1
XFILLER_172_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30306_ _35399_/Q _29481_/X _30306_/S VGND VGND VPWR VPWR _30307_/A sky130_fd_sc_hd__mux2_1
X_18028_ _17709_/X _18026_/X _18027_/X _17712_/X VGND VGND VPWR VPWR _18028_/X sky130_fd_sc_hd__a22o_1
XFILLER_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31286_ _31286_/A VGND VGND VPWR VPWR _35862_/D sky130_fd_sc_hd__clkbuf_1
X_34074_ _36219_/CLK _34074_/D VGND VGND VPWR VPWR _34074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33025_ _36033_/CLK _33025_/D VGND VGND VPWR VPWR _33025_/Q sky130_fd_sc_hd__dfxtp_1
X_30237_ _35366_/Q _29379_/X _30243_/S VGND VGND VPWR VPWR _30238_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1019 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30168_ _30168_/A VGND VGND VPWR VPWR _35333_/D sky130_fd_sc_hd__clkbuf_1
X_19979_ _34691_/Q _34627_/Q _34563_/Q _34499_/Q _19945_/X _19946_/X VGND VGND VPWR
+ VPWR _19979_/X sky130_fd_sc_hd__mux4_1
XFILLER_140_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_429_CLK clkbuf_6_38__f_CLK/X VGND VGND VPWR VPWR _34612_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_101_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22990_ input27/X VGND VGND VPWR VPWR _22990_/X sky130_fd_sc_hd__clkbuf_4
X_34976_ _35177_/CLK _34976_/D VGND VGND VPWR VPWR _34976_/Q sky130_fd_sc_hd__dfxtp_1
X_30099_ _30099_/A VGND VGND VPWR VPWR _35300_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_227_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33927_ _36159_/CLK _33927_/D VGND VGND VPWR VPWR _33927_/Q sky130_fd_sc_hd__dfxtp_1
X_21941_ _21937_/X _21940_/X _21732_/X VGND VGND VPWR VPWR _21971_/A sky130_fd_sc_hd__o21ba_1
XFILLER_55_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24660_ _24660_/A VGND VGND VPWR VPWR _32853_/D sky130_fd_sc_hd__clkbuf_1
X_33858_ _36099_/CLK _33858_/D VGND VGND VPWR VPWR _33858_/Q sky130_fd_sc_hd__dfxtp_1
X_21872_ _33400_/Q _33336_/Q _33272_/Q _33208_/Q _21727_/X _21728_/X VGND VGND VPWR
+ VPWR _21872_/X sky130_fd_sc_hd__mux4_1
XFILLER_242_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23611_ _23611_/A VGND VGND VPWR VPWR _32297_/D sky130_fd_sc_hd__clkbuf_1
X_20823_ _32858_/Q _32794_/Q _32730_/Q _32666_/Q _20637_/X _20639_/X VGND VGND VPWR
+ VPWR _20823_/X sky130_fd_sc_hd__mux4_1
X_32809_ _32875_/CLK _32809_/D VGND VGND VPWR VPWR _32809_/Q sky130_fd_sc_hd__dfxtp_1
X_24591_ _22980_/X _32820_/Q _24609_/S VGND VGND VPWR VPWR _24592_/A sky130_fd_sc_hd__mux2_1
X_33789_ _36093_/CLK _33789_/D VGND VGND VPWR VPWR _33789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26330_ _24964_/X _33611_/Q _26342_/S VGND VGND VPWR VPWR _26331_/A sky130_fd_sc_hd__mux2_1
X_23542_ _23542_/A VGND VGND VPWR VPWR _32265_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35528_ _35721_/CLK _35528_/D VGND VGND VPWR VPWR _35528_/Q sky130_fd_sc_hd__dfxtp_1
X_20754_ _33112_/Q _35992_/Q _32984_/Q _32920_/Q _20624_/X _20625_/X VGND VGND VPWR
+ VPWR _20754_/X sky130_fd_sc_hd__mux4_1
XFILLER_211_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26261_ _24861_/X _33578_/Q _26279_/S VGND VGND VPWR VPWR _26262_/A sky130_fd_sc_hd__mux2_1
X_23473_ _32236_/Q _23472_/X _23485_/S VGND VGND VPWR VPWR _23474_/A sky130_fd_sc_hd__mux2_1
X_35459_ _35841_/CLK _35459_/D VGND VGND VPWR VPWR _35459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20685_ _21611_/A VGND VGND VPWR VPWR _20685_/X sky130_fd_sc_hd__buf_4
XFILLER_210_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28000_ _34337_/Q _27069_/X _28016_/S VGND VGND VPWR VPWR _28001_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25212_ _25212_/A VGND VGND VPWR VPWR _33082_/D sky130_fd_sc_hd__clkbuf_1
X_22424_ _34439_/Q _36167_/Q _34311_/Q _34247_/Q _22182_/X _22183_/X VGND VGND VPWR
+ VPWR _22424_/X sky130_fd_sc_hd__mux4_1
X_26192_ _26192_/A VGND VGND VPWR VPWR _33545_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_1382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25143_ _25143_/A VGND VGND VPWR VPWR _33049_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22355_ _22351_/X _22354_/X _22118_/X VGND VGND VPWR VPWR _22356_/D sky130_fd_sc_hd__o21ba_1
XFILLER_163_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21306_ _22505_/A VGND VGND VPWR VPWR _21306_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_108_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29951_ _29951_/A VGND VGND VPWR VPWR _35230_/D sky130_fd_sc_hd__clkbuf_1
X_25074_ _24911_/X _33018_/Q _25080_/S VGND VGND VPWR VPWR _25075_/A sky130_fd_sc_hd__mux2_1
X_22286_ _22286_/A _22286_/B _22286_/C _22286_/D VGND VGND VPWR VPWR _22287_/A sky130_fd_sc_hd__or4_4
X_28902_ _28902_/A VGND VGND VPWR VPWR _34763_/D sky130_fd_sc_hd__clkbuf_1
X_24025_ _24025_/A VGND VGND VPWR VPWR _32554_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21237_ _33126_/Q _36006_/Q _32998_/Q _32934_/Q _20956_/X _20957_/X VGND VGND VPWR
+ VPWR _21237_/X sky130_fd_sc_hd__mux4_1
X_29882_ _29930_/S VGND VGND VPWR VPWR _29901_/S sky130_fd_sc_hd__buf_4
XFILLER_160_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28833_ _28833_/A VGND VGND VPWR VPWR _34730_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21168_ _21100_/X _21166_/X _21167_/X _21103_/X VGND VGND VPWR VPWR _21168_/X sky130_fd_sc_hd__a22o_1
XFILLER_78_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20119_ _20009_/X _20117_/X _20118_/X _20012_/X VGND VGND VPWR VPWR _20119_/X sky130_fd_sc_hd__a22o_1
X_28764_ _34699_/Q _27199_/X _28776_/S VGND VGND VPWR VPWR _28765_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21099_ _21093_/X _21096_/X _21097_/X _21098_/X VGND VGND VPWR VPWR _21099_/X sky130_fd_sc_hd__a22o_1
X_25976_ _24840_/X _33443_/Q _25988_/S VGND VGND VPWR VPWR _25977_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_10 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24927_ input36/X VGND VGND VPWR VPWR _24927_/X sky130_fd_sc_hd__clkbuf_4
X_27715_ _27714_/X _34221_/Q _27733_/S VGND VGND VPWR VPWR _27716_/A sky130_fd_sc_hd__mux2_1
XTAP_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28695_ _34666_/Q _27096_/X _28713_/S VGND VGND VPWR VPWR _28696_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_944 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27646_ input12/X VGND VGND VPWR VPWR _27646_/X sky130_fd_sc_hd__clkbuf_4
X_24858_ input11/X VGND VGND VPWR VPWR _24858_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23809_ _23036_/X _32390_/Q _23811_/S VGND VGND VPWR VPWR _23810_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27577_ _34168_/Q _27140_/X _27587_/S VGND VGND VPWR VPWR _27578_/A sky130_fd_sc_hd__mux2_1
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24789_ _24789_/A VGND VGND VPWR VPWR _32914_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17330_ _34937_/Q _34873_/Q _34809_/Q _34745_/Q _17160_/X _17161_/X VGND VGND VPWR
+ VPWR _17330_/X sky130_fd_sc_hd__mux4_1
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29316_ _34960_/Q _27214_/X _29318_/S VGND VGND VPWR VPWR _29317_/A sky130_fd_sc_hd__mux2_1
XFILLER_202_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26528_ _24855_/X _33704_/Q _26530_/S VGND VGND VPWR VPWR _26529_/A sky130_fd_sc_hd__mux2_1
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17261_ _35191_/Q _35127_/Q _35063_/Q _32247_/Q _17010_/X _17011_/X VGND VGND VPWR
+ VPWR _17261_/X sky130_fd_sc_hd__mux4_1
XFILLER_70_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26459_ _26486_/S VGND VGND VPWR VPWR _26478_/S sky130_fd_sc_hd__buf_4
XFILLER_198_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29247_ _34927_/Q _27112_/X _29255_/S VGND VGND VPWR VPWR _29248_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16212_ _16140_/X _16210_/X _16211_/X _16145_/X VGND VGND VPWR VPWR _16212_/X sky130_fd_sc_hd__a22o_1
X_19000_ _34152_/Q _34088_/Q _34024_/Q _33960_/Q _18687_/X _18688_/X VGND VGND VPWR
+ VPWR _19000_/X sky130_fd_sc_hd__mux4_2
XFILLER_186_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29178_ _29178_/A VGND VGND VPWR VPWR _34894_/D sky130_fd_sc_hd__clkbuf_1
X_17192_ _17153_/X _17190_/X _17191_/X _17156_/X VGND VGND VPWR VPWR _17192_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28129_ _28129_/A VGND VGND VPWR VPWR _34398_/D sky130_fd_sc_hd__clkbuf_1
X_16143_ _33624_/Q _33560_/Q _33496_/Q _33432_/Q _16141_/X _16142_/X VGND VGND VPWR
+ VPWR _16143_/X sky130_fd_sc_hd__mux4_1
XFILLER_10_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31140_ _31140_/A VGND VGND VPWR VPWR _35794_/D sky130_fd_sc_hd__clkbuf_1
X_16074_ input69/X input70/X VGND VGND VPWR VPWR _17857_/A sky130_fd_sc_hd__or2_4
XFILLER_170_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19902_ _19720_/X _19900_/X _19901_/X _19724_/X VGND VGND VPWR VPWR _19902_/X sky130_fd_sc_hd__a22o_1
XFILLER_114_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31071_ _31071_/A VGND VGND VPWR VPWR _35761_/D sky130_fd_sc_hd__clkbuf_1
X_30022_ _35264_/Q _29460_/X _30036_/S VGND VGND VPWR VPWR _30023_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19833_ _32895_/Q _32831_/Q _32767_/Q _32703_/Q _19646_/X _19647_/X VGND VGND VPWR
+ VPWR _19833_/X sky130_fd_sc_hd__mux4_1
XFILLER_64_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34830_ _34961_/CLK _34830_/D VGND VGND VPWR VPWR _34830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_1188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19764_ _35453_/Q _35389_/Q _35325_/Q _35261_/Q _19554_/X _19555_/X VGND VGND VPWR
+ VPWR _19764_/X sky130_fd_sc_hd__mux4_1
XFILLER_111_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16976_ _34415_/Q _36143_/Q _34287_/Q _34223_/Q _16876_/X _16877_/X VGND VGND VPWR
+ VPWR _16976_/X sky130_fd_sc_hd__mux4_1
X_18715_ _18711_/X _18714_/X _18404_/X VGND VGND VPWR VPWR _18716_/D sky130_fd_sc_hd__o21ba_2
XFILLER_37_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34761_ _34957_/CLK _34761_/D VGND VGND VPWR VPWR _34761_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput6 DW[14] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__buf_6
XTAP_5091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31973_ _34085_/CLK _31973_/D VGND VGND VPWR VPWR _31973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19695_ _19691_/X _19694_/X _19451_/X VGND VGND VPWR VPWR _19703_/C sky130_fd_sc_hd__o21ba_1
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33712_ _35439_/CLK _33712_/D VGND VGND VPWR VPWR _33712_/Q sky130_fd_sc_hd__dfxtp_1
X_18646_ _33630_/Q _33566_/Q _33502_/Q _33438_/Q _18441_/X _18442_/X VGND VGND VPWR
+ VPWR _18646_/X sky130_fd_sc_hd__mux4_1
XFILLER_25_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30924_ _30924_/A VGND VGND VPWR VPWR _35691_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_224_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34692_ _36164_/CLK _34692_/D VGND VGND VPWR VPWR _34692_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33643_ _34091_/CLK _33643_/D VGND VGND VPWR VPWR _33643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30855_ _35659_/Q input49/X _30867_/S VGND VGND VPWR VPWR _30856_/A sky130_fd_sc_hd__mux2_1
X_18577_ _34140_/Q _34076_/Q _34012_/Q _33948_/Q _18309_/X _18311_/X VGND VGND VPWR
+ VPWR _18577_/X sky130_fd_sc_hd__mux4_1
XFILLER_91_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17528_ _17524_/X _17527_/X _17485_/X VGND VGND VPWR VPWR _17550_/A sky130_fd_sc_hd__o21ba_1
XFILLER_162_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33574_ _34146_/CLK _33574_/D VGND VGND VPWR VPWR _33574_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30786_ _35626_/Q input13/X _30804_/S VGND VGND VPWR VPWR _30787_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35313_ _35377_/CLK _35313_/D VGND VGND VPWR VPWR _35313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32525_ _35983_/CLK _32525_/D VGND VGND VPWR VPWR _32525_/Q sky130_fd_sc_hd__dfxtp_1
X_17459_ _17420_/X _17457_/X _17458_/X _17424_/X VGND VGND VPWR VPWR _17459_/X sky130_fd_sc_hd__a22o_1
XFILLER_20_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35244_ _35691_/CLK _35244_/D VGND VGND VPWR VPWR _35244_/Q sky130_fd_sc_hd__dfxtp_1
X_20470_ _32914_/Q _32850_/Q _32786_/Q _32722_/Q _18284_/X _18287_/X VGND VGND VPWR
+ VPWR _20470_/X sky130_fd_sc_hd__mux4_1
X_32456_ _36076_/CLK _32456_/D VGND VGND VPWR VPWR _32456_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31407_ _31407_/A VGND VGND VPWR VPWR _35920_/D sky130_fd_sc_hd__clkbuf_1
X_19129_ _19125_/X _19128_/X _19087_/X _19088_/X VGND VGND VPWR VPWR _19144_/B sky130_fd_sc_hd__o211a_1
XFILLER_146_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35175_ _35365_/CLK _35175_/D VGND VGND VPWR VPWR _35175_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32387_ _35907_/CLK _32387_/D VGND VGND VPWR VPWR _32387_/Q sky130_fd_sc_hd__dfxtp_1
X_34126_ _34192_/CLK _34126_/D VGND VGND VPWR VPWR _34126_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22140_ _33087_/Q _32063_/Q _35839_/Q _35775_/Q _22031_/X _22032_/X VGND VGND VPWR
+ VPWR _22140_/X sky130_fd_sc_hd__mux4_1
XFILLER_173_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31338_ _31338_/A VGND VGND VPWR VPWR _35887_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34057_ _34121_/CLK _34057_/D VGND VGND VPWR VPWR _34057_/Q sky130_fd_sc_hd__dfxtp_1
X_22071_ _34429_/Q _36157_/Q _34301_/Q _34237_/Q _21829_/X _21830_/X VGND VGND VPWR
+ VPWR _22071_/X sky130_fd_sc_hd__mux4_1
XFILLER_82_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31269_ _27819_/X _35855_/Q _31273_/S VGND VGND VPWR VPWR _31270_/A sky130_fd_sc_hd__mux2_1
X_21022_ _22400_/A VGND VGND VPWR VPWR _21022_/X sky130_fd_sc_hd__buf_4
X_33008_ _36016_/CLK _33008_/D VGND VGND VPWR VPWR _33008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25830_ _24824_/X _33374_/Q _25832_/S VGND VGND VPWR VPWR _25831_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25761_ _25761_/A VGND VGND VPWR VPWR _33341_/D sky130_fd_sc_hd__clkbuf_1
X_34959_ _34961_/CLK _34959_/D VGND VGND VPWR VPWR _34959_/Q sky130_fd_sc_hd__dfxtp_1
X_22973_ _22973_/A VGND VGND VPWR VPWR _32049_/D sky130_fd_sc_hd__clkbuf_1
X_27500_ _34132_/Q _27226_/X _27502_/S VGND VGND VPWR VPWR _27501_/A sky130_fd_sc_hd__mux2_1
X_24712_ _24712_/A VGND VGND VPWR VPWR _32877_/D sky130_fd_sc_hd__clkbuf_1
X_28480_ _27788_/X _34565_/Q _28484_/S VGND VGND VPWR VPWR _28481_/A sky130_fd_sc_hd__mux2_1
X_21924_ _21603_/X _21922_/X _21923_/X _21606_/X VGND VGND VPWR VPWR _21924_/X sky130_fd_sc_hd__a22o_1
X_25692_ _25692_/A VGND VGND VPWR VPWR _33308_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27431_ _34099_/Q _27124_/X _27431_/S VGND VGND VPWR VPWR _27432_/A sky130_fd_sc_hd__mux2_1
X_24643_ _23058_/X _32845_/Q _24651_/S VGND VGND VPWR VPWR _24644_/A sky130_fd_sc_hd__mux2_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21855_ _22561_/A VGND VGND VPWR VPWR _21855_/X sky130_fd_sc_hd__buf_4
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27362_ _27362_/A VGND VGND VPWR VPWR _34066_/D sky130_fd_sc_hd__clkbuf_1
X_20806_ _20691_/X _20804_/X _20805_/X _20701_/X VGND VGND VPWR VPWR _20806_/X sky130_fd_sc_hd__a22o_1
X_24574_ _22956_/X _32812_/Q _24588_/S VGND VGND VPWR VPWR _24575_/A sky130_fd_sc_hd__mux2_1
X_21786_ _35445_/Q _35381_/Q _35317_/Q _35253_/Q _21501_/X _21502_/X VGND VGND VPWR
+ VPWR _21786_/X sky130_fd_sc_hd__mux4_1
XFILLER_58_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26313_ _24939_/X _33603_/Q _26321_/S VGND VGND VPWR VPWR _26314_/A sky130_fd_sc_hd__mux2_1
XFILLER_223_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29101_ _29191_/S VGND VGND VPWR VPWR _29120_/S sky130_fd_sc_hd__buf_4
XFILLER_51_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23525_ _23525_/A VGND VGND VPWR VPWR _32257_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20737_ _20733_/X _20736_/X _20704_/X VGND VGND VPWR VPWR _20738_/D sky130_fd_sc_hd__o21ba_1
XFILLER_141_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27293_ _27293_/A VGND VGND VPWR VPWR _34033_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29032_ _34825_/Q _27193_/X _29048_/S VGND VGND VPWR VPWR _29033_/A sky130_fd_sc_hd__mux2_1
X_26244_ _24837_/X _33570_/Q _26258_/S VGND VGND VPWR VPWR _26245_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23456_ _23456_/A VGND VGND VPWR VPWR _32230_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20668_ _22366_/A VGND VGND VPWR VPWR _22536_/A sky130_fd_sc_hd__buf_12
XFILLER_109_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22407_ _32647_/Q _32583_/Q _32519_/Q _35975_/Q _22229_/X _22366_/X VGND VGND VPWR
+ VPWR _22407_/X sky130_fd_sc_hd__mux4_1
X_26175_ _26175_/A VGND VGND VPWR VPWR _33537_/D sky130_fd_sc_hd__clkbuf_1
X_23387_ input24/X VGND VGND VPWR VPWR _23387_/X sky130_fd_sc_hd__clkbuf_4
X_20599_ _20599_/A VGND VGND VPWR VPWR _22373_/A sky130_fd_sc_hd__buf_2
XFILLER_104_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25126_ _24988_/X _33043_/Q _25130_/S VGND VGND VPWR VPWR _25127_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22338_ _32133_/Q _32325_/Q _32389_/Q _35909_/Q _22233_/X _22021_/X VGND VGND VPWR
+ VPWR _22338_/X sky130_fd_sc_hd__mux4_1
XFILLER_191_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29934_ _35222_/Q _29328_/X _29952_/S VGND VGND VPWR VPWR _29935_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25057_ _24886_/X _33010_/Q _25059_/S VGND VGND VPWR VPWR _25058_/A sky130_fd_sc_hd__mux2_1
X_22269_ _22265_/X _22268_/X _22093_/X _22094_/X VGND VGND VPWR VPWR _22286_/B sky130_fd_sc_hd__o211a_1
XFILLER_3_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24008_ _24008_/A VGND VGND VPWR VPWR _32546_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29865_ _29865_/A VGND VGND VPWR VPWR _35189_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_1467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16830_ _35691_/Q _32199_/Q _35563_/Q _35499_/Q _16611_/X _16612_/X VGND VGND VPWR
+ VPWR _16830_/X sky130_fd_sc_hd__mux4_1
X_28816_ _28816_/A VGND VGND VPWR VPWR _34722_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29796_ _29796_/A VGND VGND VPWR VPWR _35157_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28747_ _34691_/Q _27174_/X _28755_/S VGND VGND VPWR VPWR _28748_/A sky130_fd_sc_hd__mux2_1
X_16761_ _16757_/X _16760_/X _16445_/X VGND VGND VPWR VPWR _16769_/C sky130_fd_sc_hd__o21ba_1
X_25959_ _24815_/X _33435_/Q _25967_/S VGND VGND VPWR VPWR _25960_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18500_ _18494_/X _18499_/X _18375_/X VGND VGND VPWR VPWR _18508_/C sky130_fd_sc_hd__o21ba_1
XFILLER_189_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16692_ _16447_/X _16690_/X _16691_/X _16450_/X VGND VGND VPWR VPWR _16692_/X sky130_fd_sc_hd__a22o_1
X_19480_ _32885_/Q _32821_/Q _32757_/Q _32693_/Q _19293_/X _19294_/X VGND VGND VPWR
+ VPWR _19480_/X sky130_fd_sc_hd__mux4_1
XFILLER_234_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_1382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28678_ _34658_/Q _27072_/X _28692_/S VGND VGND VPWR VPWR _28679_/A sky130_fd_sc_hd__mux2_1
XFILLER_206_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18431_ _34647_/Q _34583_/Q _34519_/Q _34455_/Q _18379_/X _18380_/X VGND VGND VPWR
+ VPWR _18431_/X sky130_fd_sc_hd__mux4_1
X_27629_ _34193_/Q _27217_/X _27629_/S VGND VGND VPWR VPWR _27630_/A sky130_fd_sc_hd__mux2_1
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18362_ _20150_/A VGND VGND VPWR VPWR _18362_/X sky130_fd_sc_hd__buf_6
X_30640_ _35557_/Q _29376_/X _30648_/S VGND VGND VPWR VPWR _30641_/A sky130_fd_sc_hd__mux2_1
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17313_ _32121_/Q _32313_/Q _32377_/Q _35897_/Q _17280_/X _17068_/X VGND VGND VPWR
+ VPWR _17313_/X sky130_fd_sc_hd__mux4_1
X_30571_ _30571_/A VGND VGND VPWR VPWR _35524_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18293_ _20099_/A VGND VGND VPWR VPWR _18293_/X sky130_fd_sc_hd__buf_4
XFILLER_30_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32310_ _32885_/CLK _32310_/D VGND VGND VPWR VPWR _32310_/Q sky130_fd_sc_hd__dfxtp_1
X_17244_ _32631_/Q _32567_/Q _32503_/Q _35959_/Q _16923_/X _17060_/X VGND VGND VPWR
+ VPWR _17244_/X sky130_fd_sc_hd__mux4_1
X_33290_ _33420_/CLK _33290_/D VGND VGND VPWR VPWR _33290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32241_ _35730_/CLK _32241_/D VGND VGND VPWR VPWR _32241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17175_ _17171_/X _17174_/X _17132_/X VGND VGND VPWR VPWR _17197_/A sky130_fd_sc_hd__o21ba_1
XFILLER_127_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16126_ _16048_/X _16124_/X _16125_/X _16058_/X VGND VGND VPWR VPWR _16126_/X sky130_fd_sc_hd__a22o_1
XFILLER_155_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32172_ _35180_/CLK _32172_/D VGND VGND VPWR VPWR _32172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31123_ _35786_/Q input48/X _31137_/S VGND VGND VPWR VPWR _31124_/A sky130_fd_sc_hd__mux2_1
X_16057_ _17771_/A VGND VGND VPWR VPWR _17862_/A sky130_fd_sc_hd__buf_12
XFILLER_142_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35931_ _35994_/CLK _35931_/D VGND VGND VPWR VPWR _35931_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31054_ _31054_/A VGND VGND VPWR VPWR _35753_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30005_ _35256_/Q _29435_/X _30015_/S VGND VGND VPWR VPWR _30006_/A sky130_fd_sc_hd__mux2_1
X_19816_ _20169_/A VGND VGND VPWR VPWR _19816_/X sky130_fd_sc_hd__clkbuf_4
X_35862_ _35863_/CLK _35862_/D VGND VGND VPWR VPWR _35862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34813_ _35448_/CLK _34813_/D VGND VGND VPWR VPWR _34813_/Q sky130_fd_sc_hd__dfxtp_1
X_19747_ _20261_/A VGND VGND VPWR VPWR _19747_/X sky130_fd_sc_hd__buf_8
XFILLER_238_872 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35793_ _35855_/CLK _35793_/D VGND VGND VPWR VPWR _35793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16959_ _16706_/X _16957_/X _16958_/X _16712_/X VGND VGND VPWR VPWR _16959_/X sky130_fd_sc_hd__a22o_1
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_894 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34744_ _35833_/CLK _34744_/D VGND VGND VPWR VPWR _34744_/Q sky130_fd_sc_hd__dfxtp_1
X_31956_ _23498_/X _36181_/Q _31956_/S VGND VGND VPWR VPWR _31957_/A sky130_fd_sc_hd__mux2_1
X_19678_ _20151_/A VGND VGND VPWR VPWR _19678_/X sky130_fd_sc_hd__buf_6
XFILLER_64_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_936 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18629_ _18625_/X _18628_/X _18344_/X _18346_/X VGND VGND VPWR VPWR _18644_/B sky130_fd_sc_hd__o211a_1
X_30907_ _30907_/A VGND VGND VPWR VPWR _35683_/D sky130_fd_sc_hd__clkbuf_1
X_34675_ _35377_/CLK _34675_/D VGND VGND VPWR VPWR _34675_/Q sky130_fd_sc_hd__dfxtp_1
X_31887_ _31956_/S VGND VGND VPWR VPWR _31906_/S sky130_fd_sc_hd__buf_4
XFILLER_24_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33626_ _36212_/CLK _33626_/D VGND VGND VPWR VPWR _33626_/Q sky130_fd_sc_hd__dfxtp_1
X_21640_ _33073_/Q _32049_/Q _35825_/Q _35761_/Q _21325_/X _21326_/X VGND VGND VPWR
+ VPWR _21640_/X sky130_fd_sc_hd__mux4_1
X_30838_ _35651_/Q input40/X _30846_/S VGND VGND VPWR VPWR _30839_/A sky130_fd_sc_hd__mux2_1
XFILLER_244_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33557_ _36119_/CLK _33557_/D VGND VGND VPWR VPWR _33557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21571_ _21250_/X _21569_/X _21570_/X _21253_/X VGND VGND VPWR VPWR _21571_/X sky130_fd_sc_hd__a22o_1
XFILLER_177_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30769_ _35618_/Q input4/X _30783_/S VGND VGND VPWR VPWR _30770_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23310_ _27232_/B _25132_/A _28786_/A VGND VGND VPWR VPWR _23311_/A sky130_fd_sc_hd__or3_1
X_20522_ _33428_/Q _33364_/Q _33300_/Q _33236_/Q _18337_/X _18339_/X VGND VGND VPWR
+ VPWR _20522_/X sky130_fd_sc_hd__mux4_1
XFILLER_177_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32508_ _35965_/CLK _32508_/D VGND VGND VPWR VPWR _32508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24290_ _24290_/A VGND VGND VPWR VPWR _32677_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33488_ _34064_/CLK _33488_/D VGND VGND VPWR VPWR _33488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23241_ _32153_/Q _23240_/X _23259_/S VGND VGND VPWR VPWR _23242_/A sky130_fd_sc_hd__mux2_1
XFILLER_203_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35227_ _35802_/CLK _35227_/D VGND VGND VPWR VPWR _35227_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20453_ _34449_/Q _36177_/Q _34321_/Q _34257_/Q _20235_/X _20236_/X VGND VGND VPWR
+ VPWR _20453_/X sky130_fd_sc_hd__mux4_1
XFILLER_119_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32439_ _33895_/CLK _32439_/D VGND VGND VPWR VPWR _32439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1084 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35158_ _36118_/CLK _35158_/D VGND VGND VPWR VPWR _35158_/Q sky130_fd_sc_hd__dfxtp_1
X_23172_ _23172_/A VGND VGND VPWR VPWR _32124_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20384_ _35663_/Q _35023_/Q _34383_/Q _33743_/Q _20150_/X _20151_/X VGND VGND VPWR
+ VPWR _20384_/X sky130_fd_sc_hd__mux4_1
XFILLER_133_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22123_ _34175_/Q _34111_/Q _34047_/Q _33983_/Q _22046_/X _22047_/X VGND VGND VPWR
+ VPWR _22123_/X sky130_fd_sc_hd__mux4_1
X_34109_ _34877_/CLK _34109_/D VGND VGND VPWR VPWR _34109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35089_ _36115_/CLK _35089_/D VGND VGND VPWR VPWR _35089_/Q sky130_fd_sc_hd__dfxtp_1
X_27980_ _27980_/A VGND VGND VPWR VPWR _34327_/D sky130_fd_sc_hd__clkbuf_1
Xoutput140 _32013_/Q VGND VGND VPWR VPWR D1[55] sky130_fd_sc_hd__buf_2
XTAP_6506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput151 _31965_/Q VGND VGND VPWR VPWR D1[7] sky130_fd_sc_hd__buf_2
XTAP_6517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput162 _36199_/Q VGND VGND VPWR VPWR D2[17] sky130_fd_sc_hd__buf_2
XFILLER_0_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput173 _36209_/Q VGND VGND VPWR VPWR D2[27] sky130_fd_sc_hd__buf_2
XFILLER_161_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26931_ _33893_/Q _23277_/X _26939_/S VGND VGND VPWR VPWR _26932_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22054_ _32637_/Q _32573_/Q _32509_/Q _35965_/Q _21876_/X _22013_/X VGND VGND VPWR
+ VPWR _22054_/X sky130_fd_sc_hd__mux4_1
XTAP_6539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput184 _36219_/Q VGND VGND VPWR VPWR D2[37] sky130_fd_sc_hd__buf_2
XFILLER_0_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput195 _36229_/Q VGND VGND VPWR VPWR D2[47] sky130_fd_sc_hd__buf_2
XTAP_5805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_844 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21005_ _35423_/Q _35359_/Q _35295_/Q _35231_/Q _20795_/X _20796_/X VGND VGND VPWR
+ VPWR _21005_/X sky130_fd_sc_hd__mux4_1
XFILLER_88_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29650_ _35088_/Q _29509_/X _29652_/S VGND VGND VPWR VPWR _29651_/A sky130_fd_sc_hd__mux2_1
XTAP_5838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26862_ _26862_/A VGND VGND VPWR VPWR _33860_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28601_ _27766_/X _34622_/Q _28619_/S VGND VGND VPWR VPWR _28602_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25813_ _25945_/S VGND VGND VPWR VPWR _25832_/S sky130_fd_sc_hd__buf_6
X_26793_ _26793_/A VGND VGND VPWR VPWR _33827_/D sky130_fd_sc_hd__clkbuf_1
X_29581_ _35055_/Q _29407_/X _29589_/S VGND VGND VPWR VPWR _29582_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28532_ _28532_/A VGND VGND VPWR VPWR _34589_/D sky130_fd_sc_hd__clkbuf_1
X_25744_ _24896_/X _33333_/Q _25760_/S VGND VGND VPWR VPWR _25745_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22956_ input15/X VGND VGND VPWR VPWR _22956_/X sky130_fd_sc_hd__buf_2
XFILLER_112_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21907_ _33913_/Q _33849_/Q _33785_/Q _36089_/Q _21624_/X _21625_/X VGND VGND VPWR
+ VPWR _21907_/X sky130_fd_sc_hd__mux4_1
XFILLER_28_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25675_ _24994_/X _33301_/Q _25675_/S VGND VGND VPWR VPWR _25676_/A sky130_fd_sc_hd__mux2_1
XFILLER_216_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28463_ _27763_/X _34557_/Q _28463_/S VGND VGND VPWR VPWR _28464_/A sky130_fd_sc_hd__mux2_1
X_22887_ _22887_/A VGND VGND VPWR VPWR _23083_/S sky130_fd_sc_hd__buf_8
XFILLER_71_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24626_ _23033_/X _32837_/Q _24630_/S VGND VGND VPWR VPWR _24627_/A sky130_fd_sc_hd__mux2_1
X_27414_ _27414_/A VGND VGND VPWR VPWR _34090_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28394_ _27661_/X _34524_/Q _28400_/S VGND VGND VPWR VPWR _28395_/A sky130_fd_sc_hd__mux2_1
X_21838_ _34167_/Q _34103_/Q _34039_/Q _33975_/Q _21693_/X _21694_/X VGND VGND VPWR
+ VPWR _21838_/X sky130_fd_sc_hd__mux4_1
XFILLER_231_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27345_ _34058_/Q _27196_/X _27359_/S VGND VGND VPWR VPWR _27346_/A sky130_fd_sc_hd__mux2_1
X_24557_ _22931_/X _32804_/Q _24567_/S VGND VGND VPWR VPWR _24558_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21769_ _33653_/Q _33589_/Q _33525_/Q _33461_/Q _21447_/X _21448_/X VGND VGND VPWR
+ VPWR _21769_/X sky130_fd_sc_hd__mux4_1
XFILLER_106_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23508_ _23508_/A VGND VGND VPWR VPWR _32249_/D sky130_fd_sc_hd__clkbuf_1
X_27276_ _27276_/A VGND VGND VPWR VPWR _34025_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24488_ _24488_/A VGND VGND VPWR VPWR _32771_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29015_ _34817_/Q _27168_/X _29027_/S VGND VGND VPWR VPWR _29016_/A sky130_fd_sc_hd__mux2_1
X_26227_ _24812_/X _33562_/Q _26237_/S VGND VGND VPWR VPWR _26228_/A sky130_fd_sc_hd__mux2_1
X_23439_ _32225_/Q _23438_/X _23451_/S VGND VGND VPWR VPWR _23440_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26158_ _26158_/A VGND VGND VPWR VPWR _33529_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25109_ _25109_/A VGND VGND VPWR VPWR _33034_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26089_ _26089_/A VGND VGND VPWR VPWR _33496_/D sky130_fd_sc_hd__clkbuf_1
X_18980_ _32871_/Q _32807_/Q _32743_/Q _32679_/Q _18940_/X _18941_/X VGND VGND VPWR
+ VPWR _18980_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1078 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29917_ _29917_/A VGND VGND VPWR VPWR _35214_/D sky130_fd_sc_hd__clkbuf_1
X_17931_ _17927_/X _17930_/X _17857_/X VGND VGND VPWR VPWR _17941_/C sky130_fd_sc_hd__o21ba_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17862_ _17862_/A VGND VGND VPWR VPWR _17862_/X sky130_fd_sc_hd__clkbuf_4
X_29848_ _29848_/A VGND VGND VPWR VPWR _35181_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19601_ _19601_/A _19601_/B _19601_/C _19601_/D VGND VGND VPWR VPWR _19602_/A sky130_fd_sc_hd__or4_1
XFILLER_113_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16813_ _16804_/X _16811_/X _16812_/X VGND VGND VPWR VPWR _16814_/D sky130_fd_sc_hd__o21ba_1
X_17793_ _34950_/Q _34886_/Q _34822_/Q _34758_/Q _17513_/X _17514_/X VGND VGND VPWR
+ VPWR _17793_/X sky130_fd_sc_hd__mux4_1
X_29779_ _35149_/Q _29500_/X _29787_/S VGND VGND VPWR VPWR _29780_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31810_ _31810_/A VGND VGND VPWR VPWR _36111_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19532_ _34934_/Q _34870_/Q _34806_/Q _34742_/Q _19460_/X _19461_/X VGND VGND VPWR
+ VPWR _19532_/X sky130_fd_sc_hd__mux4_1
X_16744_ _33385_/Q _33321_/Q _33257_/Q _33193_/Q _16421_/X _16422_/X VGND VGND VPWR
+ VPWR _16744_/X sky130_fd_sc_hd__mux4_1
X_32790_ _32856_/CLK _32790_/D VGND VGND VPWR VPWR _32790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31741_ _31741_/A VGND VGND VPWR VPWR _36078_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19463_ _19463_/A VGND VGND VPWR VPWR _19463_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_235_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16675_ _16669_/X _16674_/X _16426_/X VGND VGND VPWR VPWR _16697_/A sky130_fd_sc_hd__o21ba_1
XFILLER_74_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18414_ _33879_/Q _33815_/Q _33751_/Q _36055_/Q _18412_/X _18413_/X VGND VGND VPWR
+ VPWR _18414_/X sky130_fd_sc_hd__mux4_1
XFILLER_62_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34460_ _36229_/CLK _34460_/D VGND VGND VPWR VPWR _34460_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31672_ _27816_/X _36046_/Q _31678_/S VGND VGND VPWR VPWR _31673_/A sky130_fd_sc_hd__mux2_1
X_19394_ _20261_/A VGND VGND VPWR VPWR _19394_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33411_ _33415_/CLK _33411_/D VGND VGND VPWR VPWR _33411_/Q sky130_fd_sc_hd__dfxtp_1
X_18345_ input82/X VGND VGND VPWR VPWR _20147_/A sky130_fd_sc_hd__buf_6
X_30623_ _35549_/Q _29351_/X _30627_/S VGND VGND VPWR VPWR _30624_/A sky130_fd_sc_hd__mux2_1
X_34391_ _34647_/CLK _34391_/D VGND VGND VPWR VPWR _34391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_1219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36130_ _36210_/CLK _36130_/D VGND VGND VPWR VPWR _36130_/Q sky130_fd_sc_hd__dfxtp_1
X_33342_ _35648_/CLK _33342_/D VGND VGND VPWR VPWR _33342_/Q sky130_fd_sc_hd__dfxtp_1
X_18276_ _18272_/X _18275_/X _17871_/A VGND VGND VPWR VPWR _18277_/D sky130_fd_sc_hd__o21ba_1
X_30554_ _30554_/A VGND VGND VPWR VPWR _35516_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36061_ _36128_/CLK _36061_/D VGND VGND VPWR VPWR _36061_/Q sky130_fd_sc_hd__dfxtp_1
Xinput20 DW[27] VGND VGND VPWR VPWR input20/X sky130_fd_sc_hd__buf_4
X_17227_ _35190_/Q _35126_/Q _35062_/Q _32246_/Q _17010_/X _17011_/X VGND VGND VPWR
+ VPWR _17227_/X sky130_fd_sc_hd__mux4_1
Xinput31 DW[37] VGND VGND VPWR VPWR input31/X sky130_fd_sc_hd__buf_4
X_33273_ _36090_/CLK _33273_/D VGND VGND VPWR VPWR _33273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30485_ _30485_/A VGND VGND VPWR VPWR _35483_/D sky130_fd_sc_hd__clkbuf_1
Xinput42 DW[47] VGND VGND VPWR VPWR input42/X sky130_fd_sc_hd__buf_8
XFILLER_174_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35012_ _35843_/CLK _35012_/D VGND VGND VPWR VPWR _35012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput53 DW[57] VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__buf_12
X_32224_ _35646_/CLK _32224_/D VGND VGND VPWR VPWR _32224_/Q sky130_fd_sc_hd__dfxtp_1
Xinput64 DW[9] VGND VGND VPWR VPWR input64/X sky130_fd_sc_hd__buf_8
Xinput75 R2[4] VGND VGND VPWR VPWR input75/X sky130_fd_sc_hd__buf_2
XFILLER_122_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17158_ _17158_/A VGND VGND VPWR VPWR _17158_/X sky130_fd_sc_hd__clkbuf_4
Xinput86 RW[3] VGND VGND VPWR VPWR input86/X sky130_fd_sc_hd__buf_4
XFILLER_171_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16109_ _34135_/Q _34071_/Q _34007_/Q _33943_/Q _16009_/X _16011_/X VGND VGND VPWR
+ VPWR _16109_/X sky130_fd_sc_hd__mux4_1
X_32155_ _35800_/CLK _32155_/D VGND VGND VPWR VPWR _32155_/Q sky130_fd_sc_hd__dfxtp_1
X_17089_ _17085_/X _17088_/X _16812_/X VGND VGND VPWR VPWR _17090_/D sky130_fd_sc_hd__o21ba_1
XFILLER_171_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31106_ _35778_/Q input39/X _31116_/S VGND VGND VPWR VPWR _31107_/A sky130_fd_sc_hd__mux2_1
XFILLER_135_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32086_ _34708_/CLK _32086_/D VGND VGND VPWR VPWR _32086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_233_1022 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35914_ _35978_/CLK _35914_/D VGND VGND VPWR VPWR _35914_/Q sky130_fd_sc_hd__dfxtp_1
X_31037_ _35745_/Q input3/X _31053_/S VGND VGND VPWR VPWR _31038_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35845_ _35845_/CLK _35845_/D VGND VGND VPWR VPWR _35845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_217_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22810_ _34707_/Q _34643_/Q _34579_/Q _34515_/Q _22598_/X _22599_/X VGND VGND VPWR
+ VPWR _22810_/X sky130_fd_sc_hd__mux4_1
XFILLER_72_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35776_ _35839_/CLK _35776_/D VGND VGND VPWR VPWR _35776_/Q sky130_fd_sc_hd__dfxtp_1
X_23790_ _23008_/X _32381_/Q _23790_/S VGND VGND VPWR VPWR _23791_/A sky130_fd_sc_hd__mux2_1
X_32988_ _36054_/CLK _32988_/D VGND VGND VPWR VPWR _32988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22741_ _21758_/A _22739_/X _22740_/X _21763_/A VGND VGND VPWR VPWR _22741_/X sky130_fd_sc_hd__a22o_1
X_34727_ _34921_/CLK _34727_/D VGND VGND VPWR VPWR _34727_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_246_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31939_ _31939_/A VGND VGND VPWR VPWR _36172_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25460_ _25460_/A VGND VGND VPWR VPWR _33198_/D sky130_fd_sc_hd__clkbuf_1
X_22672_ _33423_/Q _33359_/Q _33295_/Q _33231_/Q _22433_/X _22434_/X VGND VGND VPWR
+ VPWR _22672_/X sky130_fd_sc_hd__mux4_2
X_34658_ _36209_/CLK _34658_/D VGND VGND VPWR VPWR _34658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24411_ _22915_/X _32735_/Q _24411_/S VGND VGND VPWR VPWR _24412_/A sky130_fd_sc_hd__mux2_1
X_33609_ _34185_/CLK _33609_/D VGND VGND VPWR VPWR _33609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21623_ _33393_/Q _33329_/Q _33265_/Q _33201_/Q _21374_/X _21375_/X VGND VGND VPWR
+ VPWR _21623_/X sky130_fd_sc_hd__mux4_1
XFILLER_240_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25391_ _33167_/Q _23478_/X _25395_/S VGND VGND VPWR VPWR _25392_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34589_ _36229_/CLK _34589_/D VGND VGND VPWR VPWR _34589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27130_ _27130_/A VGND VGND VPWR VPWR _33972_/D sky130_fd_sc_hd__clkbuf_1
X_24342_ _23011_/X _32702_/Q _24360_/S VGND VGND VPWR VPWR _24343_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21554_ _33903_/Q _33839_/Q _33775_/Q _36079_/Q _21271_/X _21272_/X VGND VGND VPWR
+ VPWR _21554_/X sky130_fd_sc_hd__mux4_1
XFILLER_103_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20505_ _18281_/X _20503_/X _20504_/X _18291_/X VGND VGND VPWR VPWR _20505_/X sky130_fd_sc_hd__a22o_1
X_27061_ _27061_/A VGND VGND VPWR VPWR _33950_/D sky130_fd_sc_hd__clkbuf_1
X_24273_ _24273_/A VGND VGND VPWR VPWR _32669_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21485_ _34157_/Q _34093_/Q _34029_/Q _33965_/Q _21340_/X _21341_/X VGND VGND VPWR
+ VPWR _21485_/X sky130_fd_sc_hd__mux4_1
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26012_ _24892_/X _33460_/Q _26030_/S VGND VGND VPWR VPWR _26013_/A sky130_fd_sc_hd__mux2_1
X_23224_ _23224_/A VGND VGND VPWR VPWR _32149_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20436_ _32657_/Q _32593_/Q _32529_/Q _35985_/Q _20282_/X _19177_/A VGND VGND VPWR
+ VPWR _20436_/X sky130_fd_sc_hd__mux4_1
XFILLER_175_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23155_ _22980_/X _32116_/Q _23173_/S VGND VGND VPWR VPWR _23156_/A sky130_fd_sc_hd__mux2_1
XTAP_7026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20367_ _20367_/A _20367_/B _20367_/C _20367_/D VGND VGND VPWR VPWR _20368_/A sky130_fd_sc_hd__or4_1
XFILLER_175_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22106_ _22459_/A VGND VGND VPWR VPWR _22106_/X sky130_fd_sc_hd__clkbuf_4
XTAP_7059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27963_ _27822_/X _34320_/Q _27965_/S VGND VGND VPWR VPWR _27964_/A sky130_fd_sc_hd__mux2_1
XTAP_6325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23086_ _23086_/A VGND VGND VPWR VPWR _31418_/A sky130_fd_sc_hd__buf_12
XTAP_6336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20298_ _20298_/A VGND VGND VPWR VPWR _20298_/X sky130_fd_sc_hd__buf_6
XFILLER_164_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29702_ _29702_/A VGND VGND VPWR VPWR _35112_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26914_ _33885_/Q _23252_/X _26918_/S VGND VGND VPWR VPWR _26915_/A sky130_fd_sc_hd__mux2_1
X_22037_ _35196_/Q _35132_/Q _35068_/Q _32252_/Q _21963_/X _21964_/X VGND VGND VPWR
+ VPWR _22037_/X sky130_fd_sc_hd__mux4_1
XTAP_6369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27894_ _27720_/X _34287_/Q _27902_/S VGND VGND VPWR VPWR _27895_/A sky130_fd_sc_hd__mux2_1
XTAP_5646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29633_ _29660_/S VGND VGND VPWR VPWR _29652_/S sky130_fd_sc_hd__buf_4
XTAP_4923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26845_ _26845_/A VGND VGND VPWR VPWR _33852_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29564_ _35047_/Q _29382_/X _29568_/S VGND VGND VPWR VPWR _29565_/A sky130_fd_sc_hd__mux2_1
X_23988_ _22897_/X _32537_/Q _24000_/S VGND VGND VPWR VPWR _23989_/A sky130_fd_sc_hd__mux2_1
X_26776_ _26776_/A VGND VGND VPWR VPWR _33819_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_228_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28515_ _31553_/A _31823_/B VGND VGND VPWR VPWR _28648_/S sky130_fd_sc_hd__nand2_8
X_25727_ _24871_/X _33325_/Q _25739_/S VGND VGND VPWR VPWR _25728_/A sky130_fd_sc_hd__mux2_1
X_22939_ _22939_/A VGND VGND VPWR VPWR _32038_/D sky130_fd_sc_hd__clkbuf_1
X_29495_ _35019_/Q _29494_/X _29513_/S VGND VGND VPWR VPWR _29496_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_244_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28446_ _28446_/A VGND VGND VPWR VPWR _34548_/D sky130_fd_sc_hd__clkbuf_1
X_16460_ _16451_/X _16458_/X _16459_/X VGND VGND VPWR VPWR _16461_/D sky130_fd_sc_hd__o21ba_1
XFILLER_243_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25658_ _25658_/A VGND VGND VPWR VPWR _33292_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16391_ _33375_/Q _33311_/Q _33247_/Q _33183_/Q _16002_/X _16003_/X VGND VGND VPWR
+ VPWR _16391_/X sky130_fd_sc_hd__mux4_1
X_24609_ _23008_/X _32829_/Q _24609_/S VGND VGND VPWR VPWR _24610_/A sky130_fd_sc_hd__mux2_1
XPHY_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28377_ _28377_/A VGND VGND VPWR VPWR _34516_/D sky130_fd_sc_hd__clkbuf_1
X_25589_ _25589_/A VGND VGND VPWR VPWR _33259_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18130_ _34193_/Q _34129_/Q _34065_/Q _34001_/Q _16049_/X _16050_/X VGND VGND VPWR
+ VPWR _18130_/X sky130_fd_sc_hd__mux4_1
XPHY_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27328_ _34050_/Q _27171_/X _27338_/S VGND VGND VPWR VPWR _27329_/A sky130_fd_sc_hd__mux2_1
XFILLER_197_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18061_ _35214_/Q _35150_/Q _35086_/Q _32270_/Q _16092_/X _16094_/X VGND VGND VPWR
+ VPWR _18061_/X sky130_fd_sc_hd__mux4_1
X_27259_ _34017_/Q _27069_/X _27275_/S VGND VGND VPWR VPWR _27260_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17012_ _35184_/Q _35120_/Q _35056_/Q _32187_/Q _17010_/X _17011_/X VGND VGND VPWR
+ VPWR _17012_/X sky130_fd_sc_hd__mux4_1
X_30270_ _30270_/A VGND VGND VPWR VPWR _35381_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_180_CLK clkbuf_6_27__f_CLK/X VGND VGND VPWR VPWR _35729_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_193_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18963_ _18752_/X _18961_/X _18962_/X _18757_/X VGND VGND VPWR VPWR _18963_/X sky130_fd_sc_hd__a22o_1
XFILLER_152_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17914_ _33930_/Q _33866_/Q _33802_/Q _36106_/Q _17730_/X _17731_/X VGND VGND VPWR
+ VPWR _17914_/X sky130_fd_sc_hd__mux4_1
X_33960_ _34920_/CLK _33960_/D VGND VGND VPWR VPWR _33960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18894_ _18890_/X _18893_/X _18759_/X VGND VGND VPWR VPWR _18895_/D sky130_fd_sc_hd__o21ba_1
XTAP_6870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32911_ _32911_/CLK _32911_/D VGND VGND VPWR VPWR _32911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17845_ _17773_/X _17843_/X _17844_/X _17777_/X VGND VGND VPWR VPWR _17845_/X sky130_fd_sc_hd__a22o_1
X_33891_ _36070_/CLK _33891_/D VGND VGND VPWR VPWR _33891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35630_ _35630_/CLK _35630_/D VGND VGND VPWR VPWR _35630_/Q sky130_fd_sc_hd__dfxtp_1
X_32842_ _32906_/CLK _32842_/D VGND VGND VPWR VPWR _32842_/Q sky130_fd_sc_hd__dfxtp_1
X_17776_ _32902_/Q _32838_/Q _32774_/Q _32710_/Q _17699_/X _17700_/X VGND VGND VPWR
+ VPWR _17776_/X sky130_fd_sc_hd__mux4_1
XFILLER_94_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19515_ _32118_/Q _32310_/Q _32374_/Q _35894_/Q _19227_/X _19368_/X VGND VGND VPWR
+ VPWR _19515_/X sky130_fd_sc_hd__mux4_1
X_35561_ _35685_/CLK _35561_/D VGND VGND VPWR VPWR _35561_/Q sky130_fd_sc_hd__dfxtp_1
X_16727_ _33064_/Q _32040_/Q _35816_/Q _35752_/Q _16725_/X _16726_/X VGND VGND VPWR
+ VPWR _16727_/X sky130_fd_sc_hd__mux4_1
X_32773_ _32903_/CLK _32773_/D VGND VGND VPWR VPWR _32773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34512_ _34705_/CLK _34512_/D VGND VGND VPWR VPWR _34512_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31724_ _31724_/A VGND VGND VPWR VPWR _36070_/D sky130_fd_sc_hd__clkbuf_1
X_19446_ _35636_/Q _34996_/Q _34356_/Q _33716_/Q _19444_/X _19445_/X VGND VGND VPWR
+ VPWR _19446_/X sky130_fd_sc_hd__mux4_1
XFILLER_35_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16658_ _17011_/A VGND VGND VPWR VPWR _16658_/X sky130_fd_sc_hd__buf_4
X_35492_ _35684_/CLK _35492_/D VGND VGND VPWR VPWR _35492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34443_ _36171_/CLK _34443_/D VGND VGND VPWR VPWR _34443_/Q sky130_fd_sc_hd__dfxtp_1
X_31655_ _27791_/X _36038_/Q _31657_/S VGND VGND VPWR VPWR _31656_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19377_ _35442_/Q _35378_/Q _35314_/Q _35250_/Q _19201_/X _19202_/X VGND VGND VPWR
+ VPWR _19377_/X sky130_fd_sc_hd__mux4_1
X_16589_ _35172_/Q _35108_/Q _35044_/Q _32164_/Q _16304_/X _16305_/X VGND VGND VPWR
+ VPWR _16589_/X sky130_fd_sc_hd__mux4_1
XFILLER_245_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18328_ _18318_/X _18323_/X _18326_/X _18327_/X VGND VGND VPWR VPWR _18328_/X sky130_fd_sc_hd__a22o_1
X_30606_ _30606_/A VGND VGND VPWR VPWR _35541_/D sky130_fd_sc_hd__clkbuf_1
X_34374_ _35717_/CLK _34374_/D VGND VGND VPWR VPWR _34374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31586_ _27689_/X _36005_/Q _31594_/S VGND VGND VPWR VPWR _31587_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_6_36__f_CLK clkbuf_5_18_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_36__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_36113_ _36113_/CLK _36113_/D VGND VGND VPWR VPWR _36113_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33325_ _36077_/CLK _33325_/D VGND VGND VPWR VPWR _33325_/Q sky130_fd_sc_hd__dfxtp_1
X_18259_ _32149_/Q _32341_/Q _32405_/Q _35925_/Q _17986_/X _17011_/A VGND VGND VPWR
+ VPWR _18259_/X sky130_fd_sc_hd__mux4_1
X_30537_ _35508_/Q _29422_/X _30555_/S VGND VGND VPWR VPWR _30538_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36044_ _36044_/CLK _36044_/D VGND VGND VPWR VPWR _36044_/Q sky130_fd_sc_hd__dfxtp_1
X_33256_ _36068_/CLK _33256_/D VGND VGND VPWR VPWR _33256_/Q sky130_fd_sc_hd__dfxtp_1
X_21270_ _33383_/Q _33319_/Q _33255_/Q _33191_/Q _21021_/X _21022_/X VGND VGND VPWR
+ VPWR _21270_/X sky130_fd_sc_hd__mux4_1
X_30468_ _35476_/Q _29521_/X _30470_/S VGND VGND VPWR VPWR _30469_/A sky130_fd_sc_hd__mux2_1
XFILLER_239_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_1076 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20221_ _32138_/Q _32330_/Q _32394_/Q _35914_/Q _19933_/X _20074_/X VGND VGND VPWR
+ VPWR _20221_/X sky130_fd_sc_hd__mux4_1
X_32207_ _35697_/CLK _32207_/D VGND VGND VPWR VPWR _32207_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_171_CLK clkbuf_6_28__f_CLK/X VGND VGND VPWR VPWR _35733_/CLK sky130_fd_sc_hd__clkbuf_16
X_33187_ _33573_/CLK _33187_/D VGND VGND VPWR VPWR _33187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_235_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30399_ _35443_/Q _29419_/X _30399_/S VGND VGND VPWR VPWR _30400_/A sky130_fd_sc_hd__mux2_1
XFILLER_239_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20152_ _35656_/Q _35016_/Q _34376_/Q _33736_/Q _20150_/X _20151_/X VGND VGND VPWR
+ VPWR _20152_/X sky130_fd_sc_hd__mux4_1
XFILLER_172_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32138_ _32907_/CLK _32138_/D VGND VGND VPWR VPWR _32138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24960_ _24960_/A VGND VGND VPWR VPWR _32969_/D sky130_fd_sc_hd__clkbuf_1
X_20083_ _35462_/Q _35398_/Q _35334_/Q _35270_/Q _19907_/X _19908_/X VGND VGND VPWR
+ VPWR _20083_/X sky130_fd_sc_hd__mux4_1
X_32069_ _35779_/CLK _32069_/D VGND VGND VPWR VPWR _32069_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23911_ _22984_/X _32501_/Q _23927_/S VGND VGND VPWR VPWR _23912_/A sky130_fd_sc_hd__mux2_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24891_ _24891_/A VGND VGND VPWR VPWR _32947_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_131_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26630_ _33750_/Q _23225_/X _26648_/S VGND VGND VPWR VPWR _26631_/A sky130_fd_sc_hd__mux2_1
X_23842_ _27232_/B input83/X input89/X _25132_/A VGND VGND VPWR VPWR _23843_/A sky130_fd_sc_hd__and4bb_1
XTAP_3529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35828_ _35828_/CLK _35828_/D VGND VGND VPWR VPWR _35828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_245_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26561_ _26561_/A VGND VGND VPWR VPWR _33719_/D sky130_fd_sc_hd__clkbuf_1
X_35759_ _36015_/CLK _35759_/D VGND VGND VPWR VPWR _35759_/Q sky130_fd_sc_hd__dfxtp_1
X_23773_ _23773_/A VGND VGND VPWR VPWR _32372_/D sky130_fd_sc_hd__clkbuf_1
X_20985_ _20985_/A VGND VGND VPWR VPWR _36190_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28300_ _28300_/A VGND VGND VPWR VPWR _34479_/D sky130_fd_sc_hd__clkbuf_1
X_22724_ _34960_/Q _34896_/Q _34832_/Q _34768_/Q _22466_/X _22467_/X VGND VGND VPWR
+ VPWR _22724_/X sky130_fd_sc_hd__mux4_1
X_25512_ _25512_/A VGND VGND VPWR VPWR _33223_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29280_ _29280_/A VGND VGND VPWR VPWR _34942_/D sky130_fd_sc_hd__clkbuf_1
X_26492_ _26492_/A VGND VGND VPWR VPWR _33686_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_240_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28231_ _27819_/X _34447_/Q _28235_/S VGND VGND VPWR VPWR _28232_/A sky130_fd_sc_hd__mux2_1
XFILLER_198_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25443_ _25443_/A VGND VGND VPWR VPWR _33190_/D sky130_fd_sc_hd__clkbuf_1
X_22655_ _20581_/X _22653_/X _22654_/X _20591_/X VGND VGND VPWR VPWR _22655_/X sky130_fd_sc_hd__a22o_1
XFILLER_240_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21606_ _22469_/A VGND VGND VPWR VPWR _21606_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_166_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25374_ _33159_/Q _23450_/X _25374_/S VGND VGND VPWR VPWR _25375_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28162_ _27717_/X _34414_/Q _28172_/S VGND VGND VPWR VPWR _28163_/A sky130_fd_sc_hd__mux2_1
X_22586_ _22586_/A VGND VGND VPWR VPWR _22586_/X sky130_fd_sc_hd__buf_6
XFILLER_220_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24325_ _22987_/X _32694_/Q _24339_/S VGND VGND VPWR VPWR _24326_/A sky130_fd_sc_hd__mux2_1
X_27113_ _33967_/Q _27112_/X _27125_/S VGND VGND VPWR VPWR _27114_/A sky130_fd_sc_hd__mux2_1
X_28093_ _28093_/A VGND VGND VPWR VPWR _34381_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_903 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21537_ _21250_/X _21535_/X _21536_/X _21253_/X VGND VGND VPWR VPWR _21537_/X sky130_fd_sc_hd__a22o_1
XFILLER_107_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_1307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27044_ input34/X VGND VGND VPWR VPWR _27044_/X sky130_fd_sc_hd__clkbuf_4
X_24256_ _31553_/B _31283_/B VGND VGND VPWR VPWR _24389_/S sky130_fd_sc_hd__nand2_8
XFILLER_119_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21468_ _21245_/X _21466_/X _21467_/X _21248_/X VGND VGND VPWR VPWR _21468_/X sky130_fd_sc_hd__a22o_1
XFILLER_153_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23207_ _23058_/X _32141_/Q _23215_/S VGND VGND VPWR VPWR _23208_/A sky130_fd_sc_hd__mux2_1
X_20419_ _20415_/X _20418_/X _20157_/X VGND VGND VPWR VPWR _20427_/C sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_162_CLK clkbuf_6_30__f_CLK/X VGND VGND VPWR VPWR _35217_/CLK sky130_fd_sc_hd__clkbuf_16
X_24187_ _32630_/Q _23396_/X _24201_/S VGND VGND VPWR VPWR _24188_/A sky130_fd_sc_hd__mux2_1
XFILLER_175_1042 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21399_ _21394_/X _21397_/X _21398_/X VGND VGND VPWR VPWR _21414_/C sky130_fd_sc_hd__o21ba_1
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23138_ _22956_/X _32108_/Q _23152_/S VGND VGND VPWR VPWR _23139_/A sky130_fd_sc_hd__mux2_1
XTAP_6111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28995_ _28995_/A VGND VGND VPWR VPWR _34807_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27946_ _27973_/S VGND VGND VPWR VPWR _27965_/S sky130_fd_sc_hd__buf_4
XTAP_6155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23069_ _23069_/A VGND VGND VPWR VPWR _32080_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_983 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27877_ _27695_/X _34279_/Q _27881_/S VGND VGND VPWR VPWR _27878_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29616_ _29616_/A VGND VGND VPWR VPWR _35071_/D sky130_fd_sc_hd__clkbuf_1
X_17630_ _32642_/Q _32578_/Q _32514_/Q _35970_/Q _17629_/X _17413_/X VGND VGND VPWR
+ VPWR _17630_/X sky130_fd_sc_hd__mux4_1
XTAP_5498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26828_ _33844_/Q _23387_/X _26846_/S VGND VGND VPWR VPWR _26829_/A sky130_fd_sc_hd__mux2_1
XFILLER_236_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29547_ _35039_/Q _29357_/X _29547_/S VGND VGND VPWR VPWR _29548_/A sky130_fd_sc_hd__mux2_1
X_17561_ _33920_/Q _33856_/Q _33792_/Q _36096_/Q _17377_/X _17378_/X VGND VGND VPWR
+ VPWR _17561_/X sky130_fd_sc_hd__mux4_1
XFILLER_29_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26759_ _33812_/Q _23495_/X _26761_/S VGND VGND VPWR VPWR _26760_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19300_ _35632_/Q _34992_/Q _34352_/Q _33712_/Q _19091_/X _19092_/X VGND VGND VPWR
+ VPWR _19300_/X sky130_fd_sc_hd__mux4_1
XFILLER_182_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16512_ _16508_/X _16511_/X _16434_/X _16435_/X VGND VGND VPWR VPWR _16529_/B sky130_fd_sc_hd__o211a_1
X_29478_ input43/X VGND VGND VPWR VPWR _29478_/X sky130_fd_sc_hd__buf_2
X_17492_ _17420_/X _17490_/X _17491_/X _17424_/X VGND VGND VPWR VPWR _17492_/X sky130_fd_sc_hd__a22o_1
XFILLER_210_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_878 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19231_ _19226_/X _19230_/X _19087_/X _19088_/X VGND VGND VPWR VPWR _19248_/B sky130_fd_sc_hd__o211a_1
XFILLER_147_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28429_ _28429_/A VGND VGND VPWR VPWR _34540_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16443_ _33056_/Q _32032_/Q _35808_/Q _35744_/Q _16372_/X _16373_/X VGND VGND VPWR
+ VPWR _16443_/X sky130_fd_sc_hd__mux4_1
XFILLER_204_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31440_ _31551_/S VGND VGND VPWR VPWR _31459_/S sky130_fd_sc_hd__buf_4
X_19162_ _32108_/Q _32300_/Q _32364_/Q _35884_/Q _18874_/X _19015_/X VGND VGND VPWR
+ VPWR _19162_/X sky130_fd_sc_hd__mux4_1
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16374_ _33054_/Q _32030_/Q _35806_/Q _35742_/Q _16372_/X _16373_/X VGND VGND VPWR
+ VPWR _16374_/X sky130_fd_sc_hd__mux4_1
XFILLER_83_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_932 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18113_ _35728_/Q _32239_/Q _35600_/Q _35536_/Q _15993_/X _15995_/X VGND VGND VPWR
+ VPWR _18113_/X sky130_fd_sc_hd__mux4_1
XFILLER_121_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31371_ _27770_/X _35903_/Q _31387_/S VGND VGND VPWR VPWR _31372_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19093_ _35626_/Q _34986_/Q _34346_/Q _33706_/Q _19091_/X _19092_/X VGND VGND VPWR
+ VPWR _19093_/X sky130_fd_sc_hd__mux4_1
XFILLER_184_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33110_ _35863_/CLK _33110_/D VGND VGND VPWR VPWR _33110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18044_ _17912_/X _18042_/X _18043_/X _17915_/X VGND VGND VPWR VPWR _18044_/X sky130_fd_sc_hd__a22o_1
X_30322_ _30322_/A VGND VGND VPWR VPWR _35406_/D sky130_fd_sc_hd__clkbuf_1
X_34090_ _35690_/CLK _34090_/D VGND VGND VPWR VPWR _34090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33041_ _35857_/CLK _33041_/D VGND VGND VPWR VPWR _33041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_153_CLK clkbuf_6_31__f_CLK/X VGND VGND VPWR VPWR _36179_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_158_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30253_ _30253_/A VGND VGND VPWR VPWR _35373_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_236_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30184_ _35341_/Q _29500_/X _30192_/S VGND VGND VPWR VPWR _30185_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19995_ _32644_/Q _32580_/Q _32516_/Q _35972_/Q _19929_/X _19713_/X VGND VGND VPWR
+ VPWR _19995_/X sky130_fd_sc_hd__mux4_1
XFILLER_63_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18946_ _35686_/Q _32193_/Q _35558_/Q _35494_/Q _18911_/X _18912_/X VGND VGND VPWR
+ VPWR _18946_/X sky130_fd_sc_hd__mux4_1
X_34992_ _35632_/CLK _34992_/D VGND VGND VPWR VPWR _34992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33943_ _34135_/CLK _33943_/D VGND VGND VPWR VPWR _33943_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18877_ _18661_/X _18875_/X _18876_/X _18665_/X VGND VGND VPWR VPWR _18877_/X sky130_fd_sc_hd__a22o_1
XFILLER_104_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17828_ _17828_/A _17828_/B _17828_/C _17828_/D VGND VGND VPWR VPWR _17829_/A sky130_fd_sc_hd__or4_1
XFILLER_227_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33874_ _36179_/CLK _33874_/D VGND VGND VPWR VPWR _33874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35613_ _35613_/CLK _35613_/D VGND VGND VPWR VPWR _35613_/Q sky130_fd_sc_hd__dfxtp_1
X_32825_ _35895_/CLK _32825_/D VGND VGND VPWR VPWR _32825_/Q sky130_fd_sc_hd__dfxtp_1
X_17759_ _34182_/Q _34118_/Q _34054_/Q _33990_/Q _17446_/X _17447_/X VGND VGND VPWR
+ VPWR _17759_/X sky130_fd_sc_hd__mux4_1
XFILLER_214_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35544_ _35544_/CLK _35544_/D VGND VGND VPWR VPWR _35544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20770_ _22316_/A VGND VGND VPWR VPWR _20770_/X sky130_fd_sc_hd__buf_6
X_32756_ _32882_/CLK _32756_/D VGND VGND VPWR VPWR _32756_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31707_ _31707_/A VGND VGND VPWR VPWR _36062_/D sky130_fd_sc_hd__clkbuf_1
X_19429_ _33396_/Q _33332_/Q _33268_/Q _33204_/Q _19427_/X _19428_/X VGND VGND VPWR
+ VPWR _19429_/X sky130_fd_sc_hd__mux4_1
X_35475_ _35666_/CLK _35475_/D VGND VGND VPWR VPWR _35475_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32687_ _32911_/CLK _32687_/D VGND VGND VPWR VPWR _32687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22440_ _32648_/Q _32584_/Q _32520_/Q _35976_/Q _22229_/X _22366_/X VGND VGND VPWR
+ VPWR _22440_/X sky130_fd_sc_hd__mux4_1
X_34426_ _36153_/CLK _34426_/D VGND VGND VPWR VPWR _34426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31638_ _31686_/S VGND VGND VPWR VPWR _31657_/S sky130_fd_sc_hd__buf_4
XFILLER_164_903 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22371_ _22371_/A VGND VGND VPWR VPWR _22371_/X sky130_fd_sc_hd__clkbuf_4
X_34357_ _35830_/CLK _34357_/D VGND VGND VPWR VPWR _34357_/Q sky130_fd_sc_hd__dfxtp_1
X_31569_ _27664_/X _35997_/Q _31573_/S VGND VGND VPWR VPWR _31570_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_392_CLK clkbuf_6_40__f_CLK/X VGND VGND VPWR VPWR _34166_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_175_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24110_ _24110_/A VGND VGND VPWR VPWR _32595_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33308_ _36188_/CLK _33308_/D VGND VGND VPWR VPWR _33308_/Q sky130_fd_sc_hd__dfxtp_1
X_21322_ _35624_/Q _34984_/Q _34344_/Q _33704_/Q _21038_/X _21039_/X VGND VGND VPWR
+ VPWR _21322_/X sky130_fd_sc_hd__mux4_1
X_25090_ _25090_/A VGND VGND VPWR VPWR _33025_/D sky130_fd_sc_hd__clkbuf_1
X_34288_ _36143_/CLK _34288_/D VGND VGND VPWR VPWR _34288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36027_ _36027_/CLK _36027_/D VGND VGND VPWR VPWR _36027_/Q sky130_fd_sc_hd__dfxtp_1
X_24041_ _24041_/A VGND VGND VPWR VPWR _32562_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_144_CLK clkbuf_6_28__f_CLK/X VGND VGND VPWR VPWR _32856_/CLK sky130_fd_sc_hd__clkbuf_16
X_33239_ _36059_/CLK _33239_/D VGND VGND VPWR VPWR _33239_/Q sky130_fd_sc_hd__dfxtp_1
X_21253_ _22469_/A VGND VGND VPWR VPWR _21253_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_176_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20204_ _20204_/A VGND VGND VPWR VPWR _32457_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_176_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21184_ _20897_/X _21182_/X _21183_/X _20900_/X VGND VGND VPWR VPWR _21184_/X sky130_fd_sc_hd__a22o_1
XFILLER_85_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27800_ _27800_/A VGND VGND VPWR VPWR _34248_/D sky130_fd_sc_hd__clkbuf_1
X_20135_ _33416_/Q _33352_/Q _33288_/Q _33224_/Q _20133_/X _20134_/X VGND VGND VPWR
+ VPWR _20135_/X sky130_fd_sc_hd__mux4_1
XFILLER_172_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28780_ _34707_/Q _27223_/X _28784_/S VGND VGND VPWR VPWR _28781_/A sky130_fd_sc_hd__mux2_1
X_25992_ _25992_/A VGND VGND VPWR VPWR _33450_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_217_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27731_ _27731_/A VGND VGND VPWR VPWR _34226_/D sky130_fd_sc_hd__clkbuf_1
X_24943_ _24942_/X _32964_/Q _24952_/S VGND VGND VPWR VPWR _24944_/A sky130_fd_sc_hd__mux2_1
X_20066_ _20066_/A VGND VGND VPWR VPWR _20066_/X sky130_fd_sc_hd__clkbuf_4
XTAP_4016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27662_ _27661_/X _34204_/Q _27671_/S VGND VGND VPWR VPWR _27663_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24874_ input17/X VGND VGND VPWR VPWR _24874_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_73_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29401_ input16/X VGND VGND VPWR VPWR _29401_/X sky130_fd_sc_hd__buf_2
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26613_ _26613_/A VGND VGND VPWR VPWR _33744_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23825_ _23825_/A VGND VGND VPWR VPWR _32397_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27593_ _27593_/A VGND VGND VPWR VPWR _34175_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29332_ _29332_/A VGND VGND VPWR VPWR _34966_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26544_ _26544_/A VGND VGND VPWR VPWR _33711_/D sky130_fd_sc_hd__clkbuf_1
X_23756_ _23756_/A VGND VGND VPWR VPWR _32364_/D sky130_fd_sc_hd__clkbuf_1
X_20968_ _35678_/Q _32184_/Q _35550_/Q _35486_/Q _20858_/X _20859_/X VGND VGND VPWR
+ VPWR _20968_/X sky130_fd_sc_hd__mux4_1
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22707_ _33168_/Q _36048_/Q _33040_/Q _32976_/Q _20632_/X _21761_/A VGND VGND VPWR
+ VPWR _22707_/X sky130_fd_sc_hd__mux4_1
XFILLER_148_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29263_ _29263_/A VGND VGND VPWR VPWR _34934_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26475_ _26475_/A VGND VGND VPWR VPWR _33679_/D sky130_fd_sc_hd__clkbuf_1
X_23687_ _23687_/A VGND VGND VPWR VPWR _32333_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20899_ _33052_/Q _32028_/Q _35804_/Q _35740_/Q _20667_/X _20669_/X VGND VGND VPWR
+ VPWR _20899_/X sky130_fd_sc_hd__mux4_1
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28214_ _27794_/X _34439_/Q _28214_/S VGND VGND VPWR VPWR _28215_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22638_ _22638_/A VGND VGND VPWR VPWR _36237_/D sky130_fd_sc_hd__clkbuf_1
X_25426_ _25426_/A VGND VGND VPWR VPWR _33182_/D sky130_fd_sc_hd__clkbuf_1
X_29194_ _29326_/S VGND VGND VPWR VPWR _29213_/S sky130_fd_sc_hd__buf_4
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25357_ _25357_/A VGND VGND VPWR VPWR _33150_/D sky130_fd_sc_hd__clkbuf_1
X_28145_ _27692_/X _34406_/Q _28151_/S VGND VGND VPWR VPWR _28146_/A sky130_fd_sc_hd__mux2_1
X_22569_ _34443_/Q _36171_/Q _34315_/Q _34251_/Q _22535_/X _22536_/X VGND VGND VPWR
+ VPWR _22569_/X sky130_fd_sc_hd__mux4_1
XFILLER_166_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_383_CLK clkbuf_6_42__f_CLK/X VGND VGND VPWR VPWR _33531_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_103_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16090_ _17773_/A VGND VGND VPWR VPWR _17158_/A sky130_fd_sc_hd__buf_12
X_24308_ _22962_/X _32686_/Q _24318_/S VGND VGND VPWR VPWR _24309_/A sky130_fd_sc_hd__mux2_1
X_28076_ _28076_/A VGND VGND VPWR VPWR _34373_/D sky130_fd_sc_hd__clkbuf_1
X_25288_ _33118_/Q _23255_/X _25290_/S VGND VGND VPWR VPWR _25289_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_997 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27027_ _33939_/Q _23492_/X _27031_/S VGND VGND VPWR VPWR _27028_/A sky130_fd_sc_hd__mux2_1
X_24239_ _32655_/Q _23478_/X _24243_/S VGND VGND VPWR VPWR _24240_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_135_CLK clkbuf_6_23__f_CLK/X VGND VGND VPWR VPWR _36118_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_141_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18800_ _20212_/A VGND VGND VPWR VPWR _18800_/X sky130_fd_sc_hd__buf_4
X_19780_ _20133_/A VGND VGND VPWR VPWR _19780_/X sky130_fd_sc_hd__buf_4
XFILLER_96_728 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28978_ _28978_/A VGND VGND VPWR VPWR _34799_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16992_ _32112_/Q _32304_/Q _32368_/Q _35888_/Q _16927_/X _16715_/X VGND VGND VPWR
+ VPWR _16992_/X sky130_fd_sc_hd__mux4_1
XFILLER_1_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18731_ _32096_/Q _32288_/Q _32352_/Q _35872_/Q _18521_/X _18662_/X VGND VGND VPWR
+ VPWR _18731_/X sky130_fd_sc_hd__mux4_1
XFILLER_77_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27929_ _27929_/A VGND VGND VPWR VPWR _34303_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18662_ _20074_/A VGND VGND VPWR VPWR _18662_/X sky130_fd_sc_hd__clkbuf_4
X_30940_ _30940_/A VGND VGND VPWR VPWR _35699_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17613_ _34689_/Q _34625_/Q _34561_/Q _34497_/Q _17292_/X _17293_/X VGND VGND VPWR
+ VPWR _17613_/X sky130_fd_sc_hd__mux4_1
XFILLER_63_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30871_ _35667_/Q input58/X _30875_/S VGND VGND VPWR VPWR _30872_/A sky130_fd_sc_hd__mux2_1
X_18593_ _35676_/Q _32182_/Q _35548_/Q _35484_/Q _18558_/X _18559_/X VGND VGND VPWR
+ VPWR _18593_/X sky130_fd_sc_hd__mux4_1
XTAP_4594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32610_ _36002_/CLK _32610_/D VGND VGND VPWR VPWR _32610_/Q sky130_fd_sc_hd__dfxtp_1
X_17544_ _35199_/Q _35135_/Q _35071_/Q _32255_/Q _17363_/X _17364_/X VGND VGND VPWR
+ VPWR _17544_/X sky130_fd_sc_hd__mux4_1
XFILLER_51_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33590_ _33911_/CLK _33590_/D VGND VGND VPWR VPWR _33590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32541_ _35998_/CLK _32541_/D VGND VGND VPWR VPWR _32541_/Q sky130_fd_sc_hd__dfxtp_1
X_17475_ _17475_/A _17475_/B _17475_/C _17475_/D VGND VGND VPWR VPWR _17476_/A sky130_fd_sc_hd__or4_4
XFILLER_189_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19214_ _19214_/A _19214_/B _19214_/C _19214_/D VGND VGND VPWR VPWR _19215_/A sky130_fd_sc_hd__or4_2
X_16426_ _17838_/A VGND VGND VPWR VPWR _16426_/X sky130_fd_sc_hd__buf_4
X_35260_ _35581_/CLK _35260_/D VGND VGND VPWR VPWR _35260_/Q sky130_fd_sc_hd__dfxtp_1
X_32472_ _35992_/CLK _32472_/D VGND VGND VPWR VPWR _32472_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_242_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34211_ _36210_/CLK _34211_/D VGND VGND VPWR VPWR _34211_/Q sky130_fd_sc_hd__dfxtp_1
X_31423_ _31423_/A VGND VGND VPWR VPWR _35927_/D sky130_fd_sc_hd__clkbuf_1
X_19145_ _19145_/A VGND VGND VPWR VPWR _32427_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16357_ _17907_/A VGND VGND VPWR VPWR _16357_/X sky130_fd_sc_hd__clkbuf_4
X_35191_ _35191_/CLK _35191_/D VGND VGND VPWR VPWR _35191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_762 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_374_CLK clkbuf_6_43__f_CLK/X VGND VGND VPWR VPWR _34941_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34142_ _36188_/CLK _34142_/D VGND VGND VPWR VPWR _34142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19076_ _33386_/Q _33322_/Q _33258_/Q _33194_/Q _19074_/X _19075_/X VGND VGND VPWR
+ VPWR _19076_/X sky130_fd_sc_hd__mux4_1
X_31354_ _27745_/X _35895_/Q _31366_/S VGND VGND VPWR VPWR _31355_/A sky130_fd_sc_hd__mux2_1
X_16288_ _17834_/A VGND VGND VPWR VPWR _16288_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_121_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_5_31_0_CLK clkbuf_2_3_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_31_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_161_906 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30305_ _30305_/A VGND VGND VPWR VPWR _35398_/D sky130_fd_sc_hd__clkbuf_1
X_18027_ _33101_/Q _32077_/Q _35853_/Q _35789_/Q _17784_/X _17785_/X VGND VGND VPWR
+ VPWR _18027_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_126_CLK clkbuf_6_21__f_CLK/X VGND VGND VPWR VPWR _34911_/CLK sky130_fd_sc_hd__clkbuf_16
X_34073_ _36219_/CLK _34073_/D VGND VGND VPWR VPWR _34073_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_236_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31285_ _27639_/X _35862_/Q _31303_/S VGND VGND VPWR VPWR _31286_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33024_ _35646_/CLK _33024_/D VGND VGND VPWR VPWR _33024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30236_ _30236_/A VGND VGND VPWR VPWR _35365_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30167_ _35333_/Q _29475_/X _30171_/S VGND VGND VPWR VPWR _30168_/A sky130_fd_sc_hd__mux2_1
X_19978_ _19974_/X _19977_/X _19804_/X VGND VGND VPWR VPWR _19986_/C sky130_fd_sc_hd__o21ba_1
XFILLER_141_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18929_ _33638_/Q _33574_/Q _33510_/Q _33446_/Q _18794_/X _18795_/X VGND VGND VPWR
+ VPWR _18929_/X sky130_fd_sc_hd__mux4_1
XFILLER_140_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34975_ _35615_/CLK _34975_/D VGND VGND VPWR VPWR _34975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30098_ _35300_/Q _29373_/X _30108_/S VGND VGND VPWR VPWR _30099_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21940_ _21806_/X _21938_/X _21939_/X _21809_/X VGND VGND VPWR VPWR _21940_/X sky130_fd_sc_hd__a22o_1
X_33926_ _34177_/CLK _33926_/D VGND VGND VPWR VPWR _33926_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33857_ _36097_/CLK _33857_/D VGND VGND VPWR VPWR _33857_/Q sky130_fd_sc_hd__dfxtp_1
X_21871_ _21799_/X _21869_/X _21870_/X _21804_/X VGND VGND VPWR VPWR _21871_/X sky130_fd_sc_hd__a22o_1
XFILLER_43_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23610_ _22946_/X _32297_/Q _23610_/S VGND VGND VPWR VPWR _23611_/A sky130_fd_sc_hd__mux2_1
X_20822_ _32090_/Q _32282_/Q _32346_/Q _35866_/Q _20821_/X _22467_/A VGND VGND VPWR
+ VPWR _20822_/X sky130_fd_sc_hd__mux4_1
X_32808_ _32808_/CLK _32808_/D VGND VGND VPWR VPWR _32808_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24590_ _24659_/S VGND VGND VPWR VPWR _24609_/S sky130_fd_sc_hd__buf_4
XFILLER_78_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33788_ _36092_/CLK _33788_/D VGND VGND VPWR VPWR _33788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23541_ _32265_/Q _23460_/X _23557_/S VGND VGND VPWR VPWR _23542_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_1003 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20753_ _32600_/Q _32536_/Q _32472_/Q _35928_/Q _22466_/A _22317_/A VGND VGND VPWR
+ VPWR _20753_/X sky130_fd_sc_hd__mux4_1
X_35527_ _35721_/CLK _35527_/D VGND VGND VPWR VPWR _35527_/Q sky130_fd_sc_hd__dfxtp_1
X_32739_ _32871_/CLK _32739_/D VGND VGND VPWR VPWR _32739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26260_ _26350_/S VGND VGND VPWR VPWR _26279_/S sky130_fd_sc_hd__buf_4
XFILLER_51_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35458_ _35458_/CLK _35458_/D VGND VGND VPWR VPWR _35458_/Q sky130_fd_sc_hd__dfxtp_1
X_23472_ input51/X VGND VGND VPWR VPWR _23472_/X sky130_fd_sc_hd__buf_6
XFILLER_196_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20684_ _22366_/A VGND VGND VPWR VPWR _21611_/A sky130_fd_sc_hd__buf_12
XFILLER_17_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25211_ _33082_/Q _23408_/X _25217_/S VGND VGND VPWR VPWR _25212_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22423_ _22106_/X _22421_/X _22422_/X _22109_/X VGND VGND VPWR VPWR _22423_/X sky130_fd_sc_hd__a22o_1
X_34409_ _34915_/CLK _34409_/D VGND VGND VPWR VPWR _34409_/Q sky130_fd_sc_hd__dfxtp_1
X_26191_ _24958_/X _33545_/Q _26207_/S VGND VGND VPWR VPWR _26192_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_1375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_365_CLK clkbuf_6_41__f_CLK/X VGND VGND VPWR VPWR _36150_/CLK sky130_fd_sc_hd__clkbuf_16
X_35389_ _35453_/CLK _35389_/D VGND VGND VPWR VPWR _35389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25142_ _33049_/Q _23240_/X _25154_/S VGND VGND VPWR VPWR _25143_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_1239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22354_ _22111_/X _22352_/X _22353_/X _22116_/X VGND VGND VPWR VPWR _22354_/X sky130_fd_sc_hd__a22o_1
XFILLER_178_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21305_ _21301_/X _21304_/X _21026_/X VGND VGND VPWR VPWR _21337_/A sky130_fd_sc_hd__o21ba_1
XFILLER_237_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_117_CLK clkbuf_6_20__f_CLK/X VGND VGND VPWR VPWR _36223_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_152_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29950_ _35230_/Q _29354_/X _29952_/S VGND VGND VPWR VPWR _29951_/A sky130_fd_sc_hd__mux2_1
X_25073_ _25073_/A VGND VGND VPWR VPWR _33017_/D sky130_fd_sc_hd__clkbuf_1
X_22285_ _22281_/X _22284_/X _22118_/X VGND VGND VPWR VPWR _22286_/D sky130_fd_sc_hd__o21ba_1
XFILLER_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28901_ _34763_/Q _27199_/X _28913_/S VGND VGND VPWR VPWR _28902_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24024_ _22949_/X _32554_/Q _24042_/S VGND VGND VPWR VPWR _24025_/A sky130_fd_sc_hd__mux2_1
X_21236_ _32614_/Q _32550_/Q _32486_/Q _35942_/Q _21170_/X _20954_/X VGND VGND VPWR
+ VPWR _21236_/X sky130_fd_sc_hd__mux4_1
XFILLER_151_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29881_ _29881_/A VGND VGND VPWR VPWR _35197_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_219_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28832_ _34730_/Q _27096_/X _28850_/S VGND VGND VPWR VPWR _28833_/A sky130_fd_sc_hd__mux2_1
X_21167_ _33892_/Q _33828_/Q _33764_/Q _36068_/Q _20918_/X _20919_/X VGND VGND VPWR
+ VPWR _21167_/X sky130_fd_sc_hd__mux4_1
XFILLER_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20118_ _33095_/Q _32071_/Q _35847_/Q _35783_/Q _20084_/X _20085_/X VGND VGND VPWR
+ VPWR _20118_/X sky130_fd_sc_hd__mux4_1
X_28763_ _28763_/A VGND VGND VPWR VPWR _34698_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25975_ _25975_/A VGND VGND VPWR VPWR _33442_/D sky130_fd_sc_hd__clkbuf_1
X_21098_ _22462_/A VGND VGND VPWR VPWR _21098_/X sky130_fd_sc_hd__buf_4
XFILLER_28_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27714_ input16/X VGND VGND VPWR VPWR _27714_/X sky130_fd_sc_hd__buf_2
X_20049_ _34693_/Q _34629_/Q _34565_/Q _34501_/Q _19945_/X _19946_/X VGND VGND VPWR
+ VPWR _20049_/X sky130_fd_sc_hd__mux4_1
X_24926_ _24926_/A VGND VGND VPWR VPWR _32958_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28694_ _28784_/S VGND VGND VPWR VPWR _28713_/S sky130_fd_sc_hd__buf_4
XFILLER_65_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27645_ _27645_/A VGND VGND VPWR VPWR _34198_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24857_ _24857_/A VGND VGND VPWR VPWR _32936_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23808_ _23808_/A VGND VGND VPWR VPWR _32389_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27576_ _27576_/A VGND VGND VPWR VPWR _34167_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24788_ _23073_/X _32914_/Q _24794_/S VGND VGND VPWR VPWR _24789_/A sky130_fd_sc_hd__mux2_1
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29315_ _29315_/A VGND VGND VPWR VPWR _34959_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26527_ _26527_/A VGND VGND VPWR VPWR _33703_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23739_ _23739_/A VGND VGND VPWR VPWR _32356_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29246_ _29246_/A VGND VGND VPWR VPWR _34926_/D sky130_fd_sc_hd__clkbuf_1
X_17260_ _34679_/Q _34615_/Q _34551_/Q _34487_/Q _16939_/X _16940_/X VGND VGND VPWR
+ VPWR _17260_/X sky130_fd_sc_hd__mux4_1
XFILLER_92_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26458_ _26458_/A VGND VGND VPWR VPWR _33671_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16211_ _34138_/Q _34074_/Q _34010_/Q _33946_/Q _16009_/X _16011_/X VGND VGND VPWR
+ VPWR _16211_/X sky130_fd_sc_hd__mux4_1
XFILLER_174_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25409_ _24796_/X _33174_/Q _25427_/S VGND VGND VPWR VPWR _25410_/A sky130_fd_sc_hd__mux2_1
X_29177_ _34894_/Q _27208_/X _29183_/S VGND VGND VPWR VPWR _29178_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17191_ _35189_/Q _35125_/Q _35061_/Q _32242_/Q _17010_/X _17011_/X VGND VGND VPWR
+ VPWR _17191_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_356_CLK clkbuf_6_46__f_CLK/X VGND VGND VPWR VPWR _35645_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_128_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26389_ _26389_/A VGND VGND VPWR VPWR _33638_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_880 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28128_ _27667_/X _34398_/Q _28130_/S VGND VGND VPWR VPWR _28129_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16142_ _17907_/A VGND VGND VPWR VPWR _16142_/X sky130_fd_sc_hd__buf_4
XFILLER_10_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16073_ _16060_/X _16065_/X _16070_/X _16072_/X VGND VGND VPWR VPWR _16073_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_108_CLK clkbuf_leaf_81_CLK/A VGND VGND VPWR VPWR _34007_/CLK sky130_fd_sc_hd__clkbuf_16
X_28059_ _28059_/A VGND VGND VPWR VPWR _34365_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19901_ _32897_/Q _32833_/Q _32769_/Q _32705_/Q _19646_/X _19647_/X VGND VGND VPWR
+ VPWR _19901_/X sky130_fd_sc_hd__mux4_1
X_31070_ _35761_/Q input20/X _31074_/S VGND VGND VPWR VPWR _31071_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_1270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30021_ _30021_/A VGND VGND VPWR VPWR _35263_/D sky130_fd_sc_hd__clkbuf_1
X_19832_ _32127_/Q _32319_/Q _32383_/Q _35903_/Q _19580_/X _19721_/X VGND VGND VPWR
+ VPWR _19832_/X sky130_fd_sc_hd__mux4_1
XFILLER_116_1227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19763_ _19651_/X _19761_/X _19762_/X _19654_/X VGND VGND VPWR VPWR _19763_/X sky130_fd_sc_hd__a22o_1
X_16975_ _16800_/X _16973_/X _16974_/X _16803_/X VGND VGND VPWR VPWR _16975_/X sky130_fd_sc_hd__a22o_1
X_18714_ _18391_/X _18712_/X _18713_/X _18401_/X VGND VGND VPWR VPWR _18714_/X sky130_fd_sc_hd__a22o_1
X_34760_ _34954_/CLK _34760_/D VGND VGND VPWR VPWR _34760_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31972_ _34085_/CLK _31972_/D VGND VGND VPWR VPWR _31972_/Q sky130_fd_sc_hd__dfxtp_1
X_19694_ _19656_/X _19692_/X _19693_/X _19659_/X VGND VGND VPWR VPWR _19694_/X sky130_fd_sc_hd__a22o_1
XTAP_5081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 DW[15] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__buf_6
XTAP_5092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33711_ _35694_/CLK _33711_/D VGND VGND VPWR VPWR _33711_/Q sky130_fd_sc_hd__dfxtp_1
X_18645_ _18645_/A VGND VGND VPWR VPWR _32413_/D sky130_fd_sc_hd__buf_2
X_30923_ _35691_/Q input14/X _30939_/S VGND VGND VPWR VPWR _30924_/A sky130_fd_sc_hd__mux2_1
X_34691_ _34691_/CLK _34691_/D VGND VGND VPWR VPWR _34691_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33642_ _35690_/CLK _33642_/D VGND VGND VPWR VPWR _33642_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30854_ _30854_/A VGND VGND VPWR VPWR _35658_/D sky130_fd_sc_hd__clkbuf_1
X_18576_ _33628_/Q _33564_/Q _33500_/Q _33436_/Q _18441_/X _18442_/X VGND VGND VPWR
+ VPWR _18576_/X sky130_fd_sc_hd__mux4_1
XTAP_3690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17527_ _17206_/X _17525_/X _17526_/X _17209_/X VGND VGND VPWR VPWR _17527_/X sky130_fd_sc_hd__a22o_1
XFILLER_127_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33573_ _33573_/CLK _33573_/D VGND VGND VPWR VPWR _33573_/Q sky130_fd_sc_hd__dfxtp_1
X_30785_ _30875_/S VGND VGND VPWR VPWR _30804_/S sky130_fd_sc_hd__buf_4
XFILLER_178_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35312_ _35633_/CLK _35312_/D VGND VGND VPWR VPWR _35312_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32524_ _32655_/CLK _32524_/D VGND VGND VPWR VPWR _32524_/Q sky130_fd_sc_hd__dfxtp_1
X_17458_ _32893_/Q _32829_/Q _32765_/Q _32701_/Q _17346_/X _17347_/X VGND VGND VPWR
+ VPWR _17458_/X sky130_fd_sc_hd__mux4_1
XFILLER_20_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16409_ _34655_/Q _34591_/Q _34527_/Q _34463_/Q _16233_/X _16234_/X VGND VGND VPWR
+ VPWR _16409_/X sky130_fd_sc_hd__mux4_1
XFILLER_203_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35243_ _35433_/CLK _35243_/D VGND VGND VPWR VPWR _35243_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_347_CLK clkbuf_6_47__f_CLK/X VGND VGND VPWR VPWR _35903_/CLK sky130_fd_sc_hd__clkbuf_16
X_32455_ _36085_/CLK _32455_/D VGND VGND VPWR VPWR _32455_/Q sky130_fd_sc_hd__dfxtp_1
X_17389_ _35707_/Q _32216_/Q _35579_/Q _35515_/Q _17317_/X _17318_/X VGND VGND VPWR
+ VPWR _17389_/X sky130_fd_sc_hd__mux4_1
XFILLER_186_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31406_ _27822_/X _35920_/Q _31408_/S VGND VGND VPWR VPWR _31407_/A sky130_fd_sc_hd__mux2_1
X_19128_ _19014_/X _19126_/X _19127_/X _19018_/X VGND VGND VPWR VPWR _19128_/X sky130_fd_sc_hd__a22o_1
XFILLER_145_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35174_ _35625_/CLK _35174_/D VGND VGND VPWR VPWR _35174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32386_ _35970_/CLK _32386_/D VGND VGND VPWR VPWR _32386_/Q sky130_fd_sc_hd__dfxtp_1
X_34125_ _34193_/CLK _34125_/D VGND VGND VPWR VPWR _34125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19059_ _33065_/Q _32041_/Q _35817_/Q _35753_/Q _19025_/X _19026_/X VGND VGND VPWR
+ VPWR _19059_/X sky130_fd_sc_hd__mux4_1
X_31337_ _27720_/X _35887_/Q _31345_/S VGND VGND VPWR VPWR _31338_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34056_ _34121_/CLK _34056_/D VGND VGND VPWR VPWR _34056_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22070_ _21753_/X _22068_/X _22069_/X _21756_/X VGND VGND VPWR VPWR _22070_/X sky130_fd_sc_hd__a22o_1
X_31268_ _31268_/A VGND VGND VPWR VPWR _35854_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21021_ _22399_/A VGND VGND VPWR VPWR _21021_/X sky130_fd_sc_hd__buf_4
X_33007_ _36015_/CLK _33007_/D VGND VGND VPWR VPWR _33007_/Q sky130_fd_sc_hd__dfxtp_1
X_30219_ _30219_/A VGND VGND VPWR VPWR _35357_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31199_ _31199_/A VGND VGND VPWR VPWR _35821_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_248_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25760_ _24920_/X _33341_/Q _25760_/S VGND VGND VPWR VPWR _25761_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22972_ _22971_/X _32049_/Q _22978_/S VGND VGND VPWR VPWR _22973_/A sky130_fd_sc_hd__mux2_1
X_34958_ _34961_/CLK _34958_/D VGND VGND VPWR VPWR _34958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_880 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24711_ _22959_/X _32877_/Q _24723_/S VGND VGND VPWR VPWR _24712_/A sky130_fd_sc_hd__mux2_1
X_33909_ _34100_/CLK _33909_/D VGND VGND VPWR VPWR _33909_/Q sky130_fd_sc_hd__dfxtp_1
X_21923_ _33081_/Q _32057_/Q _35833_/Q _35769_/Q _21678_/X _21679_/X VGND VGND VPWR
+ VPWR _21923_/X sky130_fd_sc_hd__mux4_1
XFILLER_228_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25691_ _24818_/X _33308_/Q _25697_/S VGND VGND VPWR VPWR _25692_/A sky130_fd_sc_hd__mux2_1
X_34889_ _34954_/CLK _34889_/D VGND VGND VPWR VPWR _34889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27430_ _27430_/A VGND VGND VPWR VPWR _34098_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21854_ _22560_/A VGND VGND VPWR VPWR _21854_/X sky130_fd_sc_hd__buf_6
X_24642_ _24642_/A VGND VGND VPWR VPWR _32844_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20805_ _34905_/Q _34841_/Q _34777_/Q _34713_/Q _20696_/X _20698_/X VGND VGND VPWR
+ VPWR _20805_/X sky130_fd_sc_hd__mux4_1
XFILLER_243_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27361_ _34066_/Q _27220_/X _27367_/S VGND VGND VPWR VPWR _27362_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24573_ _24573_/A VGND VGND VPWR VPWR _32811_/D sky130_fd_sc_hd__clkbuf_1
X_21785_ _21598_/X _21783_/X _21784_/X _21601_/X VGND VGND VPWR VPWR _21785_/X sky130_fd_sc_hd__a22o_1
XFILLER_180_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29100_ _29100_/A VGND VGND VPWR VPWR _34857_/D sky130_fd_sc_hd__clkbuf_1
X_26312_ _26312_/A VGND VGND VPWR VPWR _33602_/D sky130_fd_sc_hd__clkbuf_1
X_20736_ _20691_/X _20734_/X _20735_/X _20701_/X VGND VGND VPWR VPWR _20736_/X sky130_fd_sc_hd__a22o_1
X_23524_ _32257_/Q _23432_/X _23536_/S VGND VGND VPWR VPWR _23525_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27292_ _34033_/Q _27118_/X _27296_/S VGND VGND VPWR VPWR _27293_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29031_ _29031_/A VGND VGND VPWR VPWR _34824_/D sky130_fd_sc_hd__clkbuf_1
X_23455_ _32230_/Q _23453_/X _23485_/S VGND VGND VPWR VPWR _23456_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26243_ _26243_/A VGND VGND VPWR VPWR _33569_/D sky130_fd_sc_hd__clkbuf_1
X_20667_ _22535_/A VGND VGND VPWR VPWR _20667_/X sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_338_CLK clkbuf_6_45__f_CLK/X VGND VGND VPWR VPWR _32890_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_109_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22406_ _22402_/X _22405_/X _22085_/X VGND VGND VPWR VPWR _22428_/A sky130_fd_sc_hd__o21ba_1
XFILLER_167_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26174_ _24933_/X _33537_/Q _26186_/S VGND VGND VPWR VPWR _26175_/A sky130_fd_sc_hd__mux2_1
X_23386_ _23386_/A VGND VGND VPWR VPWR _32207_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20598_ input73/X input74/X VGND VGND VPWR VPWR _20599_/A sky130_fd_sc_hd__and2_1
XFILLER_221_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25125_ _25125_/A VGND VGND VPWR VPWR _33042_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22337_ _22012_/X _22335_/X _22336_/X _22018_/X VGND VGND VPWR VPWR _22337_/X sky130_fd_sc_hd__a22o_1
XFILLER_104_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29933_ _30065_/S VGND VGND VPWR VPWR _29952_/S sky130_fd_sc_hd__buf_6
X_25056_ _25056_/A VGND VGND VPWR VPWR _33009_/D sky130_fd_sc_hd__clkbuf_1
X_22268_ _22020_/X _22266_/X _22267_/X _22024_/X VGND VGND VPWR VPWR _22268_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24007_ _22925_/X _32546_/Q _24021_/S VGND VGND VPWR VPWR _24008_/A sky130_fd_sc_hd__mux2_1
X_21219_ _21215_/X _21218_/X _21045_/X VGND VGND VPWR VPWR _21227_/C sky130_fd_sc_hd__o21ba_1
X_29864_ _35189_/Q _29426_/X _29880_/S VGND VGND VPWR VPWR _29865_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_807 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22199_ _22012_/X _22197_/X _22198_/X _22018_/X VGND VGND VPWR VPWR _22199_/X sky130_fd_sc_hd__a22o_1
XFILLER_120_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28815_ _34722_/Q _27072_/X _28829_/S VGND VGND VPWR VPWR _28816_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29795_ _35157_/Q _29524_/X _29795_/S VGND VGND VPWR VPWR _29796_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28746_ _28746_/A VGND VGND VPWR VPWR _34690_/D sky130_fd_sc_hd__clkbuf_1
X_16760_ _16650_/X _16758_/X _16759_/X _16653_/X VGND VGND VPWR VPWR _16760_/X sky130_fd_sc_hd__a22o_1
XFILLER_59_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25958_ _25958_/A VGND VGND VPWR VPWR _33434_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24909_ _24908_/X _32953_/Q _24921_/S VGND VGND VPWR VPWR _24910_/A sky130_fd_sc_hd__mux2_1
X_16691_ _35175_/Q _35111_/Q _35047_/Q _32167_/Q _16657_/X _16658_/X VGND VGND VPWR
+ VPWR _16691_/X sky130_fd_sc_hd__mux4_1
X_28677_ _28677_/A VGND VGND VPWR VPWR _34657_/D sky130_fd_sc_hd__clkbuf_1
X_25889_ _24911_/X _33402_/Q _25895_/S VGND VGND VPWR VPWR _25890_/A sky130_fd_sc_hd__mux2_1
XFILLER_206_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18430_ _18426_/X _18429_/X _18375_/X VGND VGND VPWR VPWR _18438_/C sky130_fd_sc_hd__o21ba_1
XFILLER_189_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27628_ _27628_/A VGND VGND VPWR VPWR _34192_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_206_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18361_ _18361_/A VGND VGND VPWR VPWR _20150_/A sky130_fd_sc_hd__buf_12
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27559_ _27559_/A VGND VGND VPWR VPWR _34159_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17312_ _17059_/X _17310_/X _17311_/X _17065_/X VGND VGND VPWR VPWR _17312_/X sky130_fd_sc_hd__a22o_1
XFILLER_15_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30570_ _35524_/Q _29472_/X _30576_/S VGND VGND VPWR VPWR _30571_/A sky130_fd_sc_hd__mux2_1
X_18292_ _18361_/A VGND VGND VPWR VPWR _20099_/A sky130_fd_sc_hd__buf_12
XFILLER_15_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17243_ _17239_/X _17242_/X _17132_/X VGND VGND VPWR VPWR _17267_/A sky130_fd_sc_hd__o21ba_1
X_29229_ _29229_/A VGND VGND VPWR VPWR _34918_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_329_CLK clkbuf_6_38__f_CLK/X VGND VGND VPWR VPWR _35956_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_175_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32240_ _35729_/CLK _32240_/D VGND VGND VPWR VPWR _32240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17174_ _16853_/X _17172_/X _17173_/X _16856_/X VGND VGND VPWR VPWR _17174_/X sky130_fd_sc_hd__a22o_1
X_16125_ _35607_/Q _34967_/Q _34327_/Q _33687_/Q _16053_/X _16055_/X VGND VGND VPWR
+ VPWR _16125_/X sky130_fd_sc_hd__mux4_1
XFILLER_143_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32171_ _35754_/CLK _32171_/D VGND VGND VPWR VPWR _32171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31122_ _31122_/A VGND VGND VPWR VPWR _35785_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16056_ _35606_/Q _34966_/Q _34326_/Q _33686_/Q _16053_/X _16055_/X VGND VGND VPWR
+ VPWR _16056_/X sky130_fd_sc_hd__mux4_1
XFILLER_97_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35930_ _36055_/CLK _35930_/D VGND VGND VPWR VPWR _35930_/Q sky130_fd_sc_hd__dfxtp_1
X_31053_ _35753_/Q input11/X _31053_/S VGND VGND VPWR VPWR _31054_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_501_CLK clkbuf_6_2__f_CLK/X VGND VGND VPWR VPWR _36068_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_97_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30004_ _30004_/A VGND VGND VPWR VPWR _35255_/D sky130_fd_sc_hd__clkbuf_1
X_19815_ _34942_/Q _34878_/Q _34814_/Q _34750_/Q _19813_/X _19814_/X VGND VGND VPWR
+ VPWR _19815_/X sky130_fd_sc_hd__mux4_1
XFILLER_29_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35861_ _35861_/CLK _35861_/D VGND VGND VPWR VPWR _35861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_1270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34812_ _34941_/CLK _34812_/D VGND VGND VPWR VPWR _34812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19746_ _20260_/A VGND VGND VPWR VPWR _19746_/X sky130_fd_sc_hd__buf_8
X_16958_ _33135_/Q _36015_/Q _33007_/Q _32943_/Q _16709_/X _16710_/X VGND VGND VPWR
+ VPWR _16958_/X sky130_fd_sc_hd__mux4_1
X_35792_ _35855_/CLK _35792_/D VGND VGND VPWR VPWR _35792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31955_ _31955_/A VGND VGND VPWR VPWR _36180_/D sky130_fd_sc_hd__clkbuf_1
X_19677_ _20150_/A VGND VGND VPWR VPWR _19677_/X sky130_fd_sc_hd__buf_8
XFILLER_42_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34743_ _36151_/CLK _34743_/D VGND VGND VPWR VPWR _34743_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16889_ _16853_/X _16887_/X _16888_/X _16856_/X VGND VGND VPWR VPWR _16889_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18628_ _18330_/X _18626_/X _18627_/X _18341_/X VGND VGND VPWR VPWR _18628_/X sky130_fd_sc_hd__a22o_1
X_30906_ _35683_/Q input5/X _30918_/S VGND VGND VPWR VPWR _30907_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34674_ _35377_/CLK _34674_/D VGND VGND VPWR VPWR _34674_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31886_ _31886_/A VGND VGND VPWR VPWR _36147_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_213_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33625_ _34009_/CLK _33625_/D VGND VGND VPWR VPWR _33625_/Q sky130_fd_sc_hd__dfxtp_1
X_30837_ _30837_/A VGND VGND VPWR VPWR _35650_/D sky130_fd_sc_hd__clkbuf_1
X_18559_ _20100_/A VGND VGND VPWR VPWR _18559_/X sky130_fd_sc_hd__buf_4
X_33556_ _33685_/CLK _33556_/D VGND VGND VPWR VPWR _33556_/Q sky130_fd_sc_hd__dfxtp_1
X_21570_ _33071_/Q _32047_/Q _35823_/Q _35759_/Q _21325_/X _21326_/X VGND VGND VPWR
+ VPWR _21570_/X sky130_fd_sc_hd__mux4_1
X_30768_ _30768_/A VGND VGND VPWR VPWR _35617_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_1096 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20521_ _18318_/X _20519_/X _20520_/X _18327_/X VGND VGND VPWR VPWR _20521_/X sky130_fd_sc_hd__a22o_1
XFILLER_20_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32507_ _36027_/CLK _32507_/D VGND VGND VPWR VPWR _32507_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33487_ _34441_/CLK _33487_/D VGND VGND VPWR VPWR _33487_/Q sky130_fd_sc_hd__dfxtp_1
X_30699_ _35585_/Q _29463_/X _30711_/S VGND VGND VPWR VPWR _30700_/A sky130_fd_sc_hd__mux2_1
XFILLER_197_1107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23240_ input34/X VGND VGND VPWR VPWR _23240_/X sky130_fd_sc_hd__buf_4
X_20452_ _20159_/X _20450_/X _20451_/X _20162_/X VGND VGND VPWR VPWR _20452_/X sky130_fd_sc_hd__a22o_1
X_35226_ _35674_/CLK _35226_/D VGND VGND VPWR VPWR _35226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32438_ _33895_/CLK _32438_/D VGND VGND VPWR VPWR _32438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35157_ _35221_/CLK _35157_/D VGND VGND VPWR VPWR _35157_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23171_ _23005_/X _32124_/Q _23173_/S VGND VGND VPWR VPWR _23172_/A sky130_fd_sc_hd__mux2_1
X_20383_ _35727_/Q _32238_/Q _35599_/Q _35535_/Q _18293_/X _18295_/X VGND VGND VPWR
+ VPWR _20383_/X sky130_fd_sc_hd__mux4_1
XFILLER_118_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32369_ _35953_/CLK _32369_/D VGND VGND VPWR VPWR _32369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34108_ _34877_/CLK _34108_/D VGND VGND VPWR VPWR _34108_/Q sky130_fd_sc_hd__dfxtp_1
X_22122_ _33663_/Q _33599_/Q _33535_/Q _33471_/Q _21800_/X _21801_/X VGND VGND VPWR
+ VPWR _22122_/X sky130_fd_sc_hd__mux4_1
XFILLER_12_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35088_ _35217_/CLK _35088_/D VGND VGND VPWR VPWR _35088_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput130 _32004_/Q VGND VGND VPWR VPWR D1[46] sky130_fd_sc_hd__buf_2
XFILLER_216_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput141 _32014_/Q VGND VGND VPWR VPWR D1[56] sky130_fd_sc_hd__buf_2
XTAP_6507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput152 _31966_/Q VGND VGND VPWR VPWR D1[8] sky130_fd_sc_hd__buf_2
XTAP_6518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput163 _36200_/Q VGND VGND VPWR VPWR D2[18] sky130_fd_sc_hd__buf_2
X_34039_ _35703_/CLK _34039_/D VGND VGND VPWR VPWR _34039_/Q sky130_fd_sc_hd__dfxtp_1
X_26930_ _26930_/A VGND VGND VPWR VPWR _33892_/D sky130_fd_sc_hd__clkbuf_1
X_22053_ _22049_/X _22052_/X _21732_/X VGND VGND VPWR VPWR _22075_/A sky130_fd_sc_hd__o21ba_1
XTAP_6529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput174 _36210_/Q VGND VGND VPWR VPWR D2[28] sky130_fd_sc_hd__buf_2
XFILLER_47_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput185 _36220_/Q VGND VGND VPWR VPWR D2[38] sky130_fd_sc_hd__buf_2
XTAP_5806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput196 _36230_/Q VGND VGND VPWR VPWR D2[48] sky130_fd_sc_hd__buf_2
X_21004_ _20892_/X _21002_/X _21003_/X _20895_/X VGND VGND VPWR VPWR _21004_/X sky130_fd_sc_hd__a22o_1
XFILLER_43_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26861_ _33860_/Q _23441_/X _26867_/S VGND VGND VPWR VPWR _26862_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28600_ _28648_/S VGND VGND VPWR VPWR _28619_/S sky130_fd_sc_hd__buf_4
XFILLER_102_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25812_ _28110_/A _26352_/B VGND VGND VPWR VPWR _25945_/S sky130_fd_sc_hd__nand2_8
XFILLER_75_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_997 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29580_ _29580_/A VGND VGND VPWR VPWR _35054_/D sky130_fd_sc_hd__clkbuf_1
X_26792_ _33827_/Q _23271_/X _26804_/S VGND VGND VPWR VPWR _26793_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28531_ _27664_/X _34589_/Q _28535_/S VGND VGND VPWR VPWR _28532_/A sky130_fd_sc_hd__mux2_1
X_25743_ _25743_/A VGND VGND VPWR VPWR _33332_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22955_ _22955_/A VGND VGND VPWR VPWR _32043_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21906_ _33401_/Q _33337_/Q _33273_/Q _33209_/Q _21727_/X _21728_/X VGND VGND VPWR
+ VPWR _21906_/X sky130_fd_sc_hd__mux4_1
X_28462_ _28462_/A VGND VGND VPWR VPWR _34556_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25674_ _25674_/A VGND VGND VPWR VPWR _33300_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_216_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22886_ _31147_/A _30202_/A VGND VGND VPWR VPWR _22887_/A sky130_fd_sc_hd__or2_1
XFILLER_216_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27413_ _34090_/Q _27096_/X _27431_/S VGND VGND VPWR VPWR _27414_/A sky130_fd_sc_hd__mux2_1
X_24625_ _24625_/A VGND VGND VPWR VPWR _32836_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28393_ _28393_/A VGND VGND VPWR VPWR _34523_/D sky130_fd_sc_hd__clkbuf_1
X_21837_ _33655_/Q _33591_/Q _33527_/Q _33463_/Q _21800_/X _21801_/X VGND VGND VPWR
+ VPWR _21837_/X sky130_fd_sc_hd__mux4_1
XFILLER_58_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27344_ _27344_/A VGND VGND VPWR VPWR _34057_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24556_ _24556_/A VGND VGND VPWR VPWR _32803_/D sky130_fd_sc_hd__clkbuf_1
X_21768_ _21768_/A VGND VGND VPWR VPWR _36212_/D sky130_fd_sc_hd__buf_6
XFILLER_15_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20719_ _20618_/X _20717_/X _20718_/X _20627_/X VGND VGND VPWR VPWR _20719_/X sky130_fd_sc_hd__a22o_1
XFILLER_145_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23507_ _32249_/Q _23405_/X _23515_/S VGND VGND VPWR VPWR _23508_/A sky130_fd_sc_hd__mux2_1
X_27275_ _34025_/Q _27093_/X _27275_/S VGND VGND VPWR VPWR _27276_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24487_ _23027_/X _32771_/Q _24495_/S VGND VGND VPWR VPWR _24488_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21699_ _21453_/X _21697_/X _21698_/X _21456_/X VGND VGND VPWR VPWR _21699_/X sky130_fd_sc_hd__a22o_1
XFILLER_8_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_838 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29014_ _29014_/A VGND VGND VPWR VPWR _34816_/D sky130_fd_sc_hd__clkbuf_1
X_26226_ _26226_/A VGND VGND VPWR VPWR _33561_/D sky130_fd_sc_hd__clkbuf_1
X_23438_ input40/X VGND VGND VPWR VPWR _23438_/X sky130_fd_sc_hd__buf_4
XFILLER_149_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26157_ _24908_/X _33529_/Q _26165_/S VGND VGND VPWR VPWR _26158_/A sky130_fd_sc_hd__mux2_1
X_23369_ _32200_/Q _23299_/X _23385_/S VGND VGND VPWR VPWR _23370_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25108_ _24961_/X _33034_/Q _25122_/S VGND VGND VPWR VPWR _25109_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26088_ _24806_/X _33496_/Q _26102_/S VGND VGND VPWR VPWR _26089_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17930_ _17709_/X _17928_/X _17929_/X _17712_/X VGND VGND VPWR VPWR _17930_/X sky130_fd_sc_hd__a22o_1
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29916_ _35214_/Q _29503_/X _29922_/S VGND VGND VPWR VPWR _29917_/A sky130_fd_sc_hd__mux2_1
X_25039_ _25039_/A VGND VGND VPWR VPWR _33001_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17861_ _35208_/Q _35144_/Q _35080_/Q _32264_/Q _17716_/X _17717_/X VGND VGND VPWR
+ VPWR _17861_/X sky130_fd_sc_hd__mux4_1
XFILLER_121_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29847_ _35181_/Q _29401_/X _29859_/S VGND VGND VPWR VPWR _29848_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19600_ _19596_/X _19599_/X _19465_/X VGND VGND VPWR VPWR _19601_/D sky130_fd_sc_hd__o21ba_1
X_16812_ _17871_/A VGND VGND VPWR VPWR _16812_/X sky130_fd_sc_hd__buf_2
XFILLER_120_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17792_ _34438_/Q _36166_/Q _34310_/Q _34246_/Q _17582_/X _17583_/X VGND VGND VPWR
+ VPWR _17792_/X sky130_fd_sc_hd__mux4_1
X_29778_ _29778_/A VGND VGND VPWR VPWR _35148_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19531_ _34422_/Q _36150_/Q _34294_/Q _34230_/Q _19529_/X _19530_/X VGND VGND VPWR
+ VPWR _19531_/X sky130_fd_sc_hd__mux4_1
XFILLER_207_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16743_ _16493_/X _16739_/X _16742_/X _16498_/X VGND VGND VPWR VPWR _16743_/X sky130_fd_sc_hd__a22o_1
X_28729_ _28729_/A VGND VGND VPWR VPWR _34682_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_1063 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31740_ _36078_/Q input17/X _31750_/S VGND VGND VPWR VPWR _31741_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19462_ _34932_/Q _34868_/Q _34804_/Q _34740_/Q _19460_/X _19461_/X VGND VGND VPWR
+ VPWR _19462_/X sky130_fd_sc_hd__mux4_1
XFILLER_185_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16674_ _16500_/X _16670_/X _16673_/X _16503_/X VGND VGND VPWR VPWR _16674_/X sky130_fd_sc_hd__a22o_1
XFILLER_74_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18413_ _20151_/A VGND VGND VPWR VPWR _18413_/X sky130_fd_sc_hd__buf_4
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31671_ _31671_/A VGND VGND VPWR VPWR _36045_/D sky130_fd_sc_hd__clkbuf_1
X_19393_ _20260_/A VGND VGND VPWR VPWR _19393_/X sky130_fd_sc_hd__buf_4
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33410_ _36097_/CLK _33410_/D VGND VGND VPWR VPWR _33410_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30622_ _30622_/A VGND VGND VPWR VPWR _35548_/D sky130_fd_sc_hd__clkbuf_1
X_18344_ _20146_/A VGND VGND VPWR VPWR _18344_/X sky130_fd_sc_hd__buf_4
X_34390_ _34647_/CLK _34390_/D VGND VGND VPWR VPWR _34390_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33341_ _36092_/CLK _33341_/D VGND VGND VPWR VPWR _33341_/Q sky130_fd_sc_hd__dfxtp_1
X_18275_ _16060_/X _18273_/X _18274_/X _16072_/X VGND VGND VPWR VPWR _18275_/X sky130_fd_sc_hd__a22o_1
XFILLER_175_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30553_ _35516_/Q _29447_/X _30555_/S VGND VGND VPWR VPWR _30554_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36060_ _36060_/CLK _36060_/D VGND VGND VPWR VPWR _36060_/Q sky130_fd_sc_hd__dfxtp_1
X_17226_ _34678_/Q _34614_/Q _34550_/Q _34486_/Q _16939_/X _16940_/X VGND VGND VPWR
+ VPWR _17226_/X sky130_fd_sc_hd__mux4_1
XFILLER_200_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput10 DW[18] VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__buf_6
X_33272_ _33911_/CLK _33272_/D VGND VGND VPWR VPWR _33272_/Q sky130_fd_sc_hd__dfxtp_1
X_30484_ _35483_/Q _29345_/X _30492_/S VGND VGND VPWR VPWR _30485_/A sky130_fd_sc_hd__mux2_1
Xinput21 DW[28] VGND VGND VPWR VPWR input21/X sky130_fd_sc_hd__buf_4
XFILLER_156_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput32 DW[38] VGND VGND VPWR VPWR input32/X sky130_fd_sc_hd__clkbuf_8
XFILLER_174_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35011_ _35651_/CLK _35011_/D VGND VGND VPWR VPWR _35011_/Q sky130_fd_sc_hd__dfxtp_1
Xinput43 DW[48] VGND VGND VPWR VPWR input43/X sky130_fd_sc_hd__buf_8
X_32223_ _35711_/CLK _32223_/D VGND VGND VPWR VPWR _32223_/Q sky130_fd_sc_hd__dfxtp_1
Xinput54 DW[58] VGND VGND VPWR VPWR input54/X sky130_fd_sc_hd__buf_12
X_17157_ _17153_/X _17154_/X _17155_/X _17156_/X VGND VGND VPWR VPWR _17157_/X sky130_fd_sc_hd__a22o_1
Xinput65 R1[0] VGND VGND VPWR VPWR input65/X sky130_fd_sc_hd__clkbuf_2
Xinput76 R2[5] VGND VGND VPWR VPWR input76/X sky130_fd_sc_hd__clkbuf_4
Xinput87 RW[4] VGND VGND VPWR VPWR input87/X sky130_fd_sc_hd__buf_4
X_16108_ _33623_/Q _33559_/Q _33495_/Q _33431_/Q _15984_/X _15987_/X VGND VGND VPWR
+ VPWR _16108_/X sky130_fd_sc_hd__mux4_1
X_32154_ _36127_/CLK _32154_/D VGND VGND VPWR VPWR _32154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17088_ _16805_/X _17086_/X _17087_/X _16810_/X VGND VGND VPWR VPWR _17088_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31105_ _31105_/A VGND VGND VPWR VPWR _35777_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16039_ _17834_/A VGND VGND VPWR VPWR _16039_/X sky130_fd_sc_hd__buf_4
XFILLER_130_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32085_ _36052_/CLK _32085_/D VGND VGND VPWR VPWR _32085_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_30_CLK clkbuf_6_5__f_CLK/X VGND VGND VPWR VPWR _36207_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_112_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35913_ _35978_/CLK _35913_/D VGND VGND VPWR VPWR _35913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31036_ _31036_/A VGND VGND VPWR VPWR _35744_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35844_ _36038_/CLK _35844_/D VGND VGND VPWR VPWR _35844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_244_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_6_59__f_CLK clkbuf_5_29_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_59__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_19729_ _19651_/X _19727_/X _19728_/X _19654_/X VGND VGND VPWR VPWR _19729_/X sky130_fd_sc_hd__a22o_1
X_32987_ _36055_/CLK _32987_/D VGND VGND VPWR VPWR _32987_/Q sky130_fd_sc_hd__dfxtp_1
X_35775_ _35839_/CLK _35775_/D VGND VGND VPWR VPWR _35775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22740_ _32913_/Q _32849_/Q _32785_/Q _32721_/Q _20584_/X _20587_/X VGND VGND VPWR
+ VPWR _22740_/X sky130_fd_sc_hd__mux4_1
X_34726_ _34790_/CLK _34726_/D VGND VGND VPWR VPWR _34726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31938_ _23469_/X _36172_/Q _31948_/S VGND VGND VPWR VPWR _31939_/A sky130_fd_sc_hd__mux2_1
XFILLER_225_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22671_ _22505_/X _22669_/X _22670_/X _22510_/X VGND VGND VPWR VPWR _22671_/X sky130_fd_sc_hd__a22o_1
XFILLER_129_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31869_ _23296_/X _36139_/Q _31885_/S VGND VGND VPWR VPWR _31870_/A sky130_fd_sc_hd__mux2_1
X_34657_ _35297_/CLK _34657_/D VGND VGND VPWR VPWR _34657_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_97_CLK clkbuf_leaf_99_CLK/A VGND VGND VPWR VPWR _36058_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_40_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24410_ _24410_/A VGND VGND VPWR VPWR _32734_/D sky130_fd_sc_hd__clkbuf_1
X_21622_ _21446_/X _21620_/X _21621_/X _21451_/X VGND VGND VPWR VPWR _21622_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33608_ _33673_/CLK _33608_/D VGND VGND VPWR VPWR _33608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25390_ _25390_/A VGND VGND VPWR VPWR _33166_/D sky130_fd_sc_hd__clkbuf_1
X_34588_ _36229_/CLK _34588_/D VGND VGND VPWR VPWR _34588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24341_ _24389_/S VGND VGND VPWR VPWR _24360_/S sky130_fd_sc_hd__buf_4
X_21553_ _33391_/Q _33327_/Q _33263_/Q _33199_/Q _21374_/X _21375_/X VGND VGND VPWR
+ VPWR _21553_/X sky130_fd_sc_hd__mux4_1
X_33539_ _34942_/CLK _33539_/D VGND VGND VPWR VPWR _33539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_945 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20504_ _35667_/Q _35027_/Q _34387_/Q _33747_/Q _18412_/X _18413_/X VGND VGND VPWR
+ VPWR _20504_/X sky130_fd_sc_hd__mux4_1
X_27060_ _33950_/Q _27059_/X _27063_/S VGND VGND VPWR VPWR _27061_/A sky130_fd_sc_hd__mux2_1
X_24272_ _22909_/X _32669_/Q _24276_/S VGND VGND VPWR VPWR _24273_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21484_ _33645_/Q _33581_/Q _33517_/Q _33453_/Q _21447_/X _21448_/X VGND VGND VPWR
+ VPWR _21484_/X sky130_fd_sc_hd__mux4_1
XFILLER_165_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23223_ _23082_/X _32149_/Q _23223_/S VGND VGND VPWR VPWR _23224_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26011_ _26080_/S VGND VGND VPWR VPWR _26030_/S sky130_fd_sc_hd__buf_4
XFILLER_105_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20435_ _20431_/X _20434_/X _20138_/X VGND VGND VPWR VPWR _20457_/A sky130_fd_sc_hd__o21ba_2
X_35209_ _35210_/CLK _35209_/D VGND VGND VPWR VPWR _35209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_883 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36189_ _36205_/CLK _36189_/D VGND VGND VPWR VPWR _36189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23154_ _23223_/S VGND VGND VPWR VPWR _23173_/S sky130_fd_sc_hd__buf_4
XTAP_7005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20366_ _20362_/X _20365_/X _20171_/X VGND VGND VPWR VPWR _20367_/D sky130_fd_sc_hd__o21ba_1
XTAP_7016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_1298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22105_ _22100_/X _22103_/X _22104_/X VGND VGND VPWR VPWR _22120_/C sky130_fd_sc_hd__o21ba_1
XFILLER_122_717 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27962_ _27962_/A VGND VGND VPWR VPWR _34319_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23085_ input88/X input87/X input86/X VGND VGND VPWR VPWR _23086_/A sky130_fd_sc_hd__and3_1
X_20297_ _20293_/X _20296_/X _20157_/X VGND VGND VPWR VPWR _20307_/C sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_21_CLK clkbuf_6_4__f_CLK/X VGND VGND VPWR VPWR _36136_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_6326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29701_ _35112_/Q _29385_/X _29703_/S VGND VGND VPWR VPWR _29702_/A sky130_fd_sc_hd__mux2_1
XTAP_6348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26913_ _26913_/A VGND VGND VPWR VPWR _33884_/D sky130_fd_sc_hd__clkbuf_1
X_22036_ _34684_/Q _34620_/Q _34556_/Q _34492_/Q _21892_/X _21893_/X VGND VGND VPWR
+ VPWR _22036_/X sky130_fd_sc_hd__mux4_1
XTAP_6359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27893_ _27893_/A VGND VGND VPWR VPWR _34286_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29632_ _29632_/A VGND VGND VPWR VPWR _35079_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26844_ _33852_/Q _23414_/X _26846_/S VGND VGND VPWR VPWR _26845_/A sky130_fd_sc_hd__mux2_1
XTAP_5669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29563_ _29563_/A VGND VGND VPWR VPWR _35046_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26775_ _33819_/Q _23246_/X _26783_/S VGND VGND VPWR VPWR _26776_/A sky130_fd_sc_hd__mux2_1
XTAP_4968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23987_ _23987_/A VGND VGND VPWR VPWR _32536_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28514_ _28514_/A VGND VGND VPWR VPWR _34581_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_217_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25726_ _25726_/A VGND VGND VPWR VPWR _33324_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29494_ input49/X VGND VGND VPWR VPWR _29494_/X sky130_fd_sc_hd__buf_2
XFILLER_113_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22938_ _22937_/X _32038_/Q _22947_/S VGND VGND VPWR VPWR _22939_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28445_ _27735_/X _34548_/Q _28463_/S VGND VGND VPWR VPWR _28446_/A sky130_fd_sc_hd__mux2_1
X_25657_ _24967_/X _33292_/Q _25667_/S VGND VGND VPWR VPWR _25658_/A sky130_fd_sc_hd__mux2_1
X_22869_ _22865_/X _22868_/X _22457_/A VGND VGND VPWR VPWR _22877_/C sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_88_CLK clkbuf_leaf_88_CLK/A VGND VGND VPWR VPWR _35677_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_32_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24608_ _24608_/A VGND VGND VPWR VPWR _32828_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28376_ _27834_/X _34516_/Q _28378_/S VGND VGND VPWR VPWR _28377_/A sky130_fd_sc_hd__mux2_1
XPHY_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16390_ _16140_/X _16386_/X _16389_/X _16145_/X VGND VGND VPWR VPWR _16390_/X sky130_fd_sc_hd__a22o_1
XPHY_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25588_ _24865_/X _33259_/Q _25604_/S VGND VGND VPWR VPWR _25589_/A sky130_fd_sc_hd__mux2_1
XFILLER_227_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27327_ _27327_/A VGND VGND VPWR VPWR _34049_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24539_ _24539_/A VGND VGND VPWR VPWR _32795_/D sky130_fd_sc_hd__clkbuf_1
XPHY_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18060_ _34702_/Q _34638_/Q _34574_/Q _34510_/Q _17998_/X _17999_/X VGND VGND VPWR
+ VPWR _18060_/X sky130_fd_sc_hd__mux4_1
XFILLER_89_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27258_ _27258_/A VGND VGND VPWR VPWR _34016_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17011_ _17011_/A VGND VGND VPWR VPWR _17011_/X sky130_fd_sc_hd__clkbuf_4
X_26209_ _24985_/X _33554_/Q _26215_/S VGND VGND VPWR VPWR _26210_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27189_ input46/X VGND VGND VPWR VPWR _27189_/X sky130_fd_sc_hd__buf_4
XFILLER_137_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18962_ _34918_/Q _34854_/Q _34790_/Q _34726_/Q _18754_/X _18755_/X VGND VGND VPWR
+ VPWR _18962_/X sky130_fd_sc_hd__mux4_1
XFILLER_106_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_12_CLK clkbuf_6_3__f_CLK/X VGND VGND VPWR VPWR _36137_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_140_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17913_ _33418_/Q _33354_/Q _33290_/Q _33226_/Q _17833_/X _17834_/X VGND VGND VPWR
+ VPWR _17913_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18893_ _18752_/X _18891_/X _18892_/X _18757_/X VGND VGND VPWR VPWR _18893_/X sky130_fd_sc_hd__a22o_1
XTAP_6860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17844_ _32904_/Q _32840_/Q _32776_/Q _32712_/Q _17699_/X _17700_/X VGND VGND VPWR
+ VPWR _17844_/X sky130_fd_sc_hd__mux4_1
X_32910_ _32911_/CLK _32910_/D VGND VGND VPWR VPWR _32910_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33890_ _36066_/CLK _33890_/D VGND VGND VPWR VPWR _33890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32841_ _32905_/CLK _32841_/D VGND VGND VPWR VPWR _32841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17775_ _32134_/Q _32326_/Q _32390_/Q _35910_/Q _17633_/X _17774_/X VGND VGND VPWR
+ VPWR _17775_/X sky130_fd_sc_hd__mux4_1
XFILLER_82_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16726_ _17936_/A VGND VGND VPWR VPWR _16726_/X sky130_fd_sc_hd__buf_4
XFILLER_78_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19514_ _19359_/X _19512_/X _19513_/X _19365_/X VGND VGND VPWR VPWR _19514_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32772_ _35973_/CLK _32772_/D VGND VGND VPWR VPWR _32772_/Q sky130_fd_sc_hd__dfxtp_1
X_35560_ _35560_/CLK _35560_/D VGND VGND VPWR VPWR _35560_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_235_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34511_ _34705_/CLK _34511_/D VGND VGND VPWR VPWR _34511_/Q sky130_fd_sc_hd__dfxtp_1
X_31723_ _36070_/Q input8/X _31729_/S VGND VGND VPWR VPWR _31724_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19445_ _20299_/A VGND VGND VPWR VPWR _19445_/X sky130_fd_sc_hd__buf_4
X_16657_ _17716_/A VGND VGND VPWR VPWR _16657_/X sky130_fd_sc_hd__clkbuf_8
X_35491_ _36135_/CLK _35491_/D VGND VGND VPWR VPWR _35491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_79_CLK clkbuf_leaf_81_CLK/A VGND VGND VPWR VPWR _36055_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_223_868 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34442_ _36171_/CLK _34442_/D VGND VGND VPWR VPWR _34442_/Q sky130_fd_sc_hd__dfxtp_1
X_31654_ _31654_/A VGND VGND VPWR VPWR _36037_/D sky130_fd_sc_hd__clkbuf_1
X_19376_ _19298_/X _19374_/X _19375_/X _19301_/X VGND VGND VPWR VPWR _19376_/X sky130_fd_sc_hd__a22o_1
X_16588_ _34660_/Q _34596_/Q _34532_/Q _34468_/Q _16586_/X _16587_/X VGND VGND VPWR
+ VPWR _16588_/X sky130_fd_sc_hd__mux4_1
XFILLER_163_1150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18327_ _20210_/A VGND VGND VPWR VPWR _18327_/X sky130_fd_sc_hd__buf_4
X_30605_ _35541_/Q _29524_/X _30605_/S VGND VGND VPWR VPWR _30606_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34373_ _35717_/CLK _34373_/D VGND VGND VPWR VPWR _34373_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31585_ _31585_/A VGND VGND VPWR VPWR _36004_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_206_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36112_ _36113_/CLK _36112_/D VGND VGND VPWR VPWR _36112_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33324_ _36076_/CLK _33324_/D VGND VGND VPWR VPWR _33324_/Q sky130_fd_sc_hd__dfxtp_1
X_18258_ _17153_/A _18256_/X _18257_/X _17156_/A VGND VGND VPWR VPWR _18258_/X sky130_fd_sc_hd__a22o_1
X_30536_ _30605_/S VGND VGND VPWR VPWR _30555_/S sky130_fd_sc_hd__buf_6
XFILLER_204_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17209_ _17915_/A VGND VGND VPWR VPWR _17209_/X sky130_fd_sc_hd__buf_6
XFILLER_191_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36043_ _36044_/CLK _36043_/D VGND VGND VPWR VPWR _36043_/Q sky130_fd_sc_hd__dfxtp_1
X_33255_ _36072_/CLK _33255_/D VGND VGND VPWR VPWR _33255_/Q sky130_fd_sc_hd__dfxtp_1
X_18189_ _33683_/Q _33619_/Q _33555_/Q _33491_/Q _17906_/X _17907_/X VGND VGND VPWR
+ VPWR _18189_/X sky130_fd_sc_hd__mux4_1
X_30467_ _30467_/A VGND VGND VPWR VPWR _35475_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20220_ _20065_/X _20218_/X _20219_/X _20071_/X VGND VGND VPWR VPWR _20220_/X sky130_fd_sc_hd__a22o_1
XFILLER_116_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32206_ _35699_/CLK _32206_/D VGND VGND VPWR VPWR _32206_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33186_ _33827_/CLK _33186_/D VGND VGND VPWR VPWR _33186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30398_ _30398_/A VGND VGND VPWR VPWR _35442_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20151_ _20151_/A VGND VGND VPWR VPWR _20151_/X sky130_fd_sc_hd__clkbuf_4
X_32137_ _35976_/CLK _32137_/D VGND VGND VPWR VPWR _32137_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20082_ _20004_/X _20080_/X _20081_/X _20007_/X VGND VGND VPWR VPWR _20082_/X sky130_fd_sc_hd__a22o_1
X_32068_ _36038_/CLK _32068_/D VGND VGND VPWR VPWR _32068_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31019_ _31019_/A VGND VGND VPWR VPWR _35736_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23910_ _23910_/A VGND VGND VPWR VPWR _32500_/D sky130_fd_sc_hd__clkbuf_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24890_ _24889_/X _32947_/Q _24890_/S VGND VGND VPWR VPWR _24891_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_245_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23841_ _23841_/A VGND VGND VPWR VPWR _32405_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35827_ _36147_/CLK _35827_/D VGND VGND VPWR VPWR _35827_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26560_ _24902_/X _33719_/Q _26572_/S VGND VGND VPWR VPWR _26561_/A sky130_fd_sc_hd__mux2_1
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20984_ _20984_/A _20984_/B _20984_/C _20984_/D VGND VGND VPWR VPWR _20985_/A sky130_fd_sc_hd__or4_1
X_35758_ _35822_/CLK _35758_/D VGND VGND VPWR VPWR _35758_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23772_ _22980_/X _32372_/Q _23790_/S VGND VGND VPWR VPWR _23773_/A sky130_fd_sc_hd__mux2_1
XFILLER_226_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25511_ _24951_/X _33223_/Q _25511_/S VGND VGND VPWR VPWR _25512_/A sky130_fd_sc_hd__mux2_1
X_22723_ _34448_/Q _36176_/Q _34320_/Q _34256_/Q _22535_/X _22536_/X VGND VGND VPWR
+ VPWR _22723_/X sky130_fd_sc_hd__mux4_1
X_34709_ _36117_/CLK _34709_/D VGND VGND VPWR VPWR _34709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26491_ _24796_/X _33686_/Q _26509_/S VGND VGND VPWR VPWR _26492_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_246_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35689_ _35691_/CLK _35689_/D VGND VGND VPWR VPWR _35689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28230_ _28230_/A VGND VGND VPWR VPWR _34446_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25442_ _24849_/X _33190_/Q _25448_/S VGND VGND VPWR VPWR _25443_/A sky130_fd_sc_hd__mux2_1
XFILLER_241_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22654_ _35662_/Q _35022_/Q _34382_/Q _33742_/Q _22450_/X _22451_/X VGND VGND VPWR
+ VPWR _22654_/X sky130_fd_sc_hd__mux4_1
XFILLER_25_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28161_ _28161_/A VGND VGND VPWR VPWR _34413_/D sky130_fd_sc_hd__clkbuf_1
X_21605_ _33072_/Q _32048_/Q _35824_/Q _35760_/Q _21325_/X _21326_/X VGND VGND VPWR
+ VPWR _21605_/X sky130_fd_sc_hd__mux4_1
XFILLER_230_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25373_ _25373_/A VGND VGND VPWR VPWR _33158_/D sky130_fd_sc_hd__clkbuf_1
X_22585_ _22365_/X _22583_/X _22584_/X _22371_/X VGND VGND VPWR VPWR _22585_/X sky130_fd_sc_hd__a22o_1
XFILLER_107_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27112_ input18/X VGND VGND VPWR VPWR _27112_/X sky130_fd_sc_hd__buf_2
X_24324_ _24324_/A VGND VGND VPWR VPWR _32693_/D sky130_fd_sc_hd__clkbuf_1
X_28092_ _34381_/Q _27205_/X _28100_/S VGND VGND VPWR VPWR _28093_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21536_ _33070_/Q _32046_/Q _35822_/Q _35758_/Q _21325_/X _21326_/X VGND VGND VPWR
+ VPWR _21536_/X sky130_fd_sc_hd__mux4_1
XFILLER_103_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27043_ _27043_/A VGND VGND VPWR VPWR _33944_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24255_ _28786_/A _28786_/B VGND VGND VPWR VPWR _31283_/B sky130_fd_sc_hd__nor2_8
X_21467_ _35628_/Q _34988_/Q _34348_/Q _33708_/Q _21391_/X _21392_/X VGND VGND VPWR
+ VPWR _21467_/X sky130_fd_sc_hd__mux4_1
XFILLER_147_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20418_ _18301_/X _20416_/X _20417_/X _18307_/X VGND VGND VPWR VPWR _20418_/X sky130_fd_sc_hd__a22o_1
X_23206_ _23206_/A VGND VGND VPWR VPWR _32140_/D sky130_fd_sc_hd__clkbuf_1
X_21398_ _22457_/A VGND VGND VPWR VPWR _21398_/X sky130_fd_sc_hd__buf_2
X_24186_ _24186_/A VGND VGND VPWR VPWR _32629_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20349_ _32142_/Q _32334_/Q _32398_/Q _35918_/Q _20286_/X _20074_/X VGND VGND VPWR
+ VPWR _20349_/X sky130_fd_sc_hd__mux4_1
X_23137_ _23137_/A VGND VGND VPWR VPWR _32107_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28994_ _34807_/Q _27137_/X _29006_/S VGND VGND VPWR VPWR _28995_/A sky130_fd_sc_hd__mux2_1
XTAP_6112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27945_ _27945_/A VGND VGND VPWR VPWR _34311_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23068_ _23067_/X _32080_/Q _23071_/S VGND VGND VPWR VPWR _23069_/A sky130_fd_sc_hd__mux2_1
XTAP_6145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_995 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22019_ _22012_/X _22014_/X _22017_/X _22018_/X VGND VGND VPWR VPWR _22019_/X sky130_fd_sc_hd__a22o_1
XTAP_6189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27876_ _27876_/A VGND VGND VPWR VPWR _34278_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29615_ _35071_/Q _29457_/X _29631_/S VGND VGND VPWR VPWR _29616_/A sky130_fd_sc_hd__mux2_1
XTAP_4743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26827_ _26896_/S VGND VGND VPWR VPWR _26846_/S sky130_fd_sc_hd__buf_4
XTAP_5499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_6_42__f_CLK clkbuf_5_21_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_42__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_5_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29546_ _29546_/A VGND VGND VPWR VPWR _35038_/D sky130_fd_sc_hd__clkbuf_1
X_17560_ _33408_/Q _33344_/Q _33280_/Q _33216_/Q _17480_/X _17481_/X VGND VGND VPWR
+ VPWR _17560_/X sky130_fd_sc_hd__mux4_1
XTAP_4787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26758_ _26758_/A VGND VGND VPWR VPWR _33811_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16511_ _16361_/X _16509_/X _16510_/X _16365_/X VGND VGND VPWR VPWR _16511_/X sky130_fd_sc_hd__a22o_1
XFILLER_186_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25709_ _25709_/A VGND VGND VPWR VPWR _33316_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29477_ _29477_/A VGND VGND VPWR VPWR _35013_/D sky130_fd_sc_hd__clkbuf_1
X_17491_ _32894_/Q _32830_/Q _32766_/Q _32702_/Q _17346_/X _17347_/X VGND VGND VPWR
+ VPWR _17491_/X sky130_fd_sc_hd__mux4_1
XFILLER_232_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26689_ _26689_/A VGND VGND VPWR VPWR _33778_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19230_ _19014_/X _19228_/X _19229_/X _19018_/X VGND VGND VPWR VPWR _19230_/X sky130_fd_sc_hd__a22o_1
X_28428_ _27711_/X _34540_/Q _28442_/S VGND VGND VPWR VPWR _28429_/A sky130_fd_sc_hd__mux2_1
X_16442_ _35424_/Q _35360_/Q _35296_/Q _35232_/Q _16195_/X _16196_/X VGND VGND VPWR
+ VPWR _16442_/X sky130_fd_sc_hd__mux4_1
XFILLER_108_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_1_CLK clkbuf_leaf_2_CLK/A VGND VGND VPWR VPWR _34146_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19161_ _19006_/X _19159_/X _19160_/X _19012_/X VGND VGND VPWR VPWR _19161_/X sky130_fd_sc_hd__a22o_1
X_28359_ _28359_/A VGND VGND VPWR VPWR _34507_/D sky130_fd_sc_hd__clkbuf_1
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16373_ _17936_/A VGND VGND VPWR VPWR _16373_/X sky130_fd_sc_hd__buf_4
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18112_ _18108_/X _18111_/X _17846_/X _17847_/X VGND VGND VPWR VPWR _18127_/B sky130_fd_sc_hd__o211a_1
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31370_ _31370_/A VGND VGND VPWR VPWR _35902_/D sky130_fd_sc_hd__clkbuf_1
X_19092_ _20299_/A VGND VGND VPWR VPWR _19092_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_76_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18043_ _33934_/Q _33870_/Q _33806_/Q _36110_/Q _17730_/X _17731_/X VGND VGND VPWR
+ VPWR _18043_/X sky130_fd_sc_hd__mux4_1
X_30321_ _35406_/Q _29503_/X _30327_/S VGND VGND VPWR VPWR _30322_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_240_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33040_ _36049_/CLK _33040_/D VGND VGND VPWR VPWR _33040_/Q sky130_fd_sc_hd__dfxtp_1
X_30252_ _35373_/Q _29401_/X _30264_/S VGND VGND VPWR VPWR _30253_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30183_ _30183_/A VGND VGND VPWR VPWR _35340_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19994_ _19990_/X _19993_/X _19785_/X VGND VGND VPWR VPWR _20024_/A sky130_fd_sc_hd__o21ba_1
XFILLER_10_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18945_ _20159_/A VGND VGND VPWR VPWR _18945_/X sky130_fd_sc_hd__clkbuf_4
X_34991_ _34991_/CLK _34991_/D VGND VGND VPWR VPWR _34991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33942_ _34070_/CLK _33942_/D VGND VGND VPWR VPWR _33942_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18876_ _32868_/Q _32804_/Q _32740_/Q _32676_/Q _18587_/X _18588_/X VGND VGND VPWR
+ VPWR _18876_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17827_ _17823_/X _17826_/X _17518_/X VGND VGND VPWR VPWR _17828_/D sky130_fd_sc_hd__o21ba_1
X_33873_ _34441_/CLK _33873_/D VGND VGND VPWR VPWR _33873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35612_ _36060_/CLK _35612_/D VGND VGND VPWR VPWR _35612_/Q sky130_fd_sc_hd__dfxtp_1
X_32824_ _32891_/CLK _32824_/D VGND VGND VPWR VPWR _32824_/Q sky130_fd_sc_hd__dfxtp_1
X_17758_ _33670_/Q _33606_/Q _33542_/Q _33478_/Q _17553_/X _17554_/X VGND VGND VPWR
+ VPWR _17758_/X sky130_fd_sc_hd__mux4_1
XFILLER_47_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35543_ _35673_/CLK _35543_/D VGND VGND VPWR VPWR _35543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16709_ _17906_/A VGND VGND VPWR VPWR _16709_/X sky130_fd_sc_hd__buf_4
X_17689_ _34180_/Q _34116_/Q _34052_/Q _33988_/Q _17446_/X _17447_/X VGND VGND VPWR
+ VPWR _17689_/X sky130_fd_sc_hd__mux4_1
XFILLER_120_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32755_ _32906_/CLK _32755_/D VGND VGND VPWR VPWR _32755_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31706_ _36062_/Q input63/X _31708_/S VGND VGND VPWR VPWR _31707_/A sky130_fd_sc_hd__mux2_1
X_19428_ _20134_/A VGND VGND VPWR VPWR _19428_/X sky130_fd_sc_hd__clkbuf_4
X_35474_ _35666_/CLK _35474_/D VGND VGND VPWR VPWR _35474_/Q sky130_fd_sc_hd__dfxtp_1
X_32686_ _32877_/CLK _32686_/D VGND VGND VPWR VPWR _32686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34425_ _36152_/CLK _34425_/D VGND VGND VPWR VPWR _34425_/Q sky130_fd_sc_hd__dfxtp_1
X_31637_ _31637_/A VGND VGND VPWR VPWR _36029_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_241_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19359_ _20205_/A VGND VGND VPWR VPWR _19359_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_50_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22370_ _33158_/Q _36038_/Q _33030_/Q _32966_/Q _22368_/X _22369_/X VGND VGND VPWR
+ VPWR _22370_/X sky130_fd_sc_hd__mux4_1
X_31568_ _31568_/A VGND VGND VPWR VPWR _35996_/D sky130_fd_sc_hd__clkbuf_1
X_34356_ _35701_/CLK _34356_/D VGND VGND VPWR VPWR _34356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21321_ _35688_/Q _32195_/Q _35560_/Q _35496_/Q _21211_/X _21212_/X VGND VGND VPWR
+ VPWR _21321_/X sky130_fd_sc_hd__mux4_1
XFILLER_176_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33307_ _35547_/CLK _33307_/D VGND VGND VPWR VPWR _33307_/Q sky130_fd_sc_hd__dfxtp_1
X_30519_ _30519_/A VGND VGND VPWR VPWR _35499_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34287_ _35822_/CLK _34287_/D VGND VGND VPWR VPWR _34287_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31499_ _27760_/X _35964_/Q _31501_/S VGND VGND VPWR VPWR _31500_/A sky130_fd_sc_hd__mux2_1
XFILLER_198_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33238_ _35804_/CLK _33238_/D VGND VGND VPWR VPWR _33238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21252_ _33062_/Q _32038_/Q _35814_/Q _35750_/Q _20972_/X _20973_/X VGND VGND VPWR
+ VPWR _21252_/X sky130_fd_sc_hd__mux4_1
X_36026_ _36026_/CLK _36026_/D VGND VGND VPWR VPWR _36026_/Q sky130_fd_sc_hd__dfxtp_1
X_24040_ _22974_/X _32562_/Q _24042_/S VGND VGND VPWR VPWR _24041_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20203_ _20203_/A _20203_/B _20203_/C _20203_/D VGND VGND VPWR VPWR _20204_/A sky130_fd_sc_hd__or4_2
XFILLER_172_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33169_ _36047_/CLK _33169_/D VGND VGND VPWR VPWR _33169_/Q sky130_fd_sc_hd__dfxtp_1
X_21183_ _33060_/Q _32036_/Q _35812_/Q _35748_/Q _20972_/X _20973_/X VGND VGND VPWR
+ VPWR _21183_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20134_ _20134_/A VGND VGND VPWR VPWR _20134_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_132_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25991_ _24861_/X _33450_/Q _26009_/S VGND VGND VPWR VPWR _25992_/A sky130_fd_sc_hd__mux2_1
XFILLER_131_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27730_ _27729_/X _34226_/Q _27733_/S VGND VGND VPWR VPWR _27731_/A sky130_fd_sc_hd__mux2_1
X_24942_ input41/X VGND VGND VPWR VPWR _24942_/X sky130_fd_sc_hd__buf_4
X_20065_ _20065_/A VGND VGND VPWR VPWR _20065_/X sky130_fd_sc_hd__clkbuf_4
XTAP_4006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1082 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27661_ input61/X VGND VGND VPWR VPWR _27661_/X sky130_fd_sc_hd__buf_4
XTAP_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24873_ _24873_/A VGND VGND VPWR VPWR _32941_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29400_ _29400_/A VGND VGND VPWR VPWR _34988_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26612_ _24979_/X _33744_/Q _26614_/S VGND VGND VPWR VPWR _26613_/A sky130_fd_sc_hd__mux2_1
XTAP_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23824_ _23058_/X _32397_/Q _23832_/S VGND VGND VPWR VPWR _23825_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27592_ _34175_/Q _27162_/X _27608_/S VGND VGND VPWR VPWR _27593_/A sky130_fd_sc_hd__mux2_1
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29331_ _34966_/Q _29328_/X _29358_/S VGND VGND VPWR VPWR _29332_/A sky130_fd_sc_hd__mux2_1
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26543_ _24877_/X _33711_/Q _26551_/S VGND VGND VPWR VPWR _26544_/A sky130_fd_sc_hd__mux2_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23755_ _22956_/X _32364_/Q _23769_/S VGND VGND VPWR VPWR _23756_/A sky130_fd_sc_hd__mux2_1
XFILLER_242_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20967_ _20960_/X _20966_/X _20644_/X _20646_/X VGND VGND VPWR VPWR _20984_/B sky130_fd_sc_hd__o211a_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22706_ _32656_/Q _32592_/Q _32528_/Q _35984_/Q _22582_/X _21477_/A VGND VGND VPWR
+ VPWR _22706_/X sky130_fd_sc_hd__mux4_1
X_29262_ _34934_/Q _27134_/X _29276_/S VGND VGND VPWR VPWR _29263_/A sky130_fd_sc_hd__mux2_1
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26474_ _33679_/Q _23478_/X _26478_/S VGND VGND VPWR VPWR _26475_/A sky130_fd_sc_hd__mux2_1
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23686_ _23058_/X _32333_/Q _23694_/S VGND VGND VPWR VPWR _23687_/A sky130_fd_sc_hd__mux2_1
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20898_ _35420_/Q _35356_/Q _35292_/Q _35228_/Q _20795_/X _20796_/X VGND VGND VPWR
+ VPWR _20898_/X sky130_fd_sc_hd__mux4_1
XFILLER_109_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28213_ _28213_/A VGND VGND VPWR VPWR _34438_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25425_ _24824_/X _33182_/Q _25427_/S VGND VGND VPWR VPWR _25426_/A sky130_fd_sc_hd__mux2_1
X_22637_ _22637_/A _22637_/B _22637_/C _22637_/D VGND VGND VPWR VPWR _22638_/A sky130_fd_sc_hd__or4_4
XFILLER_201_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29193_ _30337_/A _29797_/A VGND VGND VPWR VPWR _29326_/S sky130_fd_sc_hd__nor2_8
XFILLER_70_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_932 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28144_ _28144_/A VGND VGND VPWR VPWR _34405_/D sky130_fd_sc_hd__clkbuf_1
X_25356_ _33150_/Q _23420_/X _25374_/S VGND VGND VPWR VPWR _25357_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22568_ _22459_/X _22566_/X _22567_/X _22462_/X VGND VGND VPWR VPWR _22568_/X sky130_fd_sc_hd__a22o_1
XFILLER_182_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24307_ _24307_/A VGND VGND VPWR VPWR _32685_/D sky130_fd_sc_hd__clkbuf_1
X_28075_ _34373_/Q _27180_/X _28079_/S VGND VGND VPWR VPWR _28076_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21519_ _33390_/Q _33326_/Q _33262_/Q _33198_/Q _21374_/X _21375_/X VGND VGND VPWR
+ VPWR _21519_/X sky130_fd_sc_hd__mux4_1
XFILLER_186_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25287_ _25287_/A VGND VGND VPWR VPWR _33117_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22499_ _34441_/Q _36169_/Q _34313_/Q _34249_/Q _22182_/X _22183_/X VGND VGND VPWR
+ VPWR _22499_/X sky130_fd_sc_hd__mux4_1
X_27026_ _27026_/A VGND VGND VPWR VPWR _33938_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24238_ _24238_/A VGND VGND VPWR VPWR _32654_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_812 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24169_ _24169_/A VGND VGND VPWR VPWR _32621_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16991_ _16706_/X _16989_/X _16990_/X _16712_/X VGND VGND VPWR VPWR _16991_/X sky130_fd_sc_hd__a22o_1
X_28977_ _34799_/Q _27112_/X _28985_/S VGND VGND VPWR VPWR _28978_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_231_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18730_ _18653_/X _18728_/X _18729_/X _18659_/X VGND VGND VPWR VPWR _18730_/X sky130_fd_sc_hd__a22o_1
X_27928_ _27770_/X _34303_/Q _27944_/S VGND VGND VPWR VPWR _27929_/A sky130_fd_sc_hd__mux2_1
XTAP_5230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18661_ _20212_/A VGND VGND VPWR VPWR _18661_/X sky130_fd_sc_hd__clkbuf_4
X_27859_ _27859_/A VGND VGND VPWR VPWR _34270_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17612_ _17606_/X _17611_/X _17504_/X VGND VGND VPWR VPWR _17620_/C sky130_fd_sc_hd__o21ba_1
XTAP_4573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30870_ _30870_/A VGND VGND VPWR VPWR _35666_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18592_ _20159_/A VGND VGND VPWR VPWR _18592_/X sky130_fd_sc_hd__buf_4
XFILLER_236_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17543_ _34687_/Q _34623_/Q _34559_/Q _34495_/Q _17292_/X _17293_/X VGND VGND VPWR
+ VPWR _17543_/X sky130_fd_sc_hd__mux4_1
XTAP_3872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29529_ _35030_/Q _29328_/X _29547_/S VGND VGND VPWR VPWR _29530_/A sky130_fd_sc_hd__mux2_1
XTAP_3883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32540_ _35998_/CLK _32540_/D VGND VGND VPWR VPWR _32540_/Q sky130_fd_sc_hd__dfxtp_1
X_17474_ _17470_/X _17473_/X _17165_/X VGND VGND VPWR VPWR _17475_/D sky130_fd_sc_hd__o21ba_1
XFILLER_220_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_242_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16425_ _16147_/X _16423_/X _16424_/X _16150_/X VGND VGND VPWR VPWR _16425_/X sky130_fd_sc_hd__a22o_1
X_19213_ _19209_/X _19212_/X _19112_/X VGND VGND VPWR VPWR _19214_/D sky130_fd_sc_hd__o21ba_1
X_32471_ _35929_/CLK _32471_/D VGND VGND VPWR VPWR _32471_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31422_ _27646_/X _35927_/Q _31438_/S VGND VGND VPWR VPWR _31423_/A sky130_fd_sc_hd__mux2_1
X_19144_ _19144_/A _19144_/B _19144_/C _19144_/D VGND VGND VPWR VPWR _19145_/A sky130_fd_sc_hd__or4_2
X_34210_ _36210_/CLK _34210_/D VGND VGND VPWR VPWR _34210_/Q sky130_fd_sc_hd__dfxtp_1
X_16356_ _17906_/A VGND VGND VPWR VPWR _16356_/X sky130_fd_sc_hd__buf_4
X_35190_ _36150_/CLK _35190_/D VGND VGND VPWR VPWR _35190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34141_ _36188_/CLK _34141_/D VGND VGND VPWR VPWR _34141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19075_ _20134_/A VGND VGND VPWR VPWR _19075_/X sky130_fd_sc_hd__clkbuf_4
X_31353_ _31353_/A VGND VGND VPWR VPWR _35894_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16287_ _17833_/A VGND VGND VPWR VPWR _16287_/X sky130_fd_sc_hd__buf_4
XFILLER_195_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30304_ _35398_/Q _29478_/X _30306_/S VGND VGND VPWR VPWR _30305_/A sky130_fd_sc_hd__mux2_1
X_18026_ _35469_/Q _35405_/Q _35341_/Q _35277_/Q _17960_/X _17961_/X VGND VGND VPWR
+ VPWR _18026_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34072_ _35610_/CLK _34072_/D VGND VGND VPWR VPWR _34072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31284_ _31416_/S VGND VGND VPWR VPWR _31303_/S sky130_fd_sc_hd__buf_4
X_33023_ _35903_/CLK _33023_/D VGND VGND VPWR VPWR _33023_/Q sky130_fd_sc_hd__dfxtp_1
X_30235_ _35365_/Q _29376_/X _30243_/S VGND VGND VPWR VPWR _30236_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30166_ _30166_/A VGND VGND VPWR VPWR _35332_/D sky130_fd_sc_hd__clkbuf_1
X_19977_ _19656_/X _19975_/X _19976_/X _19659_/X VGND VGND VPWR VPWR _19977_/X sky130_fd_sc_hd__a22o_1
XFILLER_45_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18928_ _18928_/A VGND VGND VPWR VPWR _32421_/D sky130_fd_sc_hd__clkbuf_1
X_34974_ _35677_/CLK _34974_/D VGND VGND VPWR VPWR _34974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30097_ _30097_/A VGND VGND VPWR VPWR _35299_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_189_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33925_ _34177_/CLK _33925_/D VGND VGND VPWR VPWR _33925_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18859_ _18752_/X _18857_/X _18858_/X _18757_/X VGND VGND VPWR VPWR _18859_/X sky130_fd_sc_hd__a22o_1
XFILLER_227_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_243_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33856_ _33921_/CLK _33856_/D VGND VGND VPWR VPWR _33856_/Q sky130_fd_sc_hd__dfxtp_1
X_21870_ _34168_/Q _34104_/Q _34040_/Q _33976_/Q _21693_/X _21694_/X VGND VGND VPWR
+ VPWR _21870_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20821_ _22586_/A VGND VGND VPWR VPWR _20821_/X sky130_fd_sc_hd__buf_6
X_32807_ _32871_/CLK _32807_/D VGND VGND VPWR VPWR _32807_/Q sky130_fd_sc_hd__dfxtp_1
X_30999_ _30999_/A VGND VGND VPWR VPWR _35727_/D sky130_fd_sc_hd__clkbuf_1
X_33787_ _36092_/CLK _33787_/D VGND VGND VPWR VPWR _33787_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23540_ _23540_/A VGND VGND VPWR VPWR _32264_/D sky130_fd_sc_hd__clkbuf_1
X_35526_ _35721_/CLK _35526_/D VGND VGND VPWR VPWR _35526_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20752_ _20746_/X _20751_/X _20615_/X VGND VGND VPWR VPWR _20776_/A sky130_fd_sc_hd__o21ba_1
X_32738_ _35871_/CLK _32738_/D VGND VGND VPWR VPWR _32738_/Q sky130_fd_sc_hd__dfxtp_1
X_20683_ _22316_/A VGND VGND VPWR VPWR _20683_/X sky130_fd_sc_hd__clkbuf_8
X_23471_ _23471_/A VGND VGND VPWR VPWR _32235_/D sky130_fd_sc_hd__clkbuf_1
X_35457_ _35458_/CLK _35457_/D VGND VGND VPWR VPWR _35457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32669_ _32797_/CLK _32669_/D VGND VGND VPWR VPWR _32669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25210_ _25210_/A VGND VGND VPWR VPWR _33081_/D sky130_fd_sc_hd__clkbuf_1
X_22422_ _35207_/Q _35143_/Q _35079_/Q _32263_/Q _22316_/X _22317_/X VGND VGND VPWR
+ VPWR _22422_/X sky130_fd_sc_hd__mux4_1
X_34408_ _34914_/CLK _34408_/D VGND VGND VPWR VPWR _34408_/Q sky130_fd_sc_hd__dfxtp_1
X_26190_ _26190_/A VGND VGND VPWR VPWR _33544_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35388_ _35708_/CLK _35388_/D VGND VGND VPWR VPWR _35388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25141_ _25141_/A VGND VGND VPWR VPWR _33048_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22353_ _34949_/Q _34885_/Q _34821_/Q _34757_/Q _22113_/X _22114_/X VGND VGND VPWR
+ VPWR _22353_/X sky130_fd_sc_hd__mux4_1
X_34339_ _35618_/CLK _34339_/D VGND VGND VPWR VPWR _34339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21304_ _21100_/X _21302_/X _21303_/X _21103_/X VGND VGND VPWR VPWR _21304_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_6_6__f_CLK clkbuf_5_3_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_6__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_22284_ _22111_/X _22282_/X _22283_/X _22116_/X VGND VGND VPWR VPWR _22284_/X sky130_fd_sc_hd__a22o_1
X_25072_ _24908_/X _33017_/Q _25080_/S VGND VGND VPWR VPWR _25073_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28900_ _28900_/A VGND VGND VPWR VPWR _34762_/D sky130_fd_sc_hd__clkbuf_1
X_21235_ _21231_/X _21234_/X _21026_/X VGND VGND VPWR VPWR _21265_/A sky130_fd_sc_hd__o21ba_1
XFILLER_2_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36009_ _36011_/CLK _36009_/D VGND VGND VPWR VPWR _36009_/Q sky130_fd_sc_hd__dfxtp_1
X_24023_ _24113_/S VGND VGND VPWR VPWR _24042_/S sky130_fd_sc_hd__buf_4
X_29880_ _35197_/Q _29450_/X _29880_/S VGND VGND VPWR VPWR _29881_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21166_ _33380_/Q _33316_/Q _33252_/Q _33188_/Q _21021_/X _21022_/X VGND VGND VPWR
+ VPWR _21166_/X sky130_fd_sc_hd__mux4_1
X_28831_ _28921_/S VGND VGND VPWR VPWR _28850_/S sky130_fd_sc_hd__buf_4
XFILLER_49_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20117_ _35463_/Q _35399_/Q _35335_/Q _35271_/Q _19907_/X _19908_/X VGND VGND VPWR
+ VPWR _20117_/X sky130_fd_sc_hd__mux4_1
X_28762_ _34698_/Q _27196_/X _28776_/S VGND VGND VPWR VPWR _28763_/A sky130_fd_sc_hd__mux2_1
XFILLER_131_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21097_ _34146_/Q _34082_/Q _34018_/Q _33954_/Q _20987_/X _20988_/X VGND VGND VPWR
+ VPWR _21097_/X sky130_fd_sc_hd__mux4_1
XFILLER_24_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25974_ _24837_/X _33442_/Q _25988_/S VGND VGND VPWR VPWR _25975_/A sky130_fd_sc_hd__mux2_1
X_27713_ _27713_/A VGND VGND VPWR VPWR _34220_/D sky130_fd_sc_hd__clkbuf_1
X_20048_ _20044_/X _20047_/X _19804_/X VGND VGND VPWR VPWR _20056_/C sky130_fd_sc_hd__o21ba_1
X_24925_ _24923_/X _32958_/Q _24952_/S VGND VGND VPWR VPWR _24926_/A sky130_fd_sc_hd__mux2_1
X_28693_ _28693_/A VGND VGND VPWR VPWR _34665_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_246_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27644_ _27639_/X _34198_/Q _27671_/S VGND VGND VPWR VPWR _27645_/A sky130_fd_sc_hd__mux2_1
XFILLER_206_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24856_ _24855_/X _32936_/Q _24859_/S VGND VGND VPWR VPWR _24857_/A sky130_fd_sc_hd__mux2_1
XTAP_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1071 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23807_ _23033_/X _32389_/Q _23811_/S VGND VGND VPWR VPWR _23808_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27575_ _34167_/Q _27137_/X _27587_/S VGND VGND VPWR VPWR _27576_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24787_ _24787_/A VGND VGND VPWR VPWR _32913_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21999_ _34427_/Q _36155_/Q _34299_/Q _34235_/Q _21829_/X _21830_/X VGND VGND VPWR
+ VPWR _21999_/X sky130_fd_sc_hd__mux4_1
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29314_ _34959_/Q _27211_/X _29318_/S VGND VGND VPWR VPWR _29315_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26526_ _24852_/X _33703_/Q _26530_/S VGND VGND VPWR VPWR _26527_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23738_ _22931_/X _32356_/Q _23748_/S VGND VGND VPWR VPWR _23739_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_241_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29245_ _34926_/Q _27109_/X _29255_/S VGND VGND VPWR VPWR _29246_/A sky130_fd_sc_hd__mux2_1
X_26457_ _33671_/Q _23450_/X _26457_/S VGND VGND VPWR VPWR _26458_/A sky130_fd_sc_hd__mux2_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23669_ _23033_/X _32325_/Q _23673_/S VGND VGND VPWR VPWR _23670_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16210_ _33626_/Q _33562_/Q _33498_/Q _33434_/Q _16141_/X _16142_/X VGND VGND VPWR
+ VPWR _16210_/X sky130_fd_sc_hd__mux4_1
XFILLER_224_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25408_ _25540_/S VGND VGND VPWR VPWR _25427_/S sky130_fd_sc_hd__buf_4
XFILLER_14_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29176_ _29176_/A VGND VGND VPWR VPWR _34893_/D sky130_fd_sc_hd__clkbuf_1
X_17190_ _34677_/Q _34613_/Q _34549_/Q _34485_/Q _16939_/X _16940_/X VGND VGND VPWR
+ VPWR _17190_/X sky130_fd_sc_hd__mux4_1
XFILLER_167_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26388_ _33638_/Q _23280_/X _26394_/S VGND VGND VPWR VPWR _26389_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_1356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28127_ _28127_/A VGND VGND VPWR VPWR _34397_/D sky130_fd_sc_hd__clkbuf_1
X_16141_ _17906_/A VGND VGND VPWR VPWR _16141_/X sky130_fd_sc_hd__buf_6
X_25339_ _33142_/Q _23396_/X _25353_/S VGND VGND VPWR VPWR _25340_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16072_ _17869_/A VGND VGND VPWR VPWR _16072_/X sky130_fd_sc_hd__buf_4
XFILLER_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28058_ _34365_/Q _27155_/X _28058_/S VGND VGND VPWR VPWR _28059_/A sky130_fd_sc_hd__mux2_1
X_27009_ _33930_/Q _23463_/X _27023_/S VGND VGND VPWR VPWR _27010_/A sky130_fd_sc_hd__mux2_1
X_19900_ _32129_/Q _32321_/Q _32385_/Q _35905_/Q _19580_/X _19721_/X VGND VGND VPWR
+ VPWR _19900_/X sky130_fd_sc_hd__mux4_1
XFILLER_135_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30020_ _35263_/Q _29457_/X _30036_/S VGND VGND VPWR VPWR _30021_/A sky130_fd_sc_hd__mux2_1
X_19831_ _19712_/X _19829_/X _19830_/X _19718_/X VGND VGND VPWR VPWR _19831_/X sky130_fd_sc_hd__a22o_1
XFILLER_190_1135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19762_ _35645_/Q _35005_/Q _34365_/Q _33725_/Q _19444_/X _19445_/X VGND VGND VPWR
+ VPWR _19762_/X sky130_fd_sc_hd__mux4_1
XFILLER_231_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16974_ _35183_/Q _35119_/Q _35055_/Q _32176_/Q _16657_/X _16658_/X VGND VGND VPWR
+ VPWR _16974_/X sky130_fd_sc_hd__mux4_1
X_18713_ _34911_/Q _34847_/Q _34783_/Q _34719_/Q _18396_/X _18398_/X VGND VGND VPWR
+ VPWR _18713_/X sky130_fd_sc_hd__mux4_1
XFILLER_77_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31971_ _34085_/CLK _31971_/D VGND VGND VPWR VPWR _31971_/Q sky130_fd_sc_hd__dfxtp_1
X_19693_ _33083_/Q _32059_/Q _35835_/Q _35771_/Q _19378_/X _19379_/X VGND VGND VPWR
+ VPWR _19693_/X sky130_fd_sc_hd__mux4_1
XTAP_5082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 DW[16] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__buf_6
XFILLER_64_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_292_CLK clkbuf_6_56__f_CLK/X VGND VGND VPWR VPWR _35902_/CLK sky130_fd_sc_hd__clkbuf_16
X_33710_ _35630_/CLK _33710_/D VGND VGND VPWR VPWR _33710_/Q sky130_fd_sc_hd__dfxtp_1
X_18644_ _18644_/A _18644_/B _18644_/C _18644_/D VGND VGND VPWR VPWR _18645_/A sky130_fd_sc_hd__or4_1
X_30922_ _30922_/A VGND VGND VPWR VPWR _35690_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_225_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34690_ _34690_/CLK _34690_/D VGND VGND VPWR VPWR _34690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_840 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30853_ _35658_/Q input48/X _30867_/S VGND VGND VPWR VPWR _30854_/A sky130_fd_sc_hd__mux2_1
X_33641_ _34153_/CLK _33641_/D VGND VGND VPWR VPWR _33641_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_1097 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18575_ _18575_/A VGND VGND VPWR VPWR _32411_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_75_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17526_ _33919_/Q _33855_/Q _33791_/Q _36095_/Q _17377_/X _17378_/X VGND VGND VPWR
+ VPWR _17526_/X sky130_fd_sc_hd__mux4_1
X_33572_ _34151_/CLK _33572_/D VGND VGND VPWR VPWR _33572_/Q sky130_fd_sc_hd__dfxtp_1
X_30784_ _30784_/A VGND VGND VPWR VPWR _35625_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35311_ _35438_/CLK _35311_/D VGND VGND VPWR VPWR _35311_/Q sky130_fd_sc_hd__dfxtp_1
X_32523_ _35980_/CLK _32523_/D VGND VGND VPWR VPWR _32523_/Q sky130_fd_sc_hd__dfxtp_1
X_17457_ _32125_/Q _32317_/Q _32381_/Q _35901_/Q _17280_/X _17421_/X VGND VGND VPWR
+ VPWR _17457_/X sky130_fd_sc_hd__mux4_1
XFILLER_75_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16408_ _16404_/X _16407_/X _16075_/X VGND VGND VPWR VPWR _16416_/C sky130_fd_sc_hd__o21ba_1
XFILLER_242_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35242_ _35434_/CLK _35242_/D VGND VGND VPWR VPWR _35242_/Q sky130_fd_sc_hd__dfxtp_1
X_32454_ _36085_/CLK _32454_/D VGND VGND VPWR VPWR _32454_/Q sky130_fd_sc_hd__dfxtp_1
X_17388_ _17384_/X _17387_/X _17140_/X _17141_/X VGND VGND VPWR VPWR _17403_/B sky130_fd_sc_hd__o211a_1
XFILLER_146_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16339_ _16078_/X _16337_/X _16338_/X _16088_/X VGND VGND VPWR VPWR _16339_/X sky130_fd_sc_hd__a22o_1
X_31405_ _31405_/A VGND VGND VPWR VPWR _35919_/D sky130_fd_sc_hd__clkbuf_1
X_19127_ _32875_/Q _32811_/Q _32747_/Q _32683_/Q _18940_/X _18941_/X VGND VGND VPWR
+ VPWR _19127_/X sky130_fd_sc_hd__mux4_1
X_32385_ _35902_/CLK _32385_/D VGND VGND VPWR VPWR _32385_/Q sky130_fd_sc_hd__dfxtp_1
X_35173_ _35490_/CLK _35173_/D VGND VGND VPWR VPWR _35173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34124_ _34188_/CLK _34124_/D VGND VGND VPWR VPWR _34124_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19058_ _35433_/Q _35369_/Q _35305_/Q _35241_/Q _18848_/X _18849_/X VGND VGND VPWR
+ VPWR _19058_/X sky130_fd_sc_hd__mux4_1
X_31336_ _31336_/A VGND VGND VPWR VPWR _35886_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18009_ _33677_/Q _33613_/Q _33549_/Q _33485_/Q _17906_/X _17907_/X VGND VGND VPWR
+ VPWR _18009_/X sky130_fd_sc_hd__mux4_1
XFILLER_160_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34055_ _34945_/CLK _34055_/D VGND VGND VPWR VPWR _34055_/Q sky130_fd_sc_hd__dfxtp_1
X_31267_ _27816_/X _35854_/Q _31273_/S VGND VGND VPWR VPWR _31268_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_940 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21020_ _20740_/X _21018_/X _21019_/X _20745_/X VGND VGND VPWR VPWR _21020_/X sky130_fd_sc_hd__a22o_1
X_30218_ _35357_/Q _29351_/X _30222_/S VGND VGND VPWR VPWR _30219_/A sky130_fd_sc_hd__mux2_1
X_33006_ _36015_/CLK _33006_/D VGND VGND VPWR VPWR _33006_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31198_ _27714_/X _35821_/Q _31210_/S VGND VGND VPWR VPWR _31199_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_1238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30149_ _30149_/A VGND VGND VPWR VPWR _35324_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34957_ _34957_/CLK _34957_/D VGND VGND VPWR VPWR _34957_/Q sky130_fd_sc_hd__dfxtp_1
X_22971_ input20/X VGND VGND VPWR VPWR _22971_/X sky130_fd_sc_hd__buf_2
XFILLER_68_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_283_CLK clkbuf_6_58__f_CLK/X VGND VGND VPWR VPWR _35713_/CLK sky130_fd_sc_hd__clkbuf_16
X_24710_ _24710_/A VGND VGND VPWR VPWR _32876_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33908_ _36085_/CLK _33908_/D VGND VGND VPWR VPWR _33908_/Q sky130_fd_sc_hd__dfxtp_1
X_21922_ _35449_/Q _35385_/Q _35321_/Q _35257_/Q _21854_/X _21855_/X VGND VGND VPWR
+ VPWR _21922_/X sky130_fd_sc_hd__mux4_1
XFILLER_56_957 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25690_ _25690_/A VGND VGND VPWR VPWR _33307_/D sky130_fd_sc_hd__clkbuf_1
X_34888_ _34954_/CLK _34888_/D VGND VGND VPWR VPWR _34888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24641_ _23055_/X _32844_/Q _24651_/S VGND VGND VPWR VPWR _24642_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33839_ _33902_/CLK _33839_/D VGND VGND VPWR VPWR _33839_/Q sky130_fd_sc_hd__dfxtp_1
X_21853_ _21598_/X _21851_/X _21852_/X _21601_/X VGND VGND VPWR VPWR _21853_/X sky130_fd_sc_hd__a22o_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27360_ _27360_/A VGND VGND VPWR VPWR _34065_/D sky130_fd_sc_hd__clkbuf_1
X_20804_ _34393_/Q _36121_/Q _34265_/Q _34201_/Q _20770_/X _20771_/X VGND VGND VPWR
+ VPWR _20804_/X sky130_fd_sc_hd__mux4_1
XFILLER_70_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24572_ _22953_/X _32811_/Q _24588_/S VGND VGND VPWR VPWR _24573_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_1304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21784_ _35637_/Q _34997_/Q _34357_/Q _33717_/Q _21744_/X _21745_/X VGND VGND VPWR
+ VPWR _21784_/X sky130_fd_sc_hd__mux4_1
XFILLER_223_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_247_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26311_ _24936_/X _33602_/Q _26321_/S VGND VGND VPWR VPWR _26312_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23523_ _23523_/A VGND VGND VPWR VPWR _32256_/D sky130_fd_sc_hd__clkbuf_1
X_35509_ _35701_/CLK _35509_/D VGND VGND VPWR VPWR _35509_/Q sky130_fd_sc_hd__dfxtp_1
X_20735_ _34903_/Q _34839_/Q _34775_/Q _34711_/Q _20696_/X _20698_/X VGND VGND VPWR
+ VPWR _20735_/X sky130_fd_sc_hd__mux4_1
XFILLER_195_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27291_ _27291_/A VGND VGND VPWR VPWR _34032_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29030_ _34824_/Q _27189_/X _29048_/S VGND VGND VPWR VPWR _29031_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26242_ _24834_/X _33569_/Q _26258_/S VGND VGND VPWR VPWR _26243_/A sky130_fd_sc_hd__mux2_1
X_23454_ _23499_/S VGND VGND VPWR VPWR _23485_/S sky130_fd_sc_hd__buf_4
X_20666_ _22582_/A VGND VGND VPWR VPWR _22535_/A sky130_fd_sc_hd__buf_12
XFILLER_17_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22405_ _22159_/X _22403_/X _22404_/X _22162_/X VGND VGND VPWR VPWR _22405_/X sky130_fd_sc_hd__a22o_1
X_26173_ _26173_/A VGND VGND VPWR VPWR _33536_/D sky130_fd_sc_hd__clkbuf_1
X_20597_ _20581_/X _20588_/X _20591_/X _20596_/X VGND VGND VPWR VPWR _20597_/X sky130_fd_sc_hd__a22o_1
XFILLER_137_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23385_ _32207_/Q _23384_/X _23385_/S VGND VGND VPWR VPWR _23386_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25124_ _24985_/X _33042_/Q _25130_/S VGND VGND VPWR VPWR _25125_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22336_ _33157_/Q _36037_/Q _33029_/Q _32965_/Q _22015_/X _22016_/X VGND VGND VPWR
+ VPWR _22336_/X sky130_fd_sc_hd__mux4_1
XFILLER_118_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29932_ _30877_/A _31688_/A VGND VGND VPWR VPWR _30065_/S sky130_fd_sc_hd__nor2_8
XFILLER_152_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25055_ _24883_/X _33009_/Q _25059_/S VGND VGND VPWR VPWR _25056_/A sky130_fd_sc_hd__mux2_1
X_22267_ _32899_/Q _32835_/Q _32771_/Q _32707_/Q _21946_/X _21947_/X VGND VGND VPWR
+ VPWR _22267_/X sky130_fd_sc_hd__mux4_1
XFILLER_2_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24006_ _24006_/A VGND VGND VPWR VPWR _32545_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21218_ _20897_/X _21216_/X _21217_/X _20900_/X VGND VGND VPWR VPWR _21218_/X sky130_fd_sc_hd__a22o_1
X_22198_ _33153_/Q _36033_/Q _33025_/Q _32961_/Q _22015_/X _22016_/X VGND VGND VPWR
+ VPWR _22198_/X sky130_fd_sc_hd__mux4_1
XFILLER_132_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29863_ _29863_/A VGND VGND VPWR VPWR _35188_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_819 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28814_ _28814_/A VGND VGND VPWR VPWR _34721_/D sky130_fd_sc_hd__clkbuf_1
X_21149_ _22561_/A VGND VGND VPWR VPWR _21149_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_232_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29794_ _29794_/A VGND VGND VPWR VPWR _35156_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28745_ _34690_/Q _27171_/X _28755_/S VGND VGND VPWR VPWR _28746_/A sky130_fd_sc_hd__mux2_1
X_25957_ _24812_/X _33434_/Q _25967_/S VGND VGND VPWR VPWR _25958_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_274_CLK clkbuf_6_59__f_CLK/X VGND VGND VPWR VPWR _35777_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_207_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24908_ input29/X VGND VGND VPWR VPWR _24908_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_58_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_246_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16690_ _34663_/Q _34599_/Q _34535_/Q _34471_/Q _16586_/X _16587_/X VGND VGND VPWR
+ VPWR _16690_/X sky130_fd_sc_hd__mux4_1
X_28676_ _34657_/Q _27069_/X _28692_/S VGND VGND VPWR VPWR _28677_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25888_ _25888_/A VGND VGND VPWR VPWR _33401_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_749 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27627_ _34192_/Q _27214_/X _27629_/S VGND VGND VPWR VPWR _27628_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_5_30_0_CLK clkbuf_2_3_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_30_0_CLK/X sky130_fd_sc_hd__clkbuf_8
X_24839_ _24839_/A VGND VGND VPWR VPWR _32930_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18360_ _20164_/A VGND VGND VPWR VPWR _18360_/X sky130_fd_sc_hd__buf_4
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27558_ _34159_/Q _27112_/X _27566_/S VGND VGND VPWR VPWR _27559_/A sky130_fd_sc_hd__mux2_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ _33145_/Q _36025_/Q _33017_/Q _32953_/Q _17062_/X _17063_/X VGND VGND VPWR
+ VPWR _17311_/X sky130_fd_sc_hd__mux4_1
X_26509_ _24827_/X _33695_/Q _26509_/S VGND VGND VPWR VPWR _26510_/A sky130_fd_sc_hd__mux2_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18291_ _20210_/A VGND VGND VPWR VPWR _18291_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27489_ _27489_/A VGND VGND VPWR VPWR _34126_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17242_ _17206_/X _17240_/X _17241_/X _17209_/X VGND VGND VPWR VPWR _17242_/X sky130_fd_sc_hd__a22o_1
XFILLER_147_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29228_ _34918_/Q _27084_/X _29234_/S VGND VGND VPWR VPWR _29229_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29159_ _29159_/A VGND VGND VPWR VPWR _34885_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17173_ _33909_/Q _33845_/Q _33781_/Q _36085_/Q _17024_/X _17025_/X VGND VGND VPWR
+ VPWR _17173_/X sky130_fd_sc_hd__mux4_1
XFILLER_200_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16124_ _35671_/Q _32177_/Q _35543_/Q _35479_/Q _16049_/X _16050_/X VGND VGND VPWR
+ VPWR _16124_/X sky130_fd_sc_hd__mux4_1
X_32170_ _35434_/CLK _32170_/D VGND VGND VPWR VPWR _32170_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31121_ _35785_/Q input47/X _31137_/S VGND VGND VPWR VPWR _31122_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16055_ _17999_/A VGND VGND VPWR VPWR _16055_/X sky130_fd_sc_hd__buf_4
XFILLER_143_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31052_ _31052_/A VGND VGND VPWR VPWR _35752_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30003_ _35255_/Q _29432_/X _30015_/S VGND VGND VPWR VPWR _30004_/A sky130_fd_sc_hd__mux2_1
X_19814_ _20167_/A VGND VGND VPWR VPWR _19814_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_233_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35860_ _35860_/CLK _35860_/D VGND VGND VPWR VPWR _35860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_1096 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34811_ _34941_/CLK _34811_/D VGND VGND VPWR VPWR _34811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19745_ _33661_/Q _33597_/Q _33533_/Q _33469_/Q _19500_/X _19501_/X VGND VGND VPWR
+ VPWR _19745_/X sky130_fd_sc_hd__mux4_1
XFILLER_81_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35791_ _35853_/CLK _35791_/D VGND VGND VPWR VPWR _35791_/Q sky130_fd_sc_hd__dfxtp_1
X_16957_ _32623_/Q _32559_/Q _32495_/Q _35951_/Q _16923_/X _16707_/X VGND VGND VPWR
+ VPWR _16957_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_265_CLK clkbuf_6_62__f_CLK/X VGND VGND VPWR VPWR _36103_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_77_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34742_ _36151_/CLK _34742_/D VGND VGND VPWR VPWR _34742_/Q sky130_fd_sc_hd__dfxtp_1
X_31954_ _23495_/X _36180_/Q _31956_/S VGND VGND VPWR VPWR _31955_/A sky130_fd_sc_hd__mux2_1
X_19676_ _33403_/Q _33339_/Q _33275_/Q _33211_/Q _19427_/X _19428_/X VGND VGND VPWR
+ VPWR _19676_/X sky130_fd_sc_hd__mux4_1
X_16888_ _33901_/Q _33837_/Q _33773_/Q _36077_/Q _16671_/X _16672_/X VGND VGND VPWR
+ VPWR _16888_/X sky130_fd_sc_hd__mux4_1
XFILLER_53_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18627_ _32861_/Q _32797_/Q _32733_/Q _32669_/Q _18587_/X _18588_/X VGND VGND VPWR
+ VPWR _18627_/X sky130_fd_sc_hd__mux4_1
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30905_ _30905_/A VGND VGND VPWR VPWR _35682_/D sky130_fd_sc_hd__clkbuf_1
X_34673_ _35633_/CLK _34673_/D VGND VGND VPWR VPWR _34673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31885_ _23384_/X _36147_/Q _31885_/S VGND VGND VPWR VPWR _31886_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33624_ _34331_/CLK _33624_/D VGND VGND VPWR VPWR _33624_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_212_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30836_ _35650_/Q input39/X _30846_/S VGND VGND VPWR VPWR _30837_/A sky130_fd_sc_hd__mux2_1
X_18558_ _20099_/A VGND VGND VPWR VPWR _18558_/X sky130_fd_sc_hd__buf_6
XFILLER_127_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17509_ _17862_/A VGND VGND VPWR VPWR _17509_/X sky130_fd_sc_hd__clkbuf_4
X_33555_ _33875_/CLK _33555_/D VGND VGND VPWR VPWR _33555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18489_ _32857_/Q _32793_/Q _32729_/Q _32665_/Q _18337_/X _18339_/X VGND VGND VPWR
+ VPWR _18489_/X sky130_fd_sc_hd__mux4_1
XFILLER_162_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30767_ _35617_/Q input3/X _30783_/S VGND VGND VPWR VPWR _30768_/A sky130_fd_sc_hd__mux2_1
X_20520_ _34196_/Q _34132_/Q _34068_/Q _34004_/Q _18349_/X _18350_/X VGND VGND VPWR
+ VPWR _20520_/X sky130_fd_sc_hd__mux4_1
XFILLER_123_1018 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32506_ _35962_/CLK _32506_/D VGND VGND VPWR VPWR _32506_/Q sky130_fd_sc_hd__dfxtp_1
X_33486_ _34064_/CLK _33486_/D VGND VGND VPWR VPWR _33486_/Q sky130_fd_sc_hd__dfxtp_1
X_30698_ _30698_/A VGND VGND VPWR VPWR _35584_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_1198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20451_ _35217_/Q _35153_/Q _35089_/Q _32273_/Q _18392_/X _18394_/X VGND VGND VPWR
+ VPWR _20451_/X sky130_fd_sc_hd__mux4_1
XFILLER_203_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35225_ _35674_/CLK _35225_/D VGND VGND VPWR VPWR _35225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_19__f_CLK clkbuf_5_9_0_CLK/X VGND VGND VPWR VPWR clkbuf_leaf_81_CLK/A sky130_fd_sc_hd__clkbuf_16
XFILLER_119_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32437_ _33897_/CLK _32437_/D VGND VGND VPWR VPWR _32437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_1305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35156_ _35221_/CLK _35156_/D VGND VGND VPWR VPWR _35156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20382_ _20378_/X _20381_/X _20146_/X _20147_/X VGND VGND VPWR VPWR _20397_/B sky130_fd_sc_hd__o211a_1
X_23170_ _23170_/A VGND VGND VPWR VPWR _32123_/D sky130_fd_sc_hd__clkbuf_1
X_32368_ _35952_/CLK _32368_/D VGND VGND VPWR VPWR _32368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22121_ _22121_/A VGND VGND VPWR VPWR _36222_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34107_ _35449_/CLK _34107_/D VGND VGND VPWR VPWR _34107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31319_ _31319_/A VGND VGND VPWR VPWR _35878_/D sky130_fd_sc_hd__clkbuf_1
X_35087_ _35217_/CLK _35087_/D VGND VGND VPWR VPWR _35087_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput120 _31995_/Q VGND VGND VPWR VPWR D1[37] sky130_fd_sc_hd__buf_2
X_32299_ _32875_/CLK _32299_/D VGND VGND VPWR VPWR _32299_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput131 _32005_/Q VGND VGND VPWR VPWR D1[47] sky130_fd_sc_hd__buf_2
XFILLER_115_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput142 _32015_/Q VGND VGND VPWR VPWR D1[57] sky130_fd_sc_hd__buf_2
XTAP_6508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22052_ _21806_/X _22050_/X _22051_/X _21809_/X VGND VGND VPWR VPWR _22052_/X sky130_fd_sc_hd__a22o_1
XTAP_6519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34038_ _34166_/CLK _34038_/D VGND VGND VPWR VPWR _34038_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput153 _31967_/Q VGND VGND VPWR VPWR D1[9] sky130_fd_sc_hd__buf_2
XFILLER_86_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput164 _36201_/Q VGND VGND VPWR VPWR D2[19] sky130_fd_sc_hd__buf_2
Xoutput175 _36211_/Q VGND VGND VPWR VPWR D2[29] sky130_fd_sc_hd__buf_2
XFILLER_99_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput186 _36221_/Q VGND VGND VPWR VPWR D2[39] sky130_fd_sc_hd__buf_2
XFILLER_142_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput197 _36231_/Q VGND VGND VPWR VPWR D2[49] sky130_fd_sc_hd__buf_2
XTAP_5807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21003_ _35615_/Q _34975_/Q _34335_/Q _33695_/Q _20653_/X _20655_/X VGND VGND VPWR
+ VPWR _21003_/X sky130_fd_sc_hd__mux4_1
XTAP_5818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26860_ _26860_/A VGND VGND VPWR VPWR _33859_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25811_ _25811_/A VGND VGND VPWR VPWR _33365_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_229_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26791_ _26791_/A VGND VGND VPWR VPWR _33826_/D sky130_fd_sc_hd__clkbuf_1
X_35989_ _35989_/CLK _35989_/D VGND VGND VPWR VPWR _35989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_256_CLK clkbuf_6_63__f_CLK/X VGND VGND VPWR VPWR _33984_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_101_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28530_ _28530_/A VGND VGND VPWR VPWR _34588_/D sky130_fd_sc_hd__clkbuf_1
X_25742_ _24892_/X _33332_/Q _25760_/S VGND VGND VPWR VPWR _25743_/A sky130_fd_sc_hd__mux2_1
XFILLER_244_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22954_ _22953_/X _32043_/Q _22978_/S VGND VGND VPWR VPWR _22955_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21905_ _21799_/X _21903_/X _21904_/X _21804_/X VGND VGND VPWR VPWR _21905_/X sky130_fd_sc_hd__a22o_1
X_28461_ _27760_/X _34556_/Q _28463_/S VGND VGND VPWR VPWR _28462_/A sky130_fd_sc_hd__mux2_1
X_25673_ _24991_/X _33300_/Q _25675_/S VGND VGND VPWR VPWR _25674_/A sky130_fd_sc_hd__mux2_1
X_22885_ _22885_/A VGND VGND VPWR VPWR _30202_/A sky130_fd_sc_hd__buf_4
XFILLER_243_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27412_ _27502_/S VGND VGND VPWR VPWR _27431_/S sky130_fd_sc_hd__buf_4
X_24624_ _23030_/X _32836_/Q _24630_/S VGND VGND VPWR VPWR _24625_/A sky130_fd_sc_hd__mux2_1
X_28392_ _27658_/X _34523_/Q _28400_/S VGND VGND VPWR VPWR _28393_/A sky130_fd_sc_hd__mux2_1
X_21836_ _21836_/A VGND VGND VPWR VPWR _36214_/D sky130_fd_sc_hd__buf_6
XFILLER_145_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27343_ _34057_/Q _27193_/X _27359_/S VGND VGND VPWR VPWR _27344_/A sky130_fd_sc_hd__mux2_1
X_24555_ _22928_/X _32803_/Q _24567_/S VGND VGND VPWR VPWR _24556_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21767_ _21767_/A _21767_/B _21767_/C _21767_/D VGND VGND VPWR VPWR _21768_/A sky130_fd_sc_hd__or4_1
XFILLER_145_1254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23506_ _23506_/A VGND VGND VPWR VPWR _32248_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20718_ _33111_/Q _35991_/Q _32983_/Q _32919_/Q _20624_/X _20625_/X VGND VGND VPWR
+ VPWR _20718_/X sky130_fd_sc_hd__mux4_1
XFILLER_8_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27274_ _27274_/A VGND VGND VPWR VPWR _34024_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24486_ _24486_/A VGND VGND VPWR VPWR _32770_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21698_ _33907_/Q _33843_/Q _33779_/Q _36083_/Q _21624_/X _21625_/X VGND VGND VPWR
+ VPWR _21698_/X sky130_fd_sc_hd__mux4_1
X_29013_ _34816_/Q _27165_/X _29027_/S VGND VGND VPWR VPWR _29014_/A sky130_fd_sc_hd__mux2_1
XFILLER_200_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26225_ _24809_/X _33561_/Q _26237_/S VGND VGND VPWR VPWR _26226_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23437_ _23437_/A VGND VGND VPWR VPWR _32224_/D sky130_fd_sc_hd__clkbuf_1
X_20649_ _22399_/A VGND VGND VPWR VPWR _20649_/X sky130_fd_sc_hd__buf_6
XFILLER_165_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26156_ _26156_/A VGND VGND VPWR VPWR _33528_/D sky130_fd_sc_hd__clkbuf_1
X_23368_ _23368_/A VGND VGND VPWR VPWR _32199_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25107_ _25107_/A VGND VGND VPWR VPWR _33033_/D sky130_fd_sc_hd__clkbuf_1
X_22319_ _22106_/X _22315_/X _22318_/X _22109_/X VGND VGND VPWR VPWR _22319_/X sky130_fd_sc_hd__a22o_1
X_26087_ _26087_/A VGND VGND VPWR VPWR _33495_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23299_ input15/X VGND VGND VPWR VPWR _23299_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_65_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29915_ _29915_/A VGND VGND VPWR VPWR _35213_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25038_ _24858_/X _33001_/Q _25038_/S VGND VGND VPWR VPWR _25039_/A sky130_fd_sc_hd__mux2_1
XFILLER_191_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_495_CLK clkbuf_6_3__f_CLK/X VGND VGND VPWR VPWR _35620_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_61_1108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17860_ _34696_/Q _34632_/Q _34568_/Q _34504_/Q _17645_/X _17646_/X VGND VGND VPWR
+ VPWR _17860_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29846_ _29846_/A VGND VGND VPWR VPWR _35180_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_1296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16811_ _16805_/X _16806_/X _16809_/X _16810_/X VGND VGND VPWR VPWR _16811_/X sky130_fd_sc_hd__a22o_1
XFILLER_117_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29777_ _35148_/Q _29497_/X _29787_/S VGND VGND VPWR VPWR _29778_/A sky130_fd_sc_hd__mux2_1
X_17791_ _17506_/X _17789_/X _17790_/X _17509_/X VGND VGND VPWR VPWR _17791_/X sky130_fd_sc_hd__a22o_1
XFILLER_66_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26989_ _26989_/A VGND VGND VPWR VPWR _33920_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_247_CLK clkbuf_6_61__f_CLK/X VGND VGND VPWR VPWR _33420_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_232_1293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19530_ _20236_/A VGND VGND VPWR VPWR _19530_/X sky130_fd_sc_hd__buf_6
XFILLER_235_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16742_ _34153_/Q _34089_/Q _34025_/Q _33961_/Q _16740_/X _16741_/X VGND VGND VPWR
+ VPWR _16742_/X sky130_fd_sc_hd__mux4_1
X_28728_ _34682_/Q _27146_/X _28734_/S VGND VGND VPWR VPWR _28729_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16673_ _33895_/Q _33831_/Q _33767_/Q _36071_/Q _16671_/X _16672_/X VGND VGND VPWR
+ VPWR _16673_/X sky130_fd_sc_hd__mux4_1
X_19461_ _19461_/A VGND VGND VPWR VPWR _19461_/X sky130_fd_sc_hd__buf_4
XFILLER_62_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28659_ _34649_/Q _27044_/X _28671_/S VGND VGND VPWR VPWR _28660_/A sky130_fd_sc_hd__mux2_1
XFILLER_189_1192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1075 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18412_ _20150_/A VGND VGND VPWR VPWR _18412_/X sky130_fd_sc_hd__buf_6
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31670_ _27813_/X _36045_/Q _31678_/S VGND VGND VPWR VPWR _31671_/A sky130_fd_sc_hd__mux2_1
X_19392_ _33651_/Q _33587_/Q _33523_/Q _33459_/Q _19147_/X _19148_/X VGND VGND VPWR
+ VPWR _19392_/X sky130_fd_sc_hd__mux4_1
XFILLER_34_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30621_ _35548_/Q _29348_/X _30627_/S VGND VGND VPWR VPWR _30622_/A sky130_fd_sc_hd__mux2_1
X_18343_ input81/X VGND VGND VPWR VPWR _20146_/A sky130_fd_sc_hd__buf_6
XFILLER_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18274_ _34965_/Q _34901_/Q _34837_/Q _34773_/Q _16083_/X _16085_/X VGND VGND VPWR
+ VPWR _18274_/X sky130_fd_sc_hd__mux4_1
X_33340_ _33913_/CLK _33340_/D VGND VGND VPWR VPWR _33340_/Q sky130_fd_sc_hd__dfxtp_1
X_30552_ _30552_/A VGND VGND VPWR VPWR _35515_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_998 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17225_ _17221_/X _17224_/X _17151_/X VGND VGND VPWR VPWR _17235_/C sky130_fd_sc_hd__o21ba_1
X_30483_ _30483_/A VGND VGND VPWR VPWR _35482_/D sky130_fd_sc_hd__clkbuf_1
Xinput11 DW[19] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__buf_6
X_33271_ _36087_/CLK _33271_/D VGND VGND VPWR VPWR _33271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput22 DW[29] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__buf_4
XFILLER_238_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35010_ _35777_/CLK _35010_/D VGND VGND VPWR VPWR _35010_/Q sky130_fd_sc_hd__dfxtp_1
Xinput33 DW[39] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__clkbuf_8
X_32222_ _35711_/CLK _32222_/D VGND VGND VPWR VPWR _32222_/Q sky130_fd_sc_hd__dfxtp_1
Xinput44 DW[49] VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__buf_8
X_17156_ _17156_/A VGND VGND VPWR VPWR _17156_/X sky130_fd_sc_hd__clkbuf_4
Xinput55 DW[59] VGND VGND VPWR VPWR input55/X sky130_fd_sc_hd__buf_12
Xinput66 R1[1] VGND VGND VPWR VPWR input66/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput77 R3[0] VGND VGND VPWR VPWR input77/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16107_ _16107_/A VGND VGND VPWR VPWR _31958_/D sky130_fd_sc_hd__buf_4
Xinput88 RW[5] VGND VGND VPWR VPWR input88/X sky130_fd_sc_hd__buf_4
X_32153_ _35160_/CLK _32153_/D VGND VGND VPWR VPWR _32153_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17087_ _34930_/Q _34866_/Q _34802_/Q _34738_/Q _16807_/X _16808_/X VGND VGND VPWR
+ VPWR _17087_/X sky130_fd_sc_hd__mux4_1
XFILLER_66_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31104_ _35777_/Q input38/X _31116_/S VGND VGND VPWR VPWR _31105_/A sky130_fd_sc_hd__mux2_1
X_16038_ _16063_/A VGND VGND VPWR VPWR _17834_/A sky130_fd_sc_hd__buf_12
X_32084_ _35858_/CLK _32084_/D VGND VGND VPWR VPWR _32084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_486_CLK _35560_/CLK VGND VGND VPWR VPWR _35687_/CLK sky130_fd_sc_hd__clkbuf_16
X_35912_ _35976_/CLK _35912_/D VGND VGND VPWR VPWR _35912_/Q sky130_fd_sc_hd__dfxtp_1
X_31035_ _35744_/Q input2/X _31053_/S VGND VGND VPWR VPWR _31036_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35843_ _35843_/CLK _35843_/D VGND VGND VPWR VPWR _35843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17989_ _17773_/X _17987_/X _17988_/X _17777_/X VGND VGND VPWR VPWR _17989_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_238_CLK clkbuf_6_60__f_CLK/X VGND VGND VPWR VPWR _34693_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19728_ _35644_/Q _35004_/Q _34364_/Q _33724_/Q _19444_/X _19445_/X VGND VGND VPWR
+ VPWR _19728_/X sky130_fd_sc_hd__mux4_1
X_35774_ _35903_/CLK _35774_/D VGND VGND VPWR VPWR _35774_/Q sky130_fd_sc_hd__dfxtp_1
X_32986_ _34007_/CLK _32986_/D VGND VGND VPWR VPWR _32986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34725_ _34790_/CLK _34725_/D VGND VGND VPWR VPWR _34725_/Q sky130_fd_sc_hd__dfxtp_1
X_31937_ _31937_/A VGND VGND VPWR VPWR _36171_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_938 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19659_ _20169_/A VGND VGND VPWR VPWR _19659_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_52_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_246_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22670_ _34191_/Q _34127_/Q _34063_/Q _33999_/Q _22399_/X _22400_/X VGND VGND VPWR
+ VPWR _22670_/X sky130_fd_sc_hd__mux4_1
X_34656_ _35297_/CLK _34656_/D VGND VGND VPWR VPWR _34656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31868_ _31868_/A VGND VGND VPWR VPWR _36138_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_244_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33607_ _34179_/CLK _33607_/D VGND VGND VPWR VPWR _33607_/Q sky130_fd_sc_hd__dfxtp_1
X_21621_ _34161_/Q _34097_/Q _34033_/Q _33969_/Q _21340_/X _21341_/X VGND VGND VPWR
+ VPWR _21621_/X sky130_fd_sc_hd__mux4_1
X_30819_ _35642_/Q input30/X _30825_/S VGND VGND VPWR VPWR _30820_/A sky130_fd_sc_hd__mux2_1
X_34587_ _36127_/CLK _34587_/D VGND VGND VPWR VPWR _34587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31799_ _36106_/Q input48/X _31813_/S VGND VGND VPWR VPWR _31800_/A sky130_fd_sc_hd__mux2_1
XFILLER_181_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_410_CLK clkbuf_6_32__f_CLK/X VGND VGND VPWR VPWR _34098_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_90_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24340_ _24340_/A VGND VGND VPWR VPWR _32701_/D sky130_fd_sc_hd__clkbuf_1
X_33538_ _34942_/CLK _33538_/D VGND VGND VPWR VPWR _33538_/Q sky130_fd_sc_hd__dfxtp_1
X_21552_ _21446_/X _21550_/X _21551_/X _21451_/X VGND VGND VPWR VPWR _21552_/X sky130_fd_sc_hd__a22o_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20503_ _35731_/Q _32243_/Q _35603_/Q _35539_/Q _18293_/X _18295_/X VGND VGND VPWR
+ VPWR _20503_/X sky130_fd_sc_hd__mux4_1
X_24271_ _24271_/A VGND VGND VPWR VPWR _32668_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21483_ _21483_/A VGND VGND VPWR VPWR _36204_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33469_ _35449_/CLK _33469_/D VGND VGND VPWR VPWR _33469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26010_ _26010_/A VGND VGND VPWR VPWR _33459_/D sky130_fd_sc_hd__clkbuf_1
X_35208_ _35208_/CLK _35208_/D VGND VGND VPWR VPWR _35208_/Q sky130_fd_sc_hd__dfxtp_1
X_23222_ _23222_/A VGND VGND VPWR VPWR _32148_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20434_ _20212_/X _20432_/X _20433_/X _20215_/X VGND VGND VPWR VPWR _20434_/X sky130_fd_sc_hd__a22o_1
X_36188_ _36188_/CLK _36188_/D VGND VGND VPWR VPWR _36188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35139_ _35717_/CLK _35139_/D VGND VGND VPWR VPWR _35139_/Q sky130_fd_sc_hd__dfxtp_1
X_23153_ _23153_/A VGND VGND VPWR VPWR _32115_/D sky130_fd_sc_hd__clkbuf_1
XTAP_7006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20365_ _20164_/X _20363_/X _20364_/X _20169_/X VGND VGND VPWR VPWR _20365_/X sky130_fd_sc_hd__a22o_1
XFILLER_84_1108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22104_ _22457_/A VGND VGND VPWR VPWR _22104_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_136_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27961_ _27819_/X _34319_/Q _27965_/S VGND VGND VPWR VPWR _27962_/A sky130_fd_sc_hd__mux2_1
XTAP_6305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20296_ _20009_/X _20294_/X _20295_/X _20012_/X VGND VGND VPWR VPWR _20296_/X sky130_fd_sc_hd__a22o_1
X_23084_ _23084_/A VGND VGND VPWR VPWR _32085_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_477_CLK clkbuf_6_10__f_CLK/X VGND VGND VPWR VPWR _36077_/CLK sky130_fd_sc_hd__clkbuf_16
X_29700_ _29700_/A VGND VGND VPWR VPWR _35111_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_932 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26912_ _33884_/Q _23249_/X _26918_/S VGND VGND VPWR VPWR _26913_/A sky130_fd_sc_hd__mux2_1
X_22035_ _22029_/X _22034_/X _21751_/X VGND VGND VPWR VPWR _22043_/C sky130_fd_sc_hd__o21ba_1
XTAP_6349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27892_ _27717_/X _34286_/Q _27902_/S VGND VGND VPWR VPWR _27893_/A sky130_fd_sc_hd__mux2_1
XTAP_5626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29631_ _35079_/Q _29481_/X _29631_/S VGND VGND VPWR VPWR _29632_/A sky130_fd_sc_hd__mux2_1
XTAP_4903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26843_ _26843_/A VGND VGND VPWR VPWR _33851_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_229_CLK clkbuf_6_55__f_CLK/X VGND VGND VPWR VPWR _34188_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26774_ _26774_/A VGND VGND VPWR VPWR _33818_/D sky130_fd_sc_hd__clkbuf_1
X_29562_ _35046_/Q _29379_/X _29568_/S VGND VGND VPWR VPWR _29563_/A sky130_fd_sc_hd__mux2_1
X_23986_ _22894_/X _32536_/Q _24000_/S VGND VGND VPWR VPWR _23987_/A sky130_fd_sc_hd__mux2_1
XTAP_4969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28513_ _27837_/X _34581_/Q _28513_/S VGND VGND VPWR VPWR _28514_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25725_ _24868_/X _33324_/Q _25739_/S VGND VGND VPWR VPWR _25726_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22937_ input8/X VGND VGND VPWR VPWR _22937_/X sky130_fd_sc_hd__buf_2
X_29493_ _29493_/A VGND VGND VPWR VPWR _35018_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25656_ _25656_/A VGND VGND VPWR VPWR _33291_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_204_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28444_ _28513_/S VGND VGND VPWR VPWR _28463_/S sky130_fd_sc_hd__buf_4
XFILLER_95_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22868_ _20601_/X _22866_/X _22867_/X _20607_/X VGND VGND VPWR VPWR _22868_/X sky130_fd_sc_hd__a22o_1
XFILLER_227_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24607_ _23005_/X _32828_/Q _24609_/S VGND VGND VPWR VPWR _24608_/A sky130_fd_sc_hd__mux2_1
X_28375_ _28375_/A VGND VGND VPWR VPWR _34515_/D sky130_fd_sc_hd__clkbuf_1
XPHY_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21819_ _35702_/Q _32211_/Q _35574_/Q _35510_/Q _21564_/X _21565_/X VGND VGND VPWR
+ VPWR _21819_/X sky130_fd_sc_hd__mux4_1
XFILLER_58_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25587_ _25587_/A VGND VGND VPWR VPWR _33258_/D sky130_fd_sc_hd__clkbuf_1
XPHY_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22799_ _32147_/Q _32339_/Q _32403_/Q _35923_/Q _22586_/X _21611_/A VGND VGND VPWR
+ VPWR _22799_/X sky130_fd_sc_hd__mux4_1
XFILLER_12_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_401_CLK clkbuf_6_35__f_CLK/X VGND VGND VPWR VPWR _35698_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27326_ _34049_/Q _27168_/X _27338_/S VGND VGND VPWR VPWR _27327_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24538_ _22903_/X _32795_/Q _24546_/S VGND VGND VPWR VPWR _24539_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_1046 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27257_ _34016_/Q _27065_/X _27275_/S VGND VGND VPWR VPWR _27258_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24469_ _24469_/A VGND VGND VPWR VPWR _32762_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17010_ _17716_/A VGND VGND VPWR VPWR _17010_/X sky130_fd_sc_hd__buf_4
X_26208_ _26208_/A VGND VGND VPWR VPWR _33553_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27188_ _27188_/A VGND VGND VPWR VPWR _33991_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26139_ _26139_/A VGND VGND VPWR VPWR _33520_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18961_ _34406_/Q _36134_/Q _34278_/Q _34214_/Q _18823_/X _18824_/X VGND VGND VPWR
+ VPWR _18961_/X sky130_fd_sc_hd__mux4_1
XFILLER_112_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_468_CLK clkbuf_6_11__f_CLK/X VGND VGND VPWR VPWR _34926_/CLK sky130_fd_sc_hd__clkbuf_16
X_17912_ _17912_/A VGND VGND VPWR VPWR _17912_/X sky130_fd_sc_hd__buf_4
XFILLER_79_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18892_ _34916_/Q _34852_/Q _34788_/Q _34724_/Q _18754_/X _18755_/X VGND VGND VPWR
+ VPWR _18892_/X sky130_fd_sc_hd__mux4_1
XTAP_6850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17843_ _32136_/Q _32328_/Q _32392_/Q _35912_/Q _17633_/X _17774_/X VGND VGND VPWR
+ VPWR _17843_/X sky130_fd_sc_hd__mux4_1
XFILLER_21_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29829_ _29829_/A VGND VGND VPWR VPWR _35172_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32840_ _32904_/CLK _32840_/D VGND VGND VPWR VPWR _32840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17774_ _17774_/A VGND VGND VPWR VPWR _17774_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_94_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19513_ _33142_/Q _36022_/Q _33014_/Q _32950_/Q _19362_/X _19363_/X VGND VGND VPWR
+ VPWR _19513_/X sky130_fd_sc_hd__mux4_1
XFILLER_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16725_ _17935_/A VGND VGND VPWR VPWR _16725_/X sky130_fd_sc_hd__buf_6
X_32771_ _32894_/CLK _32771_/D VGND VGND VPWR VPWR _32771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34510_ _35664_/CLK _34510_/D VGND VGND VPWR VPWR _34510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31722_ _31722_/A VGND VGND VPWR VPWR _36069_/D sky130_fd_sc_hd__clkbuf_1
X_19444_ _20298_/A VGND VGND VPWR VPWR _19444_/X sky130_fd_sc_hd__buf_6
XFILLER_90_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16656_ _34662_/Q _34598_/Q _34534_/Q _34470_/Q _16586_/X _16587_/X VGND VGND VPWR
+ VPWR _16656_/X sky130_fd_sc_hd__mux4_1
X_35490_ _35490_/CLK _35490_/D VGND VGND VPWR VPWR _35490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34441_ _34441_/CLK _34441_/D VGND VGND VPWR VPWR _34441_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31653_ _27788_/X _36037_/Q _31657_/S VGND VGND VPWR VPWR _31654_/A sky130_fd_sc_hd__mux2_1
X_19375_ _35634_/Q _34994_/Q _34354_/Q _33714_/Q _19091_/X _19092_/X VGND VGND VPWR
+ VPWR _19375_/X sky130_fd_sc_hd__mux4_1
XFILLER_188_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16587_ _17999_/A VGND VGND VPWR VPWR _16587_/X sky130_fd_sc_hd__buf_4
XFILLER_76_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18326_ _33110_/Q _35990_/Q _32982_/Q _32918_/Q _18324_/X _18325_/X VGND VGND VPWR
+ VPWR _18326_/X sky130_fd_sc_hd__mux4_1
X_30604_ _30604_/A VGND VGND VPWR VPWR _35540_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_1162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34372_ _35717_/CLK _34372_/D VGND VGND VPWR VPWR _34372_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31584_ _27686_/X _36004_/Q _31594_/S VGND VGND VPWR VPWR _31585_/A sky130_fd_sc_hd__mux2_1
XFILLER_175_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36111_ _36113_/CLK _36111_/D VGND VGND VPWR VPWR _36111_/Q sky130_fd_sc_hd__dfxtp_1
X_33323_ _36075_/CLK _33323_/D VGND VGND VPWR VPWR _33323_/Q sky130_fd_sc_hd__dfxtp_1
X_18257_ _33173_/Q _36053_/Q _33045_/Q _32981_/Q _16032_/X _17161_/A VGND VGND VPWR
+ VPWR _18257_/X sky130_fd_sc_hd__mux4_1
X_30535_ _30535_/A VGND VGND VPWR VPWR _35507_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_176_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36042_ _36042_/CLK _36042_/D VGND VGND VPWR VPWR _36042_/Q sky130_fd_sc_hd__dfxtp_1
X_17208_ _33910_/Q _33846_/Q _33782_/Q _36086_/Q _17024_/X _17025_/X VGND VGND VPWR
+ VPWR _17208_/X sky130_fd_sc_hd__mux4_1
XFILLER_204_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30466_ _35475_/Q _29518_/X _30470_/S VGND VGND VPWR VPWR _30467_/A sky130_fd_sc_hd__mux2_1
X_33254_ _33697_/CLK _33254_/D VGND VGND VPWR VPWR _33254_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18188_ _18188_/A VGND VGND VPWR VPWR _32018_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_11_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32205_ _35697_/CLK _32205_/D VGND VGND VPWR VPWR _32205_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17139_ _17067_/X _17137_/X _17138_/X _17071_/X VGND VGND VPWR VPWR _17139_/X sky130_fd_sc_hd__a22o_1
X_33185_ _36065_/CLK _33185_/D VGND VGND VPWR VPWR _33185_/Q sky130_fd_sc_hd__dfxtp_1
X_30397_ _35442_/Q _29416_/X _30399_/S VGND VGND VPWR VPWR _30398_/A sky130_fd_sc_hd__mux2_1
XFILLER_239_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20150_ _20150_/A VGND VGND VPWR VPWR _20150_/X sky130_fd_sc_hd__buf_4
XFILLER_89_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32136_ _32905_/CLK _32136_/D VGND VGND VPWR VPWR _32136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_459_CLK clkbuf_leaf_49_CLK/A VGND VGND VPWR VPWR _35753_/CLK sky130_fd_sc_hd__clkbuf_16
X_20081_ _35654_/Q _35014_/Q _34374_/Q _33734_/Q _19797_/X _19798_/X VGND VGND VPWR
+ VPWR _20081_/X sky130_fd_sc_hd__mux4_1
XFILLER_174_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32067_ _35779_/CLK _32067_/D VGND VGND VPWR VPWR _32067_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31018_ _35736_/Q input23/X _31032_/S VGND VGND VPWR VPWR _31019_/A sky130_fd_sc_hd__mux2_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23840_ _23082_/X _32405_/Q _23840_/S VGND VGND VPWR VPWR _23841_/A sky130_fd_sc_hd__mux2_1
XTAP_3509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35826_ _36147_/CLK _35826_/D VGND VGND VPWR VPWR _35826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_245_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35757_ _36013_/CLK _35757_/D VGND VGND VPWR VPWR _35757_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23771_ _23840_/S VGND VGND VPWR VPWR _23790_/S sky130_fd_sc_hd__buf_4
X_20983_ _20979_/X _20982_/X _20704_/X VGND VGND VPWR VPWR _20984_/D sky130_fd_sc_hd__o21ba_1
X_32969_ _36044_/CLK _32969_/D VGND VGND VPWR VPWR _32969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25510_ _25510_/A VGND VGND VPWR VPWR _33222_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22722_ _22459_/X _22720_/X _22721_/X _22462_/X VGND VGND VPWR VPWR _22722_/X sky130_fd_sc_hd__a22o_1
X_34708_ _34708_/CLK _34708_/D VGND VGND VPWR VPWR _34708_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_246_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26490_ _26622_/S VGND VGND VPWR VPWR _26509_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_25_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35688_ _35690_/CLK _35688_/D VGND VGND VPWR VPWR _35688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25441_ _25441_/A VGND VGND VPWR VPWR _33189_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_241_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34639_ _35147_/CLK _34639_/D VGND VGND VPWR VPWR _34639_/Q sky130_fd_sc_hd__dfxtp_1
X_22653_ _35726_/Q _32237_/Q _35598_/Q _35534_/Q _20593_/X _20595_/X VGND VGND VPWR
+ VPWR _22653_/X sky130_fd_sc_hd__mux4_1
XFILLER_53_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_240_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21604_ _35440_/Q _35376_/Q _35312_/Q _35248_/Q _21501_/X _21502_/X VGND VGND VPWR
+ VPWR _21604_/X sky130_fd_sc_hd__mux4_1
X_28160_ _27714_/X _34413_/Q _28172_/S VGND VGND VPWR VPWR _28161_/A sky130_fd_sc_hd__mux2_1
X_25372_ _33158_/Q _23447_/X _25374_/S VGND VGND VPWR VPWR _25373_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22584_ _33164_/Q _36044_/Q _33036_/Q _32972_/Q _22368_/X _22369_/X VGND VGND VPWR
+ VPWR _22584_/X sky130_fd_sc_hd__mux4_1
X_27111_ _27111_/A VGND VGND VPWR VPWR _33966_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24323_ _22984_/X _32693_/Q _24339_/S VGND VGND VPWR VPWR _24324_/A sky130_fd_sc_hd__mux2_1
X_28091_ _28091_/A VGND VGND VPWR VPWR _34380_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21535_ _35438_/Q _35374_/Q _35310_/Q _35246_/Q _21501_/X _21502_/X VGND VGND VPWR
+ VPWR _21535_/X sky130_fd_sc_hd__mux4_1
XFILLER_193_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27042_ _33944_/Q _27041_/X _27063_/S VGND VGND VPWR VPWR _27043_/A sky130_fd_sc_hd__mux2_1
X_24254_ _24254_/A VGND VGND VPWR VPWR _31553_/B sky130_fd_sc_hd__buf_12
XFILLER_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21466_ _35692_/Q _32200_/Q _35564_/Q _35500_/Q _21211_/X _21212_/X VGND VGND VPWR
+ VPWR _21466_/X sky130_fd_sc_hd__mux4_1
XFILLER_107_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23205_ _23055_/X _32140_/Q _23215_/S VGND VGND VPWR VPWR _23206_/A sky130_fd_sc_hd__mux2_1
X_20417_ _33104_/Q _32080_/Q _35856_/Q _35792_/Q _18379_/X _18380_/X VGND VGND VPWR
+ VPWR _20417_/X sky130_fd_sc_hd__mux4_1
X_24185_ _32629_/Q _23393_/X _24201_/S VGND VGND VPWR VPWR _24186_/A sky130_fd_sc_hd__mux2_1
XFILLER_218_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21397_ _21250_/X _21395_/X _21396_/X _21253_/X VGND VGND VPWR VPWR _21397_/X sky130_fd_sc_hd__a22o_1
XFILLER_218_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23136_ _22953_/X _32107_/Q _23152_/S VGND VGND VPWR VPWR _23137_/A sky130_fd_sc_hd__mux2_1
X_20348_ _20065_/X _20346_/X _20347_/X _20071_/X VGND VGND VPWR VPWR _20348_/X sky130_fd_sc_hd__a22o_1
XTAP_6102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28993_ _28993_/A VGND VGND VPWR VPWR _34806_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27944_ _27794_/X _34311_/Q _27944_/S VGND VGND VPWR VPWR _27945_/A sky130_fd_sc_hd__mux2_1
XFILLER_175_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23067_ input54/X VGND VGND VPWR VPWR _23067_/X sky130_fd_sc_hd__buf_2
XFILLER_0_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20279_ _33932_/Q _33868_/Q _33804_/Q _36108_/Q _20030_/X _20031_/X VGND VGND VPWR
+ VPWR _20279_/X sky130_fd_sc_hd__mux4_1
XTAP_6146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22018_ _22510_/A VGND VGND VPWR VPWR _22018_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_68_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27875_ _27692_/X _34278_/Q _27881_/S VGND VGND VPWR VPWR _27876_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29614_ _29614_/A VGND VGND VPWR VPWR _35070_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26826_ _26826_/A VGND VGND VPWR VPWR _33843_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29545_ _35038_/Q _29354_/X _29547_/S VGND VGND VPWR VPWR _29546_/A sky130_fd_sc_hd__mux2_1
XTAP_4788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26757_ _33811_/Q _23492_/X _26761_/S VGND VGND VPWR VPWR _26758_/A sky130_fd_sc_hd__mux2_1
X_23969_ _23070_/X _32529_/Q _23969_/S VGND VGND VPWR VPWR _23970_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16510_ _32866_/Q _32802_/Q _32738_/Q _32674_/Q _16287_/X _16288_/X VGND VGND VPWR
+ VPWR _16510_/X sky130_fd_sc_hd__mux4_1
X_25708_ _24843_/X _33316_/Q _25718_/S VGND VGND VPWR VPWR _25709_/A sky130_fd_sc_hd__mux2_1
X_29476_ _35013_/Q _29475_/X _29482_/S VGND VGND VPWR VPWR _29477_/A sky130_fd_sc_hd__mux2_1
X_17490_ _32126_/Q _32318_/Q _32382_/Q _35902_/Q _17280_/X _17421_/X VGND VGND VPWR
+ VPWR _17490_/X sky130_fd_sc_hd__mux4_1
X_26688_ _33778_/Q _23381_/X _26690_/S VGND VGND VPWR VPWR _26689_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28427_ _28427_/A VGND VGND VPWR VPWR _34539_/D sky130_fd_sc_hd__clkbuf_1
X_16441_ _16292_/X _16437_/X _16440_/X _16295_/X VGND VGND VPWR VPWR _16441_/X sky130_fd_sc_hd__a22o_1
X_25639_ _25639_/A VGND VGND VPWR VPWR _33283_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_1048 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16372_ _17935_/A VGND VGND VPWR VPWR _16372_/X sky130_fd_sc_hd__buf_6
X_19160_ _33132_/Q _36012_/Q _33004_/Q _32940_/Q _19009_/X _19010_/X VGND VGND VPWR
+ VPWR _19160_/X sky130_fd_sc_hd__mux4_1
X_28358_ _27807_/X _34507_/Q _28370_/S VGND VGND VPWR VPWR _28359_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18111_ _17158_/A _18109_/X _18110_/X _17163_/A VGND VGND VPWR VPWR _18111_/X sky130_fd_sc_hd__a22o_1
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27309_ _34041_/Q _27143_/X _27317_/S VGND VGND VPWR VPWR _27310_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_1477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19091_ _20298_/A VGND VGND VPWR VPWR _19091_/X sky130_fd_sc_hd__buf_6
X_28289_ _27704_/X _34474_/Q _28307_/S VGND VGND VPWR VPWR _28290_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30320_ _30320_/A VGND VGND VPWR VPWR _35405_/D sky130_fd_sc_hd__clkbuf_1
X_18042_ _33422_/Q _33358_/Q _33294_/Q _33230_/Q _17833_/X _17834_/X VGND VGND VPWR
+ VPWR _18042_/X sky130_fd_sc_hd__mux4_1
XFILLER_201_1332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30251_ _30251_/A VGND VGND VPWR VPWR _35372_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_1406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30182_ _35340_/Q _29497_/X _30192_/S VGND VGND VPWR VPWR _30183_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19993_ _19859_/X _19991_/X _19992_/X _19862_/X VGND VGND VPWR VPWR _19993_/X sky130_fd_sc_hd__a22o_1
XFILLER_28_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18944_ _18938_/X _18943_/X _18734_/X _18735_/X VGND VGND VPWR VPWR _18965_/B sky130_fd_sc_hd__o211a_2
X_34990_ _35694_/CLK _34990_/D VGND VGND VPWR VPWR _34990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33941_ _33941_/CLK _33941_/D VGND VGND VPWR VPWR _33941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18875_ _32100_/Q _32292_/Q _32356_/Q _35876_/Q _18874_/X _18662_/X VGND VGND VPWR
+ VPWR _18875_/X sky130_fd_sc_hd__mux4_1
XTAP_6680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17826_ _17511_/X _17824_/X _17825_/X _17516_/X VGND VGND VPWR VPWR _17826_/X sky130_fd_sc_hd__a22o_1
X_33872_ _34440_/CLK _33872_/D VGND VGND VPWR VPWR _33872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35611_ _35802_/CLK _35611_/D VGND VGND VPWR VPWR _35611_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_616 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32823_ _32885_/CLK _32823_/D VGND VGND VPWR VPWR _32823_/Q sky130_fd_sc_hd__dfxtp_1
X_17757_ _17757_/A VGND VGND VPWR VPWR _32005_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_94_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35542_ _35735_/CLK _35542_/D VGND VGND VPWR VPWR _35542_/Q sky130_fd_sc_hd__dfxtp_1
X_16708_ _32616_/Q _32552_/Q _32488_/Q _35944_/Q _16570_/X _16707_/X VGND VGND VPWR
+ VPWR _16708_/X sky130_fd_sc_hd__mux4_1
X_32754_ _32818_/CLK _32754_/D VGND VGND VPWR VPWR _32754_/Q sky130_fd_sc_hd__dfxtp_1
X_17688_ _33668_/Q _33604_/Q _33540_/Q _33476_/Q _17553_/X _17554_/X VGND VGND VPWR
+ VPWR _17688_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31705_ _31705_/A VGND VGND VPWR VPWR _36061_/D sky130_fd_sc_hd__clkbuf_1
X_19427_ _20133_/A VGND VGND VPWR VPWR _19427_/X sky130_fd_sc_hd__buf_4
X_35473_ _35855_/CLK _35473_/D VGND VGND VPWR VPWR _35473_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16639_ _32102_/Q _32294_/Q _32358_/Q _35878_/Q _16574_/X _16362_/X VGND VGND VPWR
+ VPWR _16639_/X sky130_fd_sc_hd__mux4_1
X_32685_ _32877_/CLK _32685_/D VGND VGND VPWR VPWR _32685_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34424_ _35192_/CLK _34424_/D VGND VGND VPWR VPWR _34424_/Q sky130_fd_sc_hd__dfxtp_1
X_19358_ _19354_/X _19357_/X _19079_/X VGND VGND VPWR VPWR _19390_/A sky130_fd_sc_hd__o21ba_1
X_31636_ _27763_/X _36029_/Q _31636_/S VGND VGND VPWR VPWR _31637_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18309_ _20260_/A VGND VGND VPWR VPWR _18309_/X sky130_fd_sc_hd__buf_6
XFILLER_200_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34355_ _35632_/CLK _34355_/D VGND VGND VPWR VPWR _34355_/Q sky130_fd_sc_hd__dfxtp_1
X_31567_ _27661_/X _35996_/Q _31573_/S VGND VGND VPWR VPWR _31568_/A sky130_fd_sc_hd__mux2_1
X_19289_ _32624_/Q _32560_/Q _32496_/Q _35952_/Q _19223_/X _19007_/X VGND VGND VPWR
+ VPWR _19289_/X sky130_fd_sc_hd__mux4_1
XFILLER_176_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33306_ _33818_/CLK _33306_/D VGND VGND VPWR VPWR _33306_/Q sky130_fd_sc_hd__dfxtp_1
X_21320_ _21313_/X _21319_/X _21034_/X _21035_/X VGND VGND VPWR VPWR _21337_/B sky130_fd_sc_hd__o211a_1
XFILLER_108_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30518_ _35499_/Q _29395_/X _30534_/S VGND VGND VPWR VPWR _30519_/A sky130_fd_sc_hd__mux2_1
X_34286_ _36142_/CLK _34286_/D VGND VGND VPWR VPWR _34286_/Q sky130_fd_sc_hd__dfxtp_1
X_31498_ _31498_/A VGND VGND VPWR VPWR _35963_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36025_ _36025_/CLK _36025_/D VGND VGND VPWR VPWR _36025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33237_ _33685_/CLK _33237_/D VGND VGND VPWR VPWR _33237_/Q sky130_fd_sc_hd__dfxtp_1
X_21251_ _35430_/Q _35366_/Q _35302_/Q _35238_/Q _21148_/X _21149_/X VGND VGND VPWR
+ VPWR _21251_/X sky130_fd_sc_hd__mux4_1
X_30449_ _30449_/A VGND VGND VPWR VPWR _35466_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20202_ _20198_/X _20201_/X _20171_/X VGND VGND VPWR VPWR _20203_/D sky130_fd_sc_hd__o21ba_1
XFILLER_132_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33168_ _36047_/CLK _33168_/D VGND VGND VPWR VPWR _33168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21182_ _35428_/Q _35364_/Q _35300_/Q _35236_/Q _21148_/X _21149_/X VGND VGND VPWR
+ VPWR _21182_/X sky130_fd_sc_hd__mux4_1
XFILLER_144_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20133_ _20133_/A VGND VGND VPWR VPWR _20133_/X sky130_fd_sc_hd__buf_4
XFILLER_137_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32119_ _35895_/CLK _32119_/D VGND VGND VPWR VPWR _32119_/Q sky130_fd_sc_hd__dfxtp_1
X_25990_ _26080_/S VGND VGND VPWR VPWR _26009_/S sky130_fd_sc_hd__buf_4
X_33099_ _35852_/CLK _33099_/D VGND VGND VPWR VPWR _33099_/Q sky130_fd_sc_hd__dfxtp_1
X_20064_ _20060_/X _20063_/X _19785_/X VGND VGND VPWR VPWR _20096_/A sky130_fd_sc_hd__o21ba_2
X_24941_ _24941_/A VGND VGND VPWR VPWR _32963_/D sky130_fd_sc_hd__clkbuf_1
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27660_ _27660_/A VGND VGND VPWR VPWR _34203_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24872_ _24871_/X _32941_/Q _24890_/S VGND VGND VPWR VPWR _24873_/A sky130_fd_sc_hd__mux2_1
XTAP_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1018 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26611_ _26611_/A VGND VGND VPWR VPWR _33743_/D sky130_fd_sc_hd__clkbuf_1
X_23823_ _23823_/A VGND VGND VPWR VPWR _32396_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27591_ _27591_/A VGND VGND VPWR VPWR _34174_/D sky130_fd_sc_hd__clkbuf_1
X_35809_ _36007_/CLK _35809_/D VGND VGND VPWR VPWR _35809_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29330_ _29525_/S VGND VGND VPWR VPWR _29358_/S sky130_fd_sc_hd__clkbuf_8
X_26542_ _26542_/A VGND VGND VPWR VPWR _33710_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23754_ _23754_/A VGND VGND VPWR VPWR _32363_/D sky130_fd_sc_hd__clkbuf_1
X_20966_ _20961_/X _20963_/X _20964_/X _20965_/X VGND VGND VPWR VPWR _20966_/X sky130_fd_sc_hd__a22o_1
XFILLER_187_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22705_ _22701_/X _22704_/X _22438_/X VGND VGND VPWR VPWR _22727_/A sky130_fd_sc_hd__o21ba_1
XFILLER_26_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26473_ _26473_/A VGND VGND VPWR VPWR _33678_/D sky130_fd_sc_hd__clkbuf_1
X_29261_ _29261_/A VGND VGND VPWR VPWR _34933_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23685_ _23685_/A VGND VGND VPWR VPWR _32332_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20897_ _22464_/A VGND VGND VPWR VPWR _20897_/X sky130_fd_sc_hd__buf_4
XFILLER_213_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28212_ _27791_/X _34438_/Q _28214_/S VGND VGND VPWR VPWR _28213_/A sky130_fd_sc_hd__mux2_1
X_25424_ _25424_/A VGND VGND VPWR VPWR _33181_/D sky130_fd_sc_hd__clkbuf_1
X_29192_ _29192_/A VGND VGND VPWR VPWR _34901_/D sky130_fd_sc_hd__clkbuf_1
X_22636_ _22632_/X _22635_/X _22471_/X VGND VGND VPWR VPWR _22637_/D sky130_fd_sc_hd__o21ba_1
XFILLER_16_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_1354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25355_ _25403_/S VGND VGND VPWR VPWR _25374_/S sky130_fd_sc_hd__buf_4
X_28143_ _27689_/X _34405_/Q _28151_/S VGND VGND VPWR VPWR _28144_/A sky130_fd_sc_hd__mux2_1
X_22567_ _35211_/Q _35147_/Q _35083_/Q _32267_/Q _22316_/X _22317_/X VGND VGND VPWR
+ VPWR _22567_/X sky130_fd_sc_hd__mux4_1
XFILLER_194_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24306_ _22959_/X _32685_/Q _24318_/S VGND VGND VPWR VPWR _24307_/A sky130_fd_sc_hd__mux2_1
X_28074_ _28074_/A VGND VGND VPWR VPWR _34372_/D sky130_fd_sc_hd__clkbuf_1
X_21518_ _21446_/X _21516_/X _21517_/X _21451_/X VGND VGND VPWR VPWR _21518_/X sky130_fd_sc_hd__a22o_1
X_25286_ _33117_/Q _23252_/X _25290_/S VGND VGND VPWR VPWR _25287_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_1371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22498_ _22459_/X _22496_/X _22497_/X _22462_/X VGND VGND VPWR VPWR _22498_/X sky130_fd_sc_hd__a22o_1
XFILLER_177_1106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27025_ _33938_/Q _23487_/X _27031_/S VGND VGND VPWR VPWR _27026_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24237_ _32654_/Q _23475_/X _24243_/S VGND VGND VPWR VPWR _24238_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21449_ _33644_/Q _33580_/Q _33516_/Q _33452_/Q _21447_/X _21448_/X VGND VGND VPWR
+ VPWR _21449_/X sky130_fd_sc_hd__mux4_1
XFILLER_163_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_824 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24168_ _32621_/Q _23302_/X _24180_/S VGND VGND VPWR VPWR _24169_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23119_ _22928_/X _32099_/Q _23131_/S VGND VGND VPWR VPWR _23120_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24099_ _23061_/X _32590_/Q _24105_/S VGND VGND VPWR VPWR _24100_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28976_ _28976_/A VGND VGND VPWR VPWR _34798_/D sky130_fd_sc_hd__clkbuf_1
X_16990_ _33136_/Q _36016_/Q _33008_/Q _32944_/Q _16709_/X _16710_/X VGND VGND VPWR
+ VPWR _16990_/X sky130_fd_sc_hd__mux4_1
X_27927_ _27927_/A VGND VGND VPWR VPWR _34302_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18660_ _18653_/X _18655_/X _18658_/X _18659_/X VGND VGND VPWR VPWR _18660_/X sky130_fd_sc_hd__a22o_1
X_27858_ _27667_/X _34270_/Q _27860_/S VGND VGND VPWR VPWR _27859_/A sky130_fd_sc_hd__mux2_1
XFILLER_188_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17611_ _17356_/X _17609_/X _17610_/X _17359_/X VGND VGND VPWR VPWR _17611_/X sky130_fd_sc_hd__a22o_1
XFILLER_36_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26809_ _33835_/Q _23296_/X _26825_/S VGND VGND VPWR VPWR _26810_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18591_ _18585_/X _18590_/X _18344_/X _18346_/X VGND VGND VPWR VPWR _18612_/B sky130_fd_sc_hd__o211a_1
XTAP_4574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27789_ _27788_/X _34245_/Q _27795_/S VGND VGND VPWR VPWR _27790_/A sky130_fd_sc_hd__mux2_1
XTAP_4585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29528_ _29660_/S VGND VGND VPWR VPWR _29547_/S sky130_fd_sc_hd__buf_6
X_17542_ _17538_/X _17541_/X _17504_/X VGND VGND VPWR VPWR _17550_/C sky130_fd_sc_hd__o21ba_1
XTAP_3873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_225_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29459_ _29459_/A VGND VGND VPWR VPWR _35007_/D sky130_fd_sc_hd__clkbuf_1
X_17473_ _17158_/X _17471_/X _17472_/X _17163_/X VGND VGND VPWR VPWR _17473_/X sky130_fd_sc_hd__a22o_1
XFILLER_233_986 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19212_ _19105_/X _19210_/X _19211_/X _19110_/X VGND VGND VPWR VPWR _19212_/X sky130_fd_sc_hd__a22o_1
X_16424_ _33888_/Q _33824_/Q _33760_/Q _36064_/Q _16318_/X _16319_/X VGND VGND VPWR
+ VPWR _16424_/X sky130_fd_sc_hd__mux4_1
XFILLER_73_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32470_ _35990_/CLK _32470_/D VGND VGND VPWR VPWR _32470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31421_ _31421_/A VGND VGND VPWR VPWR _35926_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_1132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19143_ _19139_/X _19142_/X _19112_/X VGND VGND VPWR VPWR _19144_/D sky130_fd_sc_hd__o21ba_1
X_16355_ _32606_/Q _32542_/Q _32478_/Q _35934_/Q _16217_/X _16354_/X VGND VGND VPWR
+ VPWR _16355_/X sky130_fd_sc_hd__mux4_1
XFILLER_199_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34140_ _36211_/CLK _34140_/D VGND VGND VPWR VPWR _34140_/Q sky130_fd_sc_hd__dfxtp_1
X_16286_ _32092_/Q _32284_/Q _32348_/Q _35868_/Q _16221_/X _17867_/A VGND VGND VPWR
+ VPWR _16286_/X sky130_fd_sc_hd__mux4_1
X_19074_ _20133_/A VGND VGND VPWR VPWR _19074_/X sky130_fd_sc_hd__buf_4
X_31352_ _27742_/X _35894_/Q _31366_/S VGND VGND VPWR VPWR _31353_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18025_ _17704_/X _18023_/X _18024_/X _17707_/X VGND VGND VPWR VPWR _18025_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30303_ _30303_/A VGND VGND VPWR VPWR _35397_/D sky130_fd_sc_hd__clkbuf_1
X_34071_ _34135_/CLK _34071_/D VGND VGND VPWR VPWR _34071_/Q sky130_fd_sc_hd__dfxtp_1
X_31283_ _31418_/A _31283_/B VGND VGND VPWR VPWR _31416_/S sky130_fd_sc_hd__nand2_8
XFILLER_160_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33022_ _35839_/CLK _33022_/D VGND VGND VPWR VPWR _33022_/Q sky130_fd_sc_hd__dfxtp_1
X_30234_ _30234_/A VGND VGND VPWR VPWR _35364_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30165_ _35332_/Q _29472_/X _30171_/S VGND VGND VPWR VPWR _30166_/A sky130_fd_sc_hd__mux2_1
X_19976_ _33091_/Q _32067_/Q _35843_/Q _35779_/Q _19731_/X _19732_/X VGND VGND VPWR
+ VPWR _19976_/X sky130_fd_sc_hd__mux4_1
XFILLER_113_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18927_ _18927_/A _18927_/B _18927_/C _18927_/D VGND VGND VPWR VPWR _18928_/A sky130_fd_sc_hd__or4_2
X_34973_ _36060_/CLK _34973_/D VGND VGND VPWR VPWR _34973_/Q sky130_fd_sc_hd__dfxtp_1
X_30096_ _35299_/Q _29370_/X _30108_/S VGND VGND VPWR VPWR _30097_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_955 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33924_ _33924_/CLK _33924_/D VGND VGND VPWR VPWR _33924_/Q sky130_fd_sc_hd__dfxtp_1
X_18858_ _34915_/Q _34851_/Q _34787_/Q _34723_/Q _18754_/X _18755_/X VGND VGND VPWR
+ VPWR _18858_/X sky130_fd_sc_hd__mux4_1
XFILLER_68_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17809_ _17765_/X _17807_/X _17808_/X _17771_/X VGND VGND VPWR VPWR _17809_/X sky130_fd_sc_hd__a22o_1
XFILLER_209_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33855_ _36095_/CLK _33855_/D VGND VGND VPWR VPWR _33855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18789_ _18752_/X _18787_/X _18788_/X _18757_/X VGND VGND VPWR VPWR _18789_/X sky130_fd_sc_hd__a22o_1
XFILLER_227_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_247_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20820_ _20618_/X _20818_/X _20819_/X _20627_/X VGND VGND VPWR VPWR _20820_/X sky130_fd_sc_hd__a22o_1
X_32806_ _32808_/CLK _32806_/D VGND VGND VPWR VPWR _32806_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33786_ _36090_/CLK _33786_/D VGND VGND VPWR VPWR _33786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_247_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30998_ _35727_/Q input53/X _31002_/S VGND VGND VPWR VPWR _30999_/A sky130_fd_sc_hd__mux2_1
XFILLER_223_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35525_ _35525_/CLK _35525_/D VGND VGND VPWR VPWR _35525_/Q sky130_fd_sc_hd__dfxtp_1
X_20751_ _20747_/X _20748_/X _20749_/X _20750_/X VGND VGND VPWR VPWR _20751_/X sky130_fd_sc_hd__a22o_1
X_32737_ _35875_/CLK _32737_/D VGND VGND VPWR VPWR _32737_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_997 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23470_ _32235_/Q _23469_/X _23485_/S VGND VGND VPWR VPWR _23471_/A sky130_fd_sc_hd__mux2_1
X_35456_ _35456_/CLK _35456_/D VGND VGND VPWR VPWR _35456_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32668_ _36053_/CLK _32668_/D VGND VGND VPWR VPWR _32668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20682_ _22582_/A VGND VGND VPWR VPWR _22316_/A sky130_fd_sc_hd__buf_12
XFILLER_195_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22421_ _34695_/Q _34631_/Q _34567_/Q _34503_/Q _22245_/X _22246_/X VGND VGND VPWR
+ VPWR _22421_/X sky130_fd_sc_hd__mux4_1
X_34407_ _36135_/CLK _34407_/D VGND VGND VPWR VPWR _34407_/Q sky130_fd_sc_hd__dfxtp_1
X_31619_ _31619_/A VGND VGND VPWR VPWR _36020_/D sky130_fd_sc_hd__clkbuf_1
X_35387_ _35581_/CLK _35387_/D VGND VGND VPWR VPWR _35387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32599_ _35929_/CLK _32599_/D VGND VGND VPWR VPWR _32599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25140_ _33048_/Q _23237_/X _25154_/S VGND VGND VPWR VPWR _25141_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22352_ _34437_/Q _36165_/Q _34309_/Q _34245_/Q _22182_/X _22183_/X VGND VGND VPWR
+ VPWR _22352_/X sky130_fd_sc_hd__mux4_1
X_34338_ _34921_/CLK _34338_/D VGND VGND VPWR VPWR _34338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21303_ _33896_/Q _33832_/Q _33768_/Q _36072_/Q _21271_/X _21272_/X VGND VGND VPWR
+ VPWR _21303_/X sky130_fd_sc_hd__mux4_1
XFILLER_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25071_ _25071_/A VGND VGND VPWR VPWR _33016_/D sky130_fd_sc_hd__clkbuf_1
X_34269_ _36235_/CLK _34269_/D VGND VGND VPWR VPWR _34269_/Q sky130_fd_sc_hd__dfxtp_1
X_22283_ _34947_/Q _34883_/Q _34819_/Q _34755_/Q _22113_/X _22114_/X VGND VGND VPWR
+ VPWR _22283_/X sky130_fd_sc_hd__mux4_1
XFILLER_156_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36008_ _36011_/CLK _36008_/D VGND VGND VPWR VPWR _36008_/Q sky130_fd_sc_hd__dfxtp_1
X_24022_ _24022_/A VGND VGND VPWR VPWR _32553_/D sky130_fd_sc_hd__clkbuf_1
X_21234_ _21100_/X _21232_/X _21233_/X _21103_/X VGND VGND VPWR VPWR _21234_/X sky130_fd_sc_hd__a22o_1
XFILLER_102_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28830_ _28830_/A VGND VGND VPWR VPWR _34729_/D sky130_fd_sc_hd__clkbuf_1
X_21165_ _21093_/X _21163_/X _21164_/X _21098_/X VGND VGND VPWR VPWR _21165_/X sky130_fd_sc_hd__a22o_1
XFILLER_104_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20116_ _20004_/X _20114_/X _20115_/X _20007_/X VGND VGND VPWR VPWR _20116_/X sky130_fd_sc_hd__a22o_1
XFILLER_132_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28761_ _28761_/A VGND VGND VPWR VPWR _34697_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21096_ _33634_/Q _33570_/Q _33506_/Q _33442_/Q _21094_/X _21095_/X VGND VGND VPWR
+ VPWR _21096_/X sky130_fd_sc_hd__mux4_1
XFILLER_28_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25973_ _25973_/A VGND VGND VPWR VPWR _33441_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_246_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27712_ _27711_/X _34220_/Q _27733_/S VGND VGND VPWR VPWR _27713_/A sky130_fd_sc_hd__mux2_1
X_20047_ _20009_/X _20045_/X _20046_/X _20012_/X VGND VGND VPWR VPWR _20047_/X sky130_fd_sc_hd__a22o_1
XFILLER_150_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24924_ _24995_/S VGND VGND VPWR VPWR _24952_/S sky130_fd_sc_hd__buf_6
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28692_ _34665_/Q _27093_/X _28692_/S VGND VGND VPWR VPWR _28693_/A sky130_fd_sc_hd__mux2_1
XTAP_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27643_ _27838_/S VGND VGND VPWR VPWR _27671_/S sky130_fd_sc_hd__buf_4
XTAP_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24855_ input10/X VGND VGND VPWR VPWR _24855_/X sky130_fd_sc_hd__buf_4
XTAP_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23806_ _23806_/A VGND VGND VPWR VPWR _32388_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24786_ _23070_/X _32913_/Q _24786_/S VGND VGND VPWR VPWR _24787_/A sky130_fd_sc_hd__mux2_1
X_27574_ _27574_/A VGND VGND VPWR VPWR _34166_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21998_ _21753_/X _21996_/X _21997_/X _21756_/X VGND VGND VPWR VPWR _21998_/X sky130_fd_sc_hd__a22o_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29313_ _29313_/A VGND VGND VPWR VPWR _34958_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26525_ _26525_/A VGND VGND VPWR VPWR _33702_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23737_ _23737_/A VGND VGND VPWR VPWR _32355_/D sky130_fd_sc_hd__clkbuf_1
X_20949_ _33374_/Q _33310_/Q _33246_/Q _33182_/Q _20602_/X _20603_/X VGND VGND VPWR
+ VPWR _20949_/X sky130_fd_sc_hd__mux4_1
XFILLER_54_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_1108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29244_ _29244_/A VGND VGND VPWR VPWR _34925_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26456_ _26456_/A VGND VGND VPWR VPWR _33670_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23668_ _23668_/A VGND VGND VPWR VPWR _32324_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25407_ _31283_/B _26352_/B VGND VGND VPWR VPWR _25540_/S sky130_fd_sc_hd__nand2_8
X_22619_ _32141_/Q _32333_/Q _32397_/Q _35917_/Q _22586_/X _22374_/X VGND VGND VPWR
+ VPWR _22619_/X sky130_fd_sc_hd__mux4_1
XFILLER_74_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29175_ _34893_/Q _27205_/X _29183_/S VGND VGND VPWR VPWR _29176_/A sky130_fd_sc_hd__mux2_1
XFILLER_197_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26387_ _26387_/A VGND VGND VPWR VPWR _33637_/D sky130_fd_sc_hd__clkbuf_1
X_23599_ _23599_/A VGND VGND VPWR VPWR _32291_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16140_ _17859_/A VGND VGND VPWR VPWR _16140_/X sky130_fd_sc_hd__buf_4
XFILLER_10_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28126_ _27664_/X _34397_/Q _28130_/S VGND VGND VPWR VPWR _28127_/A sky130_fd_sc_hd__mux2_1
XFILLER_220_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25338_ _25338_/A VGND VGND VPWR VPWR _33141_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16071_ _17777_/A VGND VGND VPWR VPWR _17869_/A sky130_fd_sc_hd__buf_12
XFILLER_182_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25269_ _30877_/B _31553_/B VGND VGND VPWR VPWR _25270_/A sky130_fd_sc_hd__and2b_1
X_28057_ _28057_/A VGND VGND VPWR VPWR _34364_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27008_ _27008_/A VGND VGND VPWR VPWR _33929_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19830_ _33151_/Q _36031_/Q _33023_/Q _32959_/Q _19715_/X _19716_/X VGND VGND VPWR
+ VPWR _19830_/X sky130_fd_sc_hd__mux4_1
XFILLER_64_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19761_ _35709_/Q _32218_/Q _35581_/Q _35517_/Q _19617_/X _19618_/X VGND VGND VPWR
+ VPWR _19761_/X sky130_fd_sc_hd__mux4_1
X_28959_ _28959_/A VGND VGND VPWR VPWR _34790_/D sky130_fd_sc_hd__clkbuf_1
X_16973_ _34671_/Q _34607_/Q _34543_/Q _34479_/Q _16939_/X _16940_/X VGND VGND VPWR
+ VPWR _16973_/X sky130_fd_sc_hd__mux4_1
XFILLER_49_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18712_ _34399_/Q _36127_/Q _34271_/Q _34207_/Q _18470_/X _18471_/X VGND VGND VPWR
+ VPWR _18712_/X sky130_fd_sc_hd__mux4_1
XTAP_5050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31970_ _34085_/CLK _31970_/D VGND VGND VPWR VPWR _31970_/Q sky130_fd_sc_hd__dfxtp_1
X_19692_ _35451_/Q _35387_/Q _35323_/Q _35259_/Q _19554_/X _19555_/X VGND VGND VPWR
+ VPWR _19692_/X sky130_fd_sc_hd__mux4_1
XFILLER_237_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_231_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput9 DW[17] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__buf_6
XFILLER_92_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18643_ _18639_/X _18642_/X _18404_/X VGND VGND VPWR VPWR _18644_/D sky130_fd_sc_hd__o21ba_1
XTAP_5094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30921_ _35690_/Q input13/X _30939_/S VGND VGND VPWR VPWR _30922_/A sky130_fd_sc_hd__mux2_1
XFILLER_225_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33640_ _35624_/CLK _33640_/D VGND VGND VPWR VPWR _33640_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30852_ _30852_/A VGND VGND VPWR VPWR _35657_/D sky130_fd_sc_hd__clkbuf_1
X_18574_ _18574_/A _18574_/B _18574_/C _18574_/D VGND VGND VPWR VPWR _18575_/A sky130_fd_sc_hd__or4_1
XFILLER_18_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17525_ _33407_/Q _33343_/Q _33279_/Q _33215_/Q _17480_/X _17481_/X VGND VGND VPWR
+ VPWR _17525_/X sky130_fd_sc_hd__mux4_1
XFILLER_229_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33571_ _34151_/CLK _33571_/D VGND VGND VPWR VPWR _33571_/Q sky130_fd_sc_hd__dfxtp_1
X_30783_ _35625_/Q input11/X _30783_/S VGND VGND VPWR VPWR _30784_/A sky130_fd_sc_hd__mux2_1
XFILLER_233_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_923 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35310_ _35438_/CLK _35310_/D VGND VGND VPWR VPWR _35310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32522_ _35978_/CLK _32522_/D VGND VGND VPWR VPWR _32522_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17456_ _17412_/X _17454_/X _17455_/X _17418_/X VGND VGND VPWR VPWR _17456_/X sky130_fd_sc_hd__a22o_1
XFILLER_177_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16407_ _16297_/X _16405_/X _16406_/X _16300_/X VGND VGND VPWR VPWR _16407_/X sky130_fd_sc_hd__a22o_1
X_35241_ _35433_/CLK _35241_/D VGND VGND VPWR VPWR _35241_/Q sky130_fd_sc_hd__dfxtp_1
X_32453_ _36087_/CLK _32453_/D VGND VGND VPWR VPWR _32453_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_193_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17387_ _17067_/X _17385_/X _17386_/X _17071_/X VGND VGND VPWR VPWR _17387_/X sky130_fd_sc_hd__a22o_1
XFILLER_192_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31404_ _27819_/X _35919_/Q _31408_/S VGND VGND VPWR VPWR _31405_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19126_ _32107_/Q _32299_/Q _32363_/Q _35883_/Q _18874_/X _19015_/X VGND VGND VPWR
+ VPWR _19126_/X sky130_fd_sc_hd__mux4_1
X_16338_ _35165_/Q _35101_/Q _35037_/Q _32157_/Q _16304_/X _16305_/X VGND VGND VPWR
+ VPWR _16338_/X sky130_fd_sc_hd__mux4_1
XFILLER_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35172_ _35490_/CLK _35172_/D VGND VGND VPWR VPWR _35172_/Q sky130_fd_sc_hd__dfxtp_1
X_32384_ _35969_/CLK _32384_/D VGND VGND VPWR VPWR _32384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34123_ _34187_/CLK _34123_/D VGND VGND VPWR VPWR _34123_/Q sky130_fd_sc_hd__dfxtp_1
X_19057_ _18945_/X _19055_/X _19056_/X _18948_/X VGND VGND VPWR VPWR _19057_/X sky130_fd_sc_hd__a22o_1
X_31335_ _27717_/X _35886_/Q _31345_/S VGND VGND VPWR VPWR _31336_/A sky130_fd_sc_hd__mux2_1
X_16269_ _16078_/X _16267_/X _16268_/X _16088_/X VGND VGND VPWR VPWR _16269_/X sky130_fd_sc_hd__a22o_1
XFILLER_69_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18008_ _18008_/A VGND VGND VPWR VPWR _32012_/D sky130_fd_sc_hd__buf_2
X_34054_ _34182_/CLK _34054_/D VGND VGND VPWR VPWR _34054_/Q sky130_fd_sc_hd__dfxtp_1
X_31266_ _31266_/A VGND VGND VPWR VPWR _35853_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33005_ _36013_/CLK _33005_/D VGND VGND VPWR VPWR _33005_/Q sky130_fd_sc_hd__dfxtp_1
X_30217_ _30217_/A VGND VGND VPWR VPWR _35356_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31197_ _31197_/A VGND VGND VPWR VPWR _35820_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19959_ _33411_/Q _33347_/Q _33283_/Q _33219_/Q _19780_/X _19781_/X VGND VGND VPWR
+ VPWR _19959_/X sky130_fd_sc_hd__mux4_1
XFILLER_141_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30148_ _35324_/Q _29447_/X _30150_/S VGND VGND VPWR VPWR _30149_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34956_ _34956_/CLK _34956_/D VGND VGND VPWR VPWR _34956_/Q sky130_fd_sc_hd__dfxtp_1
X_22970_ _22970_/A VGND VGND VPWR VPWR _32048_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_228_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30079_ _35291_/Q _29345_/X _30087_/S VGND VGND VPWR VPWR _30080_/A sky130_fd_sc_hd__mux2_1
X_21921_ _21598_/X _21919_/X _21920_/X _21601_/X VGND VGND VPWR VPWR _21921_/X sky130_fd_sc_hd__a22o_1
XFILLER_83_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33907_ _36085_/CLK _33907_/D VGND VGND VPWR VPWR _33907_/Q sky130_fd_sc_hd__dfxtp_1
X_34887_ _36167_/CLK _34887_/D VGND VGND VPWR VPWR _34887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24640_ _24640_/A VGND VGND VPWR VPWR _32843_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33838_ _33902_/CLK _33838_/D VGND VGND VPWR VPWR _33838_/Q sky130_fd_sc_hd__dfxtp_1
X_21852_ _35639_/Q _34999_/Q _34359_/Q _33719_/Q _21744_/X _21745_/X VGND VGND VPWR
+ VPWR _21852_/X sky130_fd_sc_hd__mux4_1
XFILLER_167_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20803_ _20678_/X _20801_/X _20802_/X _20688_/X VGND VGND VPWR VPWR _20803_/X sky130_fd_sc_hd__a22o_1
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24571_ _24571_/A VGND VGND VPWR VPWR _32810_/D sky130_fd_sc_hd__clkbuf_1
X_33769_ _35624_/CLK _33769_/D VGND VGND VPWR VPWR _33769_/Q sky130_fd_sc_hd__dfxtp_1
X_21783_ _35701_/Q _32210_/Q _35573_/Q _35509_/Q _21564_/X _21565_/X VGND VGND VPWR
+ VPWR _21783_/X sky130_fd_sc_hd__mux4_1
XFILLER_58_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26310_ _26310_/A VGND VGND VPWR VPWR _33601_/D sky130_fd_sc_hd__clkbuf_1
X_23522_ _32256_/Q _23429_/X _23536_/S VGND VGND VPWR VPWR _23523_/A sky130_fd_sc_hd__mux2_1
X_20734_ _34391_/Q _36119_/Q _34263_/Q _34199_/Q _20692_/X _20694_/X VGND VGND VPWR
+ VPWR _20734_/X sky130_fd_sc_hd__mux4_1
X_27290_ _34032_/Q _27115_/X _27296_/S VGND VGND VPWR VPWR _27291_/A sky130_fd_sc_hd__mux2_1
X_35508_ _35699_/CLK _35508_/D VGND VGND VPWR VPWR _35508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26241_ _26241_/A VGND VGND VPWR VPWR _33568_/D sky130_fd_sc_hd__clkbuf_1
X_23453_ input46/X VGND VGND VPWR VPWR _23453_/X sky130_fd_sc_hd__buf_6
X_35439_ _35439_/CLK _35439_/D VGND VGND VPWR VPWR _35439_/Q sky130_fd_sc_hd__dfxtp_1
X_20665_ _35414_/Q _35350_/Q _35286_/Q _35222_/Q _20662_/X _20664_/X VGND VGND VPWR
+ VPWR _20665_/X sky130_fd_sc_hd__mux4_1
XFILLER_195_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_225_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1043 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22404_ _33927_/Q _33863_/Q _33799_/Q _36103_/Q _22330_/X _22331_/X VGND VGND VPWR
+ VPWR _22404_/X sky130_fd_sc_hd__mux4_1
XFILLER_195_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26172_ _24930_/X _33536_/Q _26186_/S VGND VGND VPWR VPWR _26173_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23384_ input22/X VGND VGND VPWR VPWR _23384_/X sky130_fd_sc_hd__buf_4
X_20596_ _34134_/Q _34070_/Q _34006_/Q _33942_/Q _20593_/X _20595_/X VGND VGND VPWR
+ VPWR _20596_/X sky130_fd_sc_hd__mux4_1
X_25123_ _25123_/A VGND VGND VPWR VPWR _33041_/D sky130_fd_sc_hd__clkbuf_1
X_22335_ _32645_/Q _32581_/Q _32517_/Q _35973_/Q _22229_/X _22013_/X VGND VGND VPWR
+ VPWR _22335_/X sky130_fd_sc_hd__mux4_1
XFILLER_100_1008 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29931_ _29931_/A VGND VGND VPWR VPWR _35221_/D sky130_fd_sc_hd__clkbuf_1
X_25054_ _25054_/A VGND VGND VPWR VPWR _33008_/D sky130_fd_sc_hd__clkbuf_1
X_22266_ _32131_/Q _32323_/Q _32387_/Q _35907_/Q _22233_/X _22021_/X VGND VGND VPWR
+ VPWR _22266_/X sky130_fd_sc_hd__mux4_1
XFILLER_219_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24005_ _22922_/X _32545_/Q _24021_/S VGND VGND VPWR VPWR _24006_/A sky130_fd_sc_hd__mux2_1
X_21217_ _33061_/Q _32037_/Q _35813_/Q _35749_/Q _20972_/X _20973_/X VGND VGND VPWR
+ VPWR _21217_/X sky130_fd_sc_hd__mux4_1
XFILLER_132_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29862_ _35188_/Q _29422_/X _29880_/S VGND VGND VPWR VPWR _29863_/A sky130_fd_sc_hd__mux2_1
X_22197_ _32641_/Q _32577_/Q _32513_/Q _35969_/Q _21876_/X _22013_/X VGND VGND VPWR
+ VPWR _22197_/X sky130_fd_sc_hd__mux4_1
XFILLER_105_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28813_ _34721_/Q _27069_/X _28829_/S VGND VGND VPWR VPWR _28814_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21148_ _22560_/A VGND VGND VPWR VPWR _21148_/X sky130_fd_sc_hd__buf_4
X_29793_ _35156_/Q _29521_/X _29795_/S VGND VGND VPWR VPWR _29794_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28744_ _28744_/A VGND VGND VPWR VPWR _34689_/D sky130_fd_sc_hd__clkbuf_1
X_25956_ _25956_/A VGND VGND VPWR VPWR _33433_/D sky130_fd_sc_hd__clkbuf_1
X_21079_ _20892_/X _21077_/X _21078_/X _20895_/X VGND VGND VPWR VPWR _21079_/X sky130_fd_sc_hd__a22o_1
XFILLER_24_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_247_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24907_ _24907_/A VGND VGND VPWR VPWR _32952_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28675_ _28675_/A VGND VGND VPWR VPWR _34656_/D sky130_fd_sc_hd__clkbuf_1
X_25887_ _24908_/X _33401_/Q _25895_/S VGND VGND VPWR VPWR _25888_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27626_ _27626_/A VGND VGND VPWR VPWR _34191_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24838_ _24837_/X _32930_/Q _24859_/S VGND VGND VPWR VPWR _24839_/A sky130_fd_sc_hd__mux2_1
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27557_ _27557_/A VGND VGND VPWR VPWR _34158_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24769_ _24769_/A VGND VGND VPWR VPWR _32904_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17310_ _32633_/Q _32569_/Q _32505_/Q _35961_/Q _17276_/X _17060_/X VGND VGND VPWR
+ VPWR _17310_/X sky130_fd_sc_hd__mux4_1
X_26508_ _26508_/A VGND VGND VPWR VPWR _33694_/D sky130_fd_sc_hd__clkbuf_1
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18290_ _20071_/A VGND VGND VPWR VPWR _20210_/A sky130_fd_sc_hd__buf_12
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27488_ _34126_/Q _27208_/X _27494_/S VGND VGND VPWR VPWR _27489_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_226_1279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17241_ _33911_/Q _33847_/Q _33783_/Q _36087_/Q _17024_/X _17025_/X VGND VGND VPWR
+ VPWR _17241_/X sky130_fd_sc_hd__mux4_1
X_29227_ _29227_/A VGND VGND VPWR VPWR _34917_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26439_ _33662_/Q _23420_/X _26457_/S VGND VGND VPWR VPWR _26440_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29158_ _34885_/Q _27180_/X _29162_/S VGND VGND VPWR VPWR _29159_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17172_ _33397_/Q _33333_/Q _33269_/Q _33205_/Q _17127_/X _17128_/X VGND VGND VPWR
+ VPWR _17172_/X sky130_fd_sc_hd__mux4_1
XFILLER_35_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16123_ _16119_/X _16122_/X _16044_/X _16046_/X VGND VGND VPWR VPWR _16138_/B sky130_fd_sc_hd__o211a_1
X_28109_ _28109_/A VGND VGND VPWR VPWR _34389_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29089_ _34852_/Q _27078_/X _29099_/S VGND VGND VPWR VPWR _29090_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31120_ _31120_/A VGND VGND VPWR VPWR _35784_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16054_ _17766_/A VGND VGND VPWR VPWR _17999_/A sky130_fd_sc_hd__buf_12
XFILLER_142_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1012 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31051_ _35752_/Q input10/X _31053_/S VGND VGND VPWR VPWR _31052_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19813_ _20166_/A VGND VGND VPWR VPWR _19813_/X sky130_fd_sc_hd__buf_4
XFILLER_123_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30002_ _30002_/A VGND VGND VPWR VPWR _35254_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34810_ _36153_/CLK _34810_/D VGND VGND VPWR VPWR _34810_/Q sky130_fd_sc_hd__dfxtp_1
X_19744_ _19744_/A VGND VGND VPWR VPWR _32444_/D sky130_fd_sc_hd__clkbuf_4
X_35790_ _35855_/CLK _35790_/D VGND VGND VPWR VPWR _35790_/Q sky130_fd_sc_hd__dfxtp_1
X_16956_ _16952_/X _16955_/X _16779_/X VGND VGND VPWR VPWR _16980_/A sky130_fd_sc_hd__o21ba_1
XFILLER_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34741_ _35126_/CLK _34741_/D VGND VGND VPWR VPWR _34741_/Q sky130_fd_sc_hd__dfxtp_1
X_31953_ _31953_/A VGND VGND VPWR VPWR _36179_/D sky130_fd_sc_hd__clkbuf_1
X_19675_ _19499_/X _19673_/X _19674_/X _19504_/X VGND VGND VPWR VPWR _19675_/X sky130_fd_sc_hd__a22o_1
X_16887_ _33389_/Q _33325_/Q _33261_/Q _33197_/Q _16774_/X _16775_/X VGND VGND VPWR
+ VPWR _16887_/X sky130_fd_sc_hd__mux4_1
XFILLER_225_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18626_ _32093_/Q _32285_/Q _32349_/Q _35869_/Q _18521_/X _20167_/A VGND VGND VPWR
+ VPWR _18626_/X sky130_fd_sc_hd__mux4_1
X_30904_ _35682_/Q input4/X _30918_/S VGND VGND VPWR VPWR _30905_/A sky130_fd_sc_hd__mux2_1
XTAP_4190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34672_ _34927_/CLK _34672_/D VGND VGND VPWR VPWR _34672_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31884_ _31884_/A VGND VGND VPWR VPWR _36146_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_225_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33623_ _35995_/CLK _33623_/D VGND VGND VPWR VPWR _33623_/Q sky130_fd_sc_hd__dfxtp_1
X_18557_ _18553_/X _18556_/X _18344_/X _18346_/X VGND VGND VPWR VPWR _18574_/B sky130_fd_sc_hd__o211a_1
X_30835_ _30835_/A VGND VGND VPWR VPWR _35649_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17508_ _35198_/Q _35134_/Q _35070_/Q _32254_/Q _17363_/X _17364_/X VGND VGND VPWR
+ VPWR _17508_/X sky130_fd_sc_hd__mux4_1
XFILLER_33_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33554_ _33875_/CLK _33554_/D VGND VGND VPWR VPWR _33554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18488_ _32089_/Q _32281_/Q _32345_/Q _35865_/Q _18332_/X _20167_/A VGND VGND VPWR
+ VPWR _18488_/X sky130_fd_sc_hd__mux4_1
XFILLER_36_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30766_ _30766_/A VGND VGND VPWR VPWR _35616_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32505_ _36025_/CLK _32505_/D VGND VGND VPWR VPWR _32505_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17439_ _34428_/Q _36156_/Q _34300_/Q _34236_/Q _17229_/X _17230_/X VGND VGND VPWR
+ VPWR _17439_/X sky130_fd_sc_hd__mux4_1
X_33485_ _34441_/CLK _33485_/D VGND VGND VPWR VPWR _33485_/Q sky130_fd_sc_hd__dfxtp_1
X_30697_ _35584_/Q _29460_/X _30711_/S VGND VGND VPWR VPWR _30698_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35224_ _35799_/CLK _35224_/D VGND VGND VPWR VPWR _35224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20450_ _34705_/Q _34641_/Q _34577_/Q _34513_/Q _20298_/X _20299_/X VGND VGND VPWR
+ VPWR _20450_/X sky130_fd_sc_hd__mux4_1
XFILLER_165_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32436_ _33895_/CLK _32436_/D VGND VGND VPWR VPWR _32436_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19109_ _34922_/Q _34858_/Q _34794_/Q _34730_/Q _19107_/X _19108_/X VGND VGND VPWR
+ VPWR _19109_/X sky130_fd_sc_hd__mux4_1
XFILLER_101_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35155_ _36114_/CLK _35155_/D VGND VGND VPWR VPWR _35155_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20381_ _20073_/X _20379_/X _20380_/X _20077_/X VGND VGND VPWR VPWR _20381_/X sky130_fd_sc_hd__a22o_1
X_32367_ _32877_/CLK _32367_/D VGND VGND VPWR VPWR _32367_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22120_ _22120_/A _22120_/B _22120_/C _22120_/D VGND VGND VPWR VPWR _22121_/A sky130_fd_sc_hd__or4_4
X_34106_ _35320_/CLK _34106_/D VGND VGND VPWR VPWR _34106_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31318_ _27692_/X _35878_/Q _31324_/S VGND VGND VPWR VPWR _31319_/A sky130_fd_sc_hd__mux2_1
X_35086_ _35731_/CLK _35086_/D VGND VGND VPWR VPWR _35086_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput110 _31986_/Q VGND VGND VPWR VPWR D1[28] sky130_fd_sc_hd__buf_2
X_32298_ _35949_/CLK _32298_/D VGND VGND VPWR VPWR _32298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput121 _31996_/Q VGND VGND VPWR VPWR D1[38] sky130_fd_sc_hd__buf_2
Xoutput132 _32006_/Q VGND VGND VPWR VPWR D1[48] sky130_fd_sc_hd__buf_2
Xoutput143 _32016_/Q VGND VGND VPWR VPWR D1[58] sky130_fd_sc_hd__buf_2
X_34037_ _34101_/CLK _34037_/D VGND VGND VPWR VPWR _34037_/Q sky130_fd_sc_hd__dfxtp_1
X_22051_ _33917_/Q _33853_/Q _33789_/Q _36093_/Q _21977_/X _21978_/X VGND VGND VPWR
+ VPWR _22051_/X sky130_fd_sc_hd__mux4_1
XTAP_6509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31249_ _31249_/A VGND VGND VPWR VPWR _35845_/D sky130_fd_sc_hd__clkbuf_1
Xoutput154 _36182_/Q VGND VGND VPWR VPWR D2[0] sky130_fd_sc_hd__buf_2
XFILLER_82_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput165 _36183_/Q VGND VGND VPWR VPWR D2[1] sky130_fd_sc_hd__buf_2
XFILLER_115_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput176 _36184_/Q VGND VGND VPWR VPWR D2[2] sky130_fd_sc_hd__buf_2
XFILLER_130_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21002_ _35679_/Q _32185_/Q _35551_/Q _35487_/Q _20858_/X _20859_/X VGND VGND VPWR
+ VPWR _21002_/X sky130_fd_sc_hd__mux4_1
XFILLER_114_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput187 _36185_/Q VGND VGND VPWR VPWR D2[3] sky130_fd_sc_hd__buf_2
XFILLER_248_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput198 _36186_/Q VGND VGND VPWR VPWR D2[4] sky130_fd_sc_hd__buf_2
XTAP_5819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_955 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25810_ _24994_/X _33365_/Q _25810_/S VGND VGND VPWR VPWR _25811_/A sky130_fd_sc_hd__mux2_1
X_26790_ _33826_/Q _23268_/X _26804_/S VGND VGND VPWR VPWR _26791_/A sky130_fd_sc_hd__mux2_1
X_35988_ _35988_/CLK _35988_/D VGND VGND VPWR VPWR _35988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25741_ _25810_/S VGND VGND VPWR VPWR _25760_/S sky130_fd_sc_hd__buf_4
X_22953_ input14/X VGND VGND VPWR VPWR _22953_/X sky130_fd_sc_hd__buf_2
XFILLER_228_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34939_ _34941_/CLK _34939_/D VGND VGND VPWR VPWR _34939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_244_834 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21904_ _34169_/Q _34105_/Q _34041_/Q _33977_/Q _21693_/X _21694_/X VGND VGND VPWR
+ VPWR _21904_/X sky130_fd_sc_hd__mux4_1
XFILLER_28_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_906 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28460_ _28460_/A VGND VGND VPWR VPWR _34555_/D sky130_fd_sc_hd__clkbuf_1
X_25672_ _25672_/A VGND VGND VPWR VPWR _33299_/D sky130_fd_sc_hd__clkbuf_1
X_22884_ _25132_/A _28786_/A input85/X VGND VGND VPWR VPWR _22885_/A sky130_fd_sc_hd__or3b_1
X_27411_ _27411_/A VGND VGND VPWR VPWR _34089_/D sky130_fd_sc_hd__clkbuf_1
X_24623_ _24623_/A VGND VGND VPWR VPWR _32835_/D sky130_fd_sc_hd__clkbuf_1
X_21835_ _21835_/A _21835_/B _21835_/C _21835_/D VGND VGND VPWR VPWR _21836_/A sky130_fd_sc_hd__or4_1
X_28391_ _28391_/A VGND VGND VPWR VPWR _34522_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27342_ _27342_/A VGND VGND VPWR VPWR _34056_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24554_ _24554_/A VGND VGND VPWR VPWR _32802_/D sky130_fd_sc_hd__clkbuf_1
X_21766_ _21757_/X _21764_/X _21765_/X VGND VGND VPWR VPWR _21767_/D sky130_fd_sc_hd__o21ba_1
XFILLER_93_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20717_ _32599_/Q _32535_/Q _32471_/Q _35927_/Q _22466_/A _22317_/A VGND VGND VPWR
+ VPWR _20717_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_1266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23505_ _32248_/Q _23402_/X _23515_/S VGND VGND VPWR VPWR _23506_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24485_ _23024_/X _32770_/Q _24495_/S VGND VGND VPWR VPWR _24486_/A sky130_fd_sc_hd__mux2_1
X_27273_ _34024_/Q _27090_/X _27275_/S VGND VGND VPWR VPWR _27274_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21697_ _33395_/Q _33331_/Q _33267_/Q _33203_/Q _21374_/X _21375_/X VGND VGND VPWR
+ VPWR _21697_/X sky130_fd_sc_hd__mux4_1
XFILLER_106_1239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29012_ _29012_/A VGND VGND VPWR VPWR _34815_/D sky130_fd_sc_hd__clkbuf_1
X_26224_ _26224_/A VGND VGND VPWR VPWR _33560_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23436_ _32224_/Q _23435_/X _23451_/S VGND VGND VPWR VPWR _23437_/A sky130_fd_sc_hd__mux2_1
X_20648_ _22459_/A VGND VGND VPWR VPWR _20648_/X sky130_fd_sc_hd__buf_4
XFILLER_109_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26155_ _24905_/X _33528_/Q _26165_/S VGND VGND VPWR VPWR _26156_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_192_CLK clkbuf_6_48__f_CLK/X VGND VGND VPWR VPWR _36044_/CLK sky130_fd_sc_hd__clkbuf_16
X_23367_ _32199_/Q _23296_/X _23385_/S VGND VGND VPWR VPWR _23368_/A sky130_fd_sc_hd__mux2_1
X_20579_ input73/X input74/X VGND VGND VPWR VPWR _22365_/A sky130_fd_sc_hd__nor2b_4
XFILLER_180_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22318_ _35204_/Q _35140_/Q _35076_/Q _32260_/Q _22316_/X _22317_/X VGND VGND VPWR
+ VPWR _22318_/X sky130_fd_sc_hd__mux4_1
XFILLER_164_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25106_ _24958_/X _33033_/Q _25122_/S VGND VGND VPWR VPWR _25107_/A sky130_fd_sc_hd__mux2_1
X_26086_ _24803_/X _33495_/Q _26102_/S VGND VGND VPWR VPWR _26087_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_1182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23298_ _23298_/A VGND VGND VPWR VPWR _32171_/D sky130_fd_sc_hd__clkbuf_1
X_29914_ _35213_/Q _29500_/X _29922_/S VGND VGND VPWR VPWR _29915_/A sky130_fd_sc_hd__mux2_1
X_25037_ _25037_/A VGND VGND VPWR VPWR _33000_/D sky130_fd_sc_hd__clkbuf_1
X_22249_ _22106_/X _22247_/X _22248_/X _22109_/X VGND VGND VPWR VPWR _22249_/X sky130_fd_sc_hd__a22o_1
XFILLER_106_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29845_ _35180_/Q _29398_/X _29859_/S VGND VGND VPWR VPWR _29846_/A sky130_fd_sc_hd__mux2_1
XFILLER_239_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16810_ _17163_/A VGND VGND VPWR VPWR _16810_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_94_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29776_ _29776_/A VGND VGND VPWR VPWR _35147_/D sky130_fd_sc_hd__clkbuf_1
X_17790_ _35206_/Q _35142_/Q _35078_/Q _32262_/Q _17716_/X _17717_/X VGND VGND VPWR
+ VPWR _17790_/X sky130_fd_sc_hd__mux4_1
XFILLER_232_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26988_ _33920_/Q _23429_/X _27002_/S VGND VGND VPWR VPWR _26989_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16741_ _17961_/A VGND VGND VPWR VPWR _16741_/X sky130_fd_sc_hd__buf_4
X_28727_ _28727_/A VGND VGND VPWR VPWR _34681_/D sky130_fd_sc_hd__clkbuf_1
X_25939_ _24985_/X _33426_/Q _25945_/S VGND VGND VPWR VPWR _25940_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19460_ _20166_/A VGND VGND VPWR VPWR _19460_/X sky130_fd_sc_hd__buf_4
X_28658_ _28658_/A VGND VGND VPWR VPWR _34648_/D sky130_fd_sc_hd__clkbuf_1
X_16672_ _17851_/A VGND VGND VPWR VPWR _16672_/X sky130_fd_sc_hd__buf_4
XFILLER_46_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_6_25__f_CLK clkbuf_5_12_0_CLK/X VGND VGND VPWR VPWR clkbuf_leaf_77_CLK/A sky130_fd_sc_hd__clkbuf_16
XFILLER_98_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18411_ _33367_/Q _33303_/Q _33239_/Q _33175_/Q _18302_/X _18303_/X VGND VGND VPWR
+ VPWR _18411_/X sky130_fd_sc_hd__mux4_1
XFILLER_62_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27609_ _27609_/A VGND VGND VPWR VPWR _34183_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19391_ _19391_/A VGND VGND VPWR VPWR _32434_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28589_ _28589_/A VGND VGND VPWR VPWR _34616_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18342_ _18330_/X _18335_/X _18340_/X _18341_/X VGND VGND VPWR VPWR _18342_/X sky130_fd_sc_hd__a22o_1
X_30620_ _30620_/A VGND VGND VPWR VPWR _35547_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18273_ _34453_/Q _36181_/Q _34325_/Q _34261_/Q _16067_/X _16069_/X VGND VGND VPWR
+ VPWR _18273_/X sky130_fd_sc_hd__mux4_1
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30551_ _35515_/Q _29444_/X _30555_/S VGND VGND VPWR VPWR _30552_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17224_ _17003_/X _17222_/X _17223_/X _17006_/X VGND VGND VPWR VPWR _17224_/X sky130_fd_sc_hd__a22o_1
X_33270_ _36087_/CLK _33270_/D VGND VGND VPWR VPWR _33270_/Q sky130_fd_sc_hd__dfxtp_1
X_30482_ _35482_/Q _29342_/X _30492_/S VGND VGND VPWR VPWR _30483_/A sky130_fd_sc_hd__mux2_1
XFILLER_198_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput12 DW[1] VGND VGND VPWR VPWR input12/X sky130_fd_sc_hd__buf_8
Xinput23 DW[2] VGND VGND VPWR VPWR input23/X sky130_fd_sc_hd__clkbuf_16
XFILLER_204_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32221_ _35711_/CLK _32221_/D VGND VGND VPWR VPWR _32221_/Q sky130_fd_sc_hd__dfxtp_1
Xinput34 DW[3] VGND VGND VPWR VPWR input34/X sky130_fd_sc_hd__buf_8
Xinput45 DW[4] VGND VGND VPWR VPWR input45/X sky130_fd_sc_hd__buf_8
X_17155_ _35188_/Q _35124_/Q _35060_/Q _32231_/Q _17010_/X _17011_/X VGND VGND VPWR
+ VPWR _17155_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_183_CLK clkbuf_6_27__f_CLK/X VGND VGND VPWR VPWR _35857_/CLK sky130_fd_sc_hd__clkbuf_16
Xinput56 DW[5] VGND VGND VPWR VPWR input56/X sky130_fd_sc_hd__buf_8
Xinput67 R1[2] VGND VGND VPWR VPWR input67/X sky130_fd_sc_hd__buf_6
XFILLER_239_1426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput78 R3[1] VGND VGND VPWR VPWR input78/X sky130_fd_sc_hd__clkbuf_1
X_16106_ _16106_/A _16106_/B _16106_/C _16106_/D VGND VGND VPWR VPWR _16107_/A sky130_fd_sc_hd__or4_2
XFILLER_128_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput89 WE VGND VGND VPWR VPWR input89/X sky130_fd_sc_hd__buf_6
XFILLER_239_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32152_ _35162_/CLK _32152_/D VGND VGND VPWR VPWR _32152_/Q sky130_fd_sc_hd__dfxtp_1
X_17086_ _34418_/Q _36146_/Q _34290_/Q _34226_/Q _16876_/X _16877_/X VGND VGND VPWR
+ VPWR _17086_/X sky130_fd_sc_hd__mux4_1
XFILLER_48_1410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31103_ _31103_/A VGND VGND VPWR VPWR _35776_/D sky130_fd_sc_hd__clkbuf_1
X_16037_ _17833_/A VGND VGND VPWR VPWR _16037_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_170_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32083_ _35859_/CLK _32083_/D VGND VGND VPWR VPWR _32083_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35911_ _35974_/CLK _35911_/D VGND VGND VPWR VPWR _35911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31034_ _31145_/S VGND VGND VPWR VPWR _31053_/S sky130_fd_sc_hd__buf_4
XFILLER_170_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35842_ _36034_/CLK _35842_/D VGND VGND VPWR VPWR _35842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17988_ _32908_/Q _32844_/Q _32780_/Q _32716_/Q _17699_/X _17700_/X VGND VGND VPWR
+ VPWR _17988_/X sky130_fd_sc_hd__mux4_1
XFILLER_211_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19727_ _35708_/Q _32217_/Q _35580_/Q _35516_/Q _19617_/X _19618_/X VGND VGND VPWR
+ VPWR _19727_/X sky130_fd_sc_hd__mux4_1
XFILLER_211_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16939_ _17998_/A VGND VGND VPWR VPWR _16939_/X sky130_fd_sc_hd__buf_6
X_32985_ _34135_/CLK _32985_/D VGND VGND VPWR VPWR _32985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35773_ _36029_/CLK _35773_/D VGND VGND VPWR VPWR _35773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31936_ _23466_/X _36171_/Q _31948_/S VGND VGND VPWR VPWR _31937_/A sky130_fd_sc_hd__mux2_1
X_34724_ _34918_/CLK _34724_/D VGND VGND VPWR VPWR _34724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19658_ _33082_/Q _32058_/Q _35834_/Q _35770_/Q _19378_/X _19379_/X VGND VGND VPWR
+ VPWR _19658_/X sky130_fd_sc_hd__mux4_1
XFILLER_237_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18609_ _34908_/Q _34844_/Q _34780_/Q _34716_/Q _18396_/X _18398_/X VGND VGND VPWR
+ VPWR _18609_/X sky130_fd_sc_hd__mux4_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34655_ _35544_/CLK _34655_/D VGND VGND VPWR VPWR _34655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19589_ _33080_/Q _32056_/Q _35832_/Q _35768_/Q _19378_/X _19379_/X VGND VGND VPWR
+ VPWR _19589_/X sky130_fd_sc_hd__mux4_1
X_31867_ _23292_/X _36138_/Q _31885_/S VGND VGND VPWR VPWR _31868_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_1299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33606_ _34179_/CLK _33606_/D VGND VGND VPWR VPWR _33606_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21620_ _33649_/Q _33585_/Q _33521_/Q _33457_/Q _21447_/X _21448_/X VGND VGND VPWR
+ VPWR _21620_/X sky130_fd_sc_hd__mux4_1
X_30818_ _30818_/A VGND VGND VPWR VPWR _35641_/D sky130_fd_sc_hd__clkbuf_1
X_34586_ _35544_/CLK _34586_/D VGND VGND VPWR VPWR _34586_/Q sky130_fd_sc_hd__dfxtp_1
X_31798_ _31798_/A VGND VGND VPWR VPWR _36105_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33537_ _33984_/CLK _33537_/D VGND VGND VPWR VPWR _33537_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21551_ _34159_/Q _34095_/Q _34031_/Q _33967_/Q _21340_/X _21341_/X VGND VGND VPWR
+ VPWR _21551_/X sky130_fd_sc_hd__mux4_1
XFILLER_55_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30749_ _30749_/A VGND VGND VPWR VPWR _35608_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20502_ _20498_/X _20501_/X _20146_/A _20147_/A VGND VGND VPWR VPWR _20517_/B sky130_fd_sc_hd__o211a_1
XFILLER_222_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24270_ _22906_/X _32668_/Q _24276_/S VGND VGND VPWR VPWR _24271_/A sky130_fd_sc_hd__mux2_1
X_33468_ _36093_/CLK _33468_/D VGND VGND VPWR VPWR _33468_/Q sky130_fd_sc_hd__dfxtp_1
X_21482_ _21482_/A _21482_/B _21482_/C _21482_/D VGND VGND VPWR VPWR _21483_/A sky130_fd_sc_hd__or4_4
XFILLER_140_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35207_ _35718_/CLK _35207_/D VGND VGND VPWR VPWR _35207_/Q sky130_fd_sc_hd__dfxtp_1
X_23221_ _23079_/X _32148_/Q _23223_/S VGND VGND VPWR VPWR _23222_/A sky130_fd_sc_hd__mux2_1
XFILLER_222_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20433_ _33937_/Q _33873_/Q _33809_/Q _36113_/Q _18362_/X _18364_/X VGND VGND VPWR
+ VPWR _20433_/X sky130_fd_sc_hd__mux4_1
X_32419_ _33828_/CLK _32419_/D VGND VGND VPWR VPWR _32419_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_174_CLK clkbuf_leaf_77_CLK/A VGND VGND VPWR VPWR _35669_/CLK sky130_fd_sc_hd__clkbuf_16
X_36187_ _36191_/CLK _36187_/D VGND VGND VPWR VPWR _36187_/Q sky130_fd_sc_hd__dfxtp_1
X_33399_ _33911_/CLK _33399_/D VGND VGND VPWR VPWR _33399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35138_ _35655_/CLK _35138_/D VGND VGND VPWR VPWR _35138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23152_ _22977_/X _32115_/Q _23152_/S VGND VGND VPWR VPWR _23153_/A sky130_fd_sc_hd__mux2_1
X_20364_ _34958_/Q _34894_/Q _34830_/Q _34766_/Q _20166_/X _20167_/X VGND VGND VPWR
+ VPWR _20364_/X sky130_fd_sc_hd__mux4_1
XTAP_7007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22103_ _21956_/X _22101_/X _22102_/X _21959_/X VGND VGND VPWR VPWR _22103_/X sky130_fd_sc_hd__a22o_1
XTAP_7029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27960_ _27960_/A VGND VGND VPWR VPWR _34318_/D sky130_fd_sc_hd__clkbuf_1
X_23083_ _23082_/X _32085_/Q _23083_/S VGND VGND VPWR VPWR _23084_/A sky130_fd_sc_hd__mux2_1
X_35069_ _35577_/CLK _35069_/D VGND VGND VPWR VPWR _35069_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20295_ _33100_/Q _32076_/Q _35852_/Q _35788_/Q _20084_/X _20085_/X VGND VGND VPWR
+ VPWR _20295_/X sky130_fd_sc_hd__mux4_1
XTAP_6317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26911_ _26911_/A VGND VGND VPWR VPWR _33883_/D sky130_fd_sc_hd__clkbuf_1
X_22034_ _21956_/X _22030_/X _22033_/X _21959_/X VGND VGND VPWR VPWR _22034_/X sky130_fd_sc_hd__a22o_1
XTAP_6339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27891_ _27891_/A VGND VGND VPWR VPWR _34285_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29630_ _29630_/A VGND VGND VPWR VPWR _35078_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26842_ _33851_/Q _23411_/X _26846_/S VGND VGND VPWR VPWR _26843_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29561_ _29561_/A VGND VGND VPWR VPWR _35045_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26773_ _33818_/Q _23243_/X _26783_/S VGND VGND VPWR VPWR _26774_/A sky130_fd_sc_hd__mux2_1
X_23985_ _23985_/A VGND VGND VPWR VPWR _32535_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28512_ _28512_/A VGND VGND VPWR VPWR _34580_/D sky130_fd_sc_hd__clkbuf_1
X_25724_ _25724_/A VGND VGND VPWR VPWR _33323_/D sky130_fd_sc_hd__clkbuf_1
X_29492_ _35018_/Q _29491_/X _29513_/S VGND VGND VPWR VPWR _29493_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22936_ _22936_/A VGND VGND VPWR VPWR _32037_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_1333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28443_ _28443_/A VGND VGND VPWR VPWR _34547_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25655_ _24964_/X _33291_/Q _25667_/S VGND VGND VPWR VPWR _25656_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22867_ _33109_/Q _32085_/Q _35861_/Q _35797_/Q _20679_/X _20680_/X VGND VGND VPWR
+ VPWR _22867_/X sky130_fd_sc_hd__mux4_1
XFILLER_73_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24606_ _24606_/A VGND VGND VPWR VPWR _32827_/D sky130_fd_sc_hd__clkbuf_1
X_28374_ _27831_/X _34515_/Q _28378_/S VGND VGND VPWR VPWR _28375_/A sky130_fd_sc_hd__mux2_1
XPHY_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21818_ _21814_/X _21817_/X _21740_/X _21741_/X VGND VGND VPWR VPWR _21835_/B sky130_fd_sc_hd__o211a_1
XPHY_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22798_ _21753_/A _22796_/X _22797_/X _21756_/A VGND VGND VPWR VPWR _22798_/X sky130_fd_sc_hd__a22o_1
X_25586_ _24861_/X _33258_/Q _25604_/S VGND VGND VPWR VPWR _25587_/A sky130_fd_sc_hd__mux2_1
XPHY_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27325_ _27325_/A VGND VGND VPWR VPWR _34048_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24537_ _24537_/A VGND VGND VPWR VPWR _32794_/D sky130_fd_sc_hd__clkbuf_1
X_21749_ _33076_/Q _32052_/Q _35828_/Q _35764_/Q _21678_/X _21679_/X VGND VGND VPWR
+ VPWR _21749_/X sky130_fd_sc_hd__mux4_1
XPHY_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_964 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_936 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27256_ _27367_/S VGND VGND VPWR VPWR _27275_/S sky130_fd_sc_hd__buf_6
XFILLER_71_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_1058 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24468_ _22999_/X _32762_/Q _24474_/S VGND VGND VPWR VPWR _24469_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26207_ _24982_/X _33553_/Q _26207_/S VGND VGND VPWR VPWR _26208_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_165_CLK clkbuf_6_30__f_CLK/X VGND VGND VPWR VPWR _35728_/CLK sky130_fd_sc_hd__clkbuf_16
X_23419_ _23419_/A VGND VGND VPWR VPWR _32218_/D sky130_fd_sc_hd__clkbuf_1
X_27187_ _33991_/Q _27186_/X _27187_/S VGND VGND VPWR VPWR _27188_/A sky130_fd_sc_hd__mux2_1
X_24399_ _22897_/X _32729_/Q _24411_/S VGND VGND VPWR VPWR _24400_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26138_ _24880_/X _33520_/Q _26144_/S VGND VGND VPWR VPWR _26139_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_1326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18960_ _18747_/X _18956_/X _18959_/X _18750_/X VGND VGND VPWR VPWR _18960_/X sky130_fd_sc_hd__a22o_1
X_26069_ _26069_/A VGND VGND VPWR VPWR _33487_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17911_ _17905_/X _17908_/X _17909_/X _17910_/X VGND VGND VPWR VPWR _17911_/X sky130_fd_sc_hd__a22o_1
X_18891_ _34404_/Q _36132_/Q _34276_/Q _34212_/Q _18823_/X _18824_/X VGND VGND VPWR
+ VPWR _18891_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17842_ _17765_/X _17840_/X _17841_/X _17771_/X VGND VGND VPWR VPWR _17842_/X sky130_fd_sc_hd__a22o_1
X_29828_ _35172_/Q _29373_/X _29838_/S VGND VGND VPWR VPWR _29829_/A sky130_fd_sc_hd__mux2_1
XTAP_6873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29759_ _29759_/A VGND VGND VPWR VPWR _35139_/D sky130_fd_sc_hd__clkbuf_1
X_17773_ _17773_/A VGND VGND VPWR VPWR _17773_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_14_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19512_ _32630_/Q _32566_/Q _32502_/Q _35958_/Q _19223_/X _19360_/X VGND VGND VPWR
+ VPWR _19512_/X sky130_fd_sc_hd__mux4_1
X_16724_ _35432_/Q _35368_/Q _35304_/Q _35240_/Q _16548_/X _16549_/X VGND VGND VPWR
+ VPWR _16724_/X sky130_fd_sc_hd__mux4_1
X_32770_ _32894_/CLK _32770_/D VGND VGND VPWR VPWR _32770_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31721_ _36069_/Q input7/X _31729_/S VGND VGND VPWR VPWR _31722_/A sky130_fd_sc_hd__mux2_1
X_19443_ _35700_/Q _32208_/Q _35572_/Q _35508_/Q _19264_/X _19265_/X VGND VGND VPWR
+ VPWR _19443_/X sky130_fd_sc_hd__mux4_1
XFILLER_222_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16655_ _16649_/X _16654_/X _16445_/X VGND VGND VPWR VPWR _16665_/C sky130_fd_sc_hd__o21ba_1
XFILLER_62_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34440_ _34440_/CLK _34440_/D VGND VGND VPWR VPWR _34440_/Q sky130_fd_sc_hd__dfxtp_1
X_31652_ _31652_/A VGND VGND VPWR VPWR _36036_/D sky130_fd_sc_hd__clkbuf_1
X_19374_ _35698_/Q _32206_/Q _35570_/Q _35506_/Q _19264_/X _19265_/X VGND VGND VPWR
+ VPWR _19374_/X sky130_fd_sc_hd__mux4_1
XFILLER_222_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16586_ _17998_/A VGND VGND VPWR VPWR _16586_/X sky130_fd_sc_hd__buf_6
XFILLER_72_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_1463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18325_ _20207_/A VGND VGND VPWR VPWR _18325_/X sky130_fd_sc_hd__buf_4
X_30603_ _35540_/Q _29521_/X _30605_/S VGND VGND VPWR VPWR _30604_/A sky130_fd_sc_hd__mux2_1
XFILLER_188_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34371_ _35716_/CLK _34371_/D VGND VGND VPWR VPWR _34371_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_774 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31583_ _31583_/A VGND VGND VPWR VPWR _36003_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36110_ _36167_/CLK _36110_/D VGND VGND VPWR VPWR _36110_/Q sky130_fd_sc_hd__dfxtp_1
X_33322_ _36076_/CLK _33322_/D VGND VGND VPWR VPWR _33322_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18256_ _32661_/Q _32597_/Q _32533_/Q _35989_/Q _17982_/X _16877_/A VGND VGND VPWR
+ VPWR _18256_/X sky130_fd_sc_hd__mux4_1
XFILLER_124_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30534_ _35507_/Q _29419_/X _30534_/S VGND VGND VPWR VPWR _30535_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36041_ _36044_/CLK _36041_/D VGND VGND VPWR VPWR _36041_/Q sky130_fd_sc_hd__dfxtp_1
X_17207_ _33398_/Q _33334_/Q _33270_/Q _33206_/Q _17127_/X _17128_/X VGND VGND VPWR
+ VPWR _17207_/X sky130_fd_sc_hd__mux4_1
X_33253_ _36068_/CLK _33253_/D VGND VGND VPWR VPWR _33253_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_156_CLK clkbuf_6_31__f_CLK/X VGND VGND VPWR VPWR _34897_/CLK sky130_fd_sc_hd__clkbuf_16
X_18187_ _18187_/A _18187_/B _18187_/C _18187_/D VGND VGND VPWR VPWR _18188_/A sky130_fd_sc_hd__or4_4
X_30465_ _30465_/A VGND VGND VPWR VPWR _35474_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_239_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32204_ _35697_/CLK _32204_/D VGND VGND VPWR VPWR _32204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17138_ _32884_/Q _32820_/Q _32756_/Q _32692_/Q _16993_/X _16994_/X VGND VGND VPWR
+ VPWR _17138_/X sky130_fd_sc_hd__mux4_1
X_33184_ _36065_/CLK _33184_/D VGND VGND VPWR VPWR _33184_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30396_ _30396_/A VGND VGND VPWR VPWR _35441_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32135_ _35974_/CLK _32135_/D VGND VGND VPWR VPWR _32135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17069_ _32114_/Q _32306_/Q _32370_/Q _35890_/Q _16927_/X _17068_/X VGND VGND VPWR
+ VPWR _17069_/X sky130_fd_sc_hd__mux4_1
XFILLER_83_1142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20080_ _35718_/Q _32228_/Q _35590_/Q _35526_/Q _19970_/X _19971_/X VGND VGND VPWR
+ VPWR _20080_/X sky130_fd_sc_hd__mux4_1
XFILLER_170_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32066_ _36034_/CLK _32066_/D VGND VGND VPWR VPWR _32066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31017_ _31017_/A VGND VGND VPWR VPWR _35735_/D sky130_fd_sc_hd__clkbuf_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35825_ _36147_/CLK _35825_/D VGND VGND VPWR VPWR _35825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23770_ _23770_/A VGND VGND VPWR VPWR _32371_/D sky130_fd_sc_hd__clkbuf_1
X_20982_ _20691_/X _20980_/X _20981_/X _20701_/X VGND VGND VPWR VPWR _20982_/X sky130_fd_sc_hd__a22o_1
X_32968_ _36040_/CLK _32968_/D VGND VGND VPWR VPWR _32968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35756_ _35820_/CLK _35756_/D VGND VGND VPWR VPWR _35756_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22721_ _35216_/Q _35152_/Q _35088_/Q _32272_/Q _20692_/X _20694_/X VGND VGND VPWR
+ VPWR _22721_/X sky130_fd_sc_hd__mux4_1
X_34707_ _36114_/CLK _34707_/D VGND VGND VPWR VPWR _34707_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_246_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31919_ _23438_/X _36163_/Q _31927_/S VGND VGND VPWR VPWR _31920_/A sky130_fd_sc_hd__mux2_1
XFILLER_198_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32899_ _35907_/CLK _32899_/D VGND VGND VPWR VPWR _32899_/Q sky130_fd_sc_hd__dfxtp_1
X_35687_ _35687_/CLK _35687_/D VGND VGND VPWR VPWR _35687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_875 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22652_ _22648_/X _22651_/X _22446_/X _22447_/X VGND VGND VPWR VPWR _22667_/B sky130_fd_sc_hd__o211a_2
X_25440_ _24846_/X _33189_/Q _25448_/S VGND VGND VPWR VPWR _25441_/A sky130_fd_sc_hd__mux2_1
X_34638_ _35664_/CLK _34638_/D VGND VGND VPWR VPWR _34638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21603_ _22464_/A VGND VGND VPWR VPWR _21603_/X sky130_fd_sc_hd__buf_4
XFILLER_167_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34569_ _35208_/CLK _34569_/D VGND VGND VPWR VPWR _34569_/Q sky130_fd_sc_hd__dfxtp_1
X_25371_ _25371_/A VGND VGND VPWR VPWR _33157_/D sky130_fd_sc_hd__clkbuf_1
X_22583_ _32652_/Q _32588_/Q _32524_/Q _35980_/Q _22582_/X _22366_/X VGND VGND VPWR
+ VPWR _22583_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_395_CLK clkbuf_6_41__f_CLK/X VGND VGND VPWR VPWR _35768_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_240_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27110_ _33966_/Q _27109_/X _27125_/S VGND VGND VPWR VPWR _27111_/A sky130_fd_sc_hd__mux2_1
X_21534_ _21245_/X _21532_/X _21533_/X _21248_/X VGND VGND VPWR VPWR _21534_/X sky130_fd_sc_hd__a22o_1
X_24322_ _24322_/A VGND VGND VPWR VPWR _32692_/D sky130_fd_sc_hd__clkbuf_1
X_28090_ _34380_/Q _27202_/X _28100_/S VGND VGND VPWR VPWR _28091_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27041_ input23/X VGND VGND VPWR VPWR _27041_/X sky130_fd_sc_hd__clkbuf_4
X_24253_ input86/X input87/X input88/X VGND VGND VPWR VPWR _24254_/A sky130_fd_sc_hd__and3b_1
X_36239_ _36242_/CLK _36239_/D VGND VGND VPWR VPWR _36239_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_147_CLK clkbuf_6_29__f_CLK/X VGND VGND VPWR VPWR _36119_/CLK sky130_fd_sc_hd__clkbuf_16
X_21465_ _21461_/X _21464_/X _21387_/X _21388_/X VGND VGND VPWR VPWR _21482_/B sky130_fd_sc_hd__o211a_1
XFILLER_119_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23204_ _23204_/A VGND VGND VPWR VPWR _32139_/D sky130_fd_sc_hd__clkbuf_1
X_20416_ _35472_/Q _35408_/Q _35344_/Q _35280_/Q _20260_/X _20261_/X VGND VGND VPWR
+ VPWR _20416_/X sky130_fd_sc_hd__mux4_1
X_24184_ _24184_/A VGND VGND VPWR VPWR _32628_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21396_ _33066_/Q _32042_/Q _35818_/Q _35754_/Q _21325_/X _21326_/X VGND VGND VPWR
+ VPWR _21396_/X sky130_fd_sc_hd__mux4_1
XFILLER_135_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23135_ _23135_/A VGND VGND VPWR VPWR _32106_/D sky130_fd_sc_hd__clkbuf_1
X_20347_ _33166_/Q _36046_/Q _33038_/Q _32974_/Q _20068_/X _20069_/X VGND VGND VPWR
+ VPWR _20347_/X sky130_fd_sc_hd__mux4_1
XFILLER_134_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28992_ _34806_/Q _27134_/X _29006_/S VGND VGND VPWR VPWR _28993_/A sky130_fd_sc_hd__mux2_1
XFILLER_134_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27943_ _27943_/A VGND VGND VPWR VPWR _34310_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23066_ _23066_/A VGND VGND VPWR VPWR _32079_/D sky130_fd_sc_hd__clkbuf_1
X_20278_ _33420_/Q _33356_/Q _33292_/Q _33228_/Q _20133_/X _20134_/X VGND VGND VPWR
+ VPWR _20278_/X sky130_fd_sc_hd__mux4_1
XFILLER_66_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22017_ _33148_/Q _36028_/Q _33020_/Q _32956_/Q _22015_/X _22016_/X VGND VGND VPWR
+ VPWR _22017_/X sky130_fd_sc_hd__mux4_1
XTAP_6169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27874_ _27874_/A VGND VGND VPWR VPWR _34277_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29613_ _35070_/Q _29453_/X _29631_/S VGND VGND VPWR VPWR _29614_/A sky130_fd_sc_hd__mux2_1
XTAP_4712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26825_ _33843_/Q _23384_/X _26825_/S VGND VGND VPWR VPWR _26826_/A sky130_fd_sc_hd__mux2_1
XFILLER_188_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29544_ _29544_/A VGND VGND VPWR VPWR _35037_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26756_ _26756_/A VGND VGND VPWR VPWR _33810_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_962 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23968_ _23968_/A VGND VGND VPWR VPWR _32528_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25707_ _25707_/A VGND VGND VPWR VPWR _33315_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29475_ input42/X VGND VGND VPWR VPWR _29475_/X sky130_fd_sc_hd__buf_2
X_22919_ _23083_/S VGND VGND VPWR VPWR _22947_/S sky130_fd_sc_hd__buf_4
X_26687_ _26687_/A VGND VGND VPWR VPWR _33777_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23899_ _23899_/A VGND VGND VPWR VPWR _32495_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_189_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16440_ _35616_/Q _34976_/Q _34336_/Q _33696_/Q _16438_/X _16439_/X VGND VGND VPWR
+ VPWR _16440_/X sky130_fd_sc_hd__mux4_1
X_28426_ _27708_/X _34539_/Q _28442_/S VGND VGND VPWR VPWR _28427_/A sky130_fd_sc_hd__mux2_1
X_25638_ _24939_/X _33283_/Q _25646_/S VGND VGND VPWR VPWR _25639_/A sky130_fd_sc_hd__mux2_1
XFILLER_232_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28357_ _28357_/A VGND VGND VPWR VPWR _34506_/D sky130_fd_sc_hd__clkbuf_1
X_16371_ _35422_/Q _35358_/Q _35294_/Q _35230_/Q _16195_/X _16196_/X VGND VGND VPWR
+ VPWR _16371_/X sky130_fd_sc_hd__mux4_1
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_386_CLK clkbuf_6_40__f_CLK/X VGND VGND VPWR VPWR _35641_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_13_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25569_ _24837_/X _33250_/Q _25583_/S VGND VGND VPWR VPWR _25570_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18110_ _32912_/Q _32848_/Q _32784_/Q _32720_/Q _15984_/X _15987_/X VGND VGND VPWR
+ VPWR _18110_/X sky130_fd_sc_hd__mux4_1
XFILLER_185_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27308_ _27308_/A VGND VGND VPWR VPWR _34040_/D sky130_fd_sc_hd__clkbuf_1
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19090_ _35690_/Q _32197_/Q _35562_/Q _35498_/Q _18911_/X _18912_/X VGND VGND VPWR
+ VPWR _19090_/X sky130_fd_sc_hd__mux4_1
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28288_ _28378_/S VGND VGND VPWR VPWR _28307_/S sky130_fd_sc_hd__buf_4
XFILLER_219_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18041_ _17905_/X _18039_/X _18040_/X _17910_/X VGND VGND VPWR VPWR _18041_/X sky130_fd_sc_hd__a22o_1
XFILLER_185_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_138_CLK clkbuf_6_22__f_CLK/X VGND VGND VPWR VPWR _35735_/CLK sky130_fd_sc_hd__clkbuf_16
X_27239_ _27239_/A VGND VGND VPWR VPWR _34007_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30250_ _35372_/Q _29398_/X _30264_/S VGND VGND VPWR VPWR _30251_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19992_ _33924_/Q _33860_/Q _33796_/Q _36100_/Q _19677_/X _19678_/X VGND VGND VPWR
+ VPWR _19992_/X sky130_fd_sc_hd__mux4_1
X_30181_ _30181_/A VGND VGND VPWR VPWR _35339_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_858 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18943_ _18661_/X _18939_/X _18942_/X _18665_/X VGND VGND VPWR VPWR _18943_/X sky130_fd_sc_hd__a22o_1
XFILLER_3_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_1443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33940_ _36179_/CLK _33940_/D VGND VGND VPWR VPWR _33940_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_310_CLK clkbuf_6_50__f_CLK/X VGND VGND VPWR VPWR _35974_/CLK sky130_fd_sc_hd__clkbuf_16
X_18874_ _20286_/A VGND VGND VPWR VPWR _18874_/X sky130_fd_sc_hd__buf_4
XTAP_6670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17825_ _34951_/Q _34887_/Q _34823_/Q _34759_/Q _17513_/X _17514_/X VGND VGND VPWR
+ VPWR _17825_/X sky130_fd_sc_hd__mux4_1
X_33871_ _34440_/CLK _33871_/D VGND VGND VPWR VPWR _33871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35610_ _35610_/CLK _35610_/D VGND VGND VPWR VPWR _35610_/Q sky130_fd_sc_hd__dfxtp_1
X_32822_ _32901_/CLK _32822_/D VGND VGND VPWR VPWR _32822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17756_ _17756_/A _17756_/B _17756_/C _17756_/D VGND VGND VPWR VPWR _17757_/A sky130_fd_sc_hd__or4_2
XFILLER_78_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16707_ _17766_/A VGND VGND VPWR VPWR _16707_/X sky130_fd_sc_hd__clkbuf_4
X_35541_ _35733_/CLK _35541_/D VGND VGND VPWR VPWR _35541_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32753_ _35953_/CLK _32753_/D VGND VGND VPWR VPWR _32753_/Q sky130_fd_sc_hd__dfxtp_1
X_17687_ _17687_/A VGND VGND VPWR VPWR _32003_/D sky130_fd_sc_hd__buf_4
XFILLER_223_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31704_ _36061_/Q input62/X _31708_/S VGND VGND VPWR VPWR _31705_/A sky130_fd_sc_hd__mux2_1
X_19426_ _19146_/X _19424_/X _19425_/X _19151_/X VGND VGND VPWR VPWR _19426_/X sky130_fd_sc_hd__a22o_1
X_35472_ _35599_/CLK _35472_/D VGND VGND VPWR VPWR _35472_/Q sky130_fd_sc_hd__dfxtp_1
X_16638_ _16353_/X _16636_/X _16637_/X _16359_/X VGND VGND VPWR VPWR _16638_/X sky130_fd_sc_hd__a22o_1
XFILLER_222_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32684_ _32914_/CLK _32684_/D VGND VGND VPWR VPWR _32684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34423_ _36150_/CLK _34423_/D VGND VGND VPWR VPWR _34423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19357_ _19153_/X _19355_/X _19356_/X _19156_/X VGND VGND VPWR VPWR _19357_/X sky130_fd_sc_hd__a22o_1
X_31635_ _31635_/A VGND VGND VPWR VPWR _36028_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16569_ _16565_/X _16568_/X _16426_/X VGND VGND VPWR VPWR _16595_/A sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_377_CLK clkbuf_6_43__f_CLK/X VGND VGND VPWR VPWR _35448_/CLK sky130_fd_sc_hd__clkbuf_16
X_18308_ _18361_/A VGND VGND VPWR VPWR _20260_/A sky130_fd_sc_hd__buf_12
XFILLER_13_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34354_ _35633_/CLK _34354_/D VGND VGND VPWR VPWR _34354_/Q sky130_fd_sc_hd__dfxtp_1
X_31566_ _31566_/A VGND VGND VPWR VPWR _35995_/D sky130_fd_sc_hd__clkbuf_1
X_19288_ _19284_/X _19287_/X _19079_/X VGND VGND VPWR VPWR _19318_/A sky130_fd_sc_hd__o21ba_1
XFILLER_129_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33305_ _33753_/CLK _33305_/D VGND VGND VPWR VPWR _33305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_777 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18239_ _18235_/X _18238_/X _17857_/A VGND VGND VPWR VPWR _18247_/C sky130_fd_sc_hd__o21ba_1
X_30517_ _30517_/A VGND VGND VPWR VPWR _35498_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_129_CLK clkbuf_6_21__f_CLK/X VGND VGND VPWR VPWR _35162_/CLK sky130_fd_sc_hd__clkbuf_16
X_34285_ _36141_/CLK _34285_/D VGND VGND VPWR VPWR _34285_/Q sky130_fd_sc_hd__dfxtp_1
X_31497_ _27757_/X _35963_/Q _31501_/S VGND VGND VPWR VPWR _31498_/A sky130_fd_sc_hd__mux2_1
XFILLER_198_1056 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33236_ _36180_/CLK _33236_/D VGND VGND VPWR VPWR _33236_/Q sky130_fd_sc_hd__dfxtp_1
X_21250_ _22464_/A VGND VGND VPWR VPWR _21250_/X sky130_fd_sc_hd__clkbuf_4
X_36024_ _36024_/CLK _36024_/D VGND VGND VPWR VPWR _36024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_758 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30448_ _35466_/Q _29491_/X _30462_/S VGND VGND VPWR VPWR _30449_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_950 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20201_ _20164_/X _20199_/X _20200_/X _20169_/X VGND VGND VPWR VPWR _20201_/X sky130_fd_sc_hd__a22o_1
X_33167_ _36047_/CLK _33167_/D VGND VGND VPWR VPWR _33167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21181_ _20892_/X _21179_/X _21180_/X _20895_/X VGND VGND VPWR VPWR _21181_/X sky130_fd_sc_hd__a22o_1
XFILLER_137_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30379_ _30379_/A VGND VGND VPWR VPWR _35433_/D sky130_fd_sc_hd__clkbuf_1
X_20132_ _19852_/X _20130_/X _20131_/X _19857_/X VGND VGND VPWR VPWR _20132_/X sky130_fd_sc_hd__a22o_1
X_32118_ _35895_/CLK _32118_/D VGND VGND VPWR VPWR _32118_/Q sky130_fd_sc_hd__dfxtp_1
X_33098_ _35849_/CLK _33098_/D VGND VGND VPWR VPWR _33098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20063_ _19859_/X _20061_/X _20062_/X _19862_/X VGND VGND VPWR VPWR _20063_/X sky130_fd_sc_hd__a22o_1
X_24940_ _24939_/X _32963_/Q _24952_/S VGND VGND VPWR VPWR _24941_/A sky130_fd_sc_hd__mux2_1
X_32049_ _36017_/CLK _32049_/D VGND VGND VPWR VPWR _32049_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_301_CLK clkbuf_6_57__f_CLK/X VGND VGND VPWR VPWR _35716_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24871_ input16/X VGND VGND VPWR VPWR _24871_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_6_1451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_940 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26610_ _24976_/X _33743_/Q _26614_/S VGND VGND VPWR VPWR _26611_/A sky130_fd_sc_hd__mux2_1
XTAP_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23822_ _23055_/X _32396_/Q _23832_/S VGND VGND VPWR VPWR _23823_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35808_ _35810_/CLK _35808_/D VGND VGND VPWR VPWR _35808_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27590_ _34174_/Q _27158_/X _27608_/S VGND VGND VPWR VPWR _27591_/A sky130_fd_sc_hd__mux2_1
XFILLER_245_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26541_ _24874_/X _33710_/Q _26551_/S VGND VGND VPWR VPWR _26542_/A sky130_fd_sc_hd__mux2_1
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35739_ _35802_/CLK _35739_/D VGND VGND VPWR VPWR _35739_/Q sky130_fd_sc_hd__dfxtp_1
X_20965_ _22515_/A VGND VGND VPWR VPWR _20965_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_54_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23753_ _22953_/X _32363_/Q _23769_/S VGND VGND VPWR VPWR _23754_/A sky130_fd_sc_hd__mux2_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22704_ _22512_/X _22702_/X _22703_/X _22515_/X VGND VGND VPWR VPWR _22704_/X sky130_fd_sc_hd__a22o_1
XFILLER_213_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29260_ _34933_/Q _27131_/X _29276_/S VGND VGND VPWR VPWR _29261_/A sky130_fd_sc_hd__mux2_1
XFILLER_246_1057 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26472_ _33678_/Q _23475_/X _26478_/S VGND VGND VPWR VPWR _26473_/A sky130_fd_sc_hd__mux2_1
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20896_ _20892_/X _20893_/X _20894_/X _20895_/X VGND VGND VPWR VPWR _20896_/X sky130_fd_sc_hd__a22o_1
X_23684_ _23055_/X _32332_/Q _23694_/S VGND VGND VPWR VPWR _23685_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1079 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28211_ _28211_/A VGND VGND VPWR VPWR _34437_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25423_ _24821_/X _33181_/Q _25427_/S VGND VGND VPWR VPWR _25424_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29191_ _34901_/Q _27229_/X _29191_/S VGND VGND VPWR VPWR _29192_/A sky130_fd_sc_hd__mux2_1
X_22635_ _22464_/X _22633_/X _22634_/X _22469_/X VGND VGND VPWR VPWR _22635_/X sky130_fd_sc_hd__a22o_1
XFILLER_41_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_368_CLK clkbuf_6_41__f_CLK/X VGND VGND VPWR VPWR _35833_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_213_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28142_ _28142_/A VGND VGND VPWR VPWR _34404_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_224_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22566_ _34699_/Q _34635_/Q _34571_/Q _34507_/Q _22245_/X _22246_/X VGND VGND VPWR
+ VPWR _22566_/X sky130_fd_sc_hd__mux4_1
X_25354_ _25354_/A VGND VGND VPWR VPWR _33149_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24305_ _24305_/A VGND VGND VPWR VPWR _32684_/D sky130_fd_sc_hd__clkbuf_1
X_21517_ _34158_/Q _34094_/Q _34030_/Q _33966_/Q _21340_/X _21341_/X VGND VGND VPWR
+ VPWR _21517_/X sky130_fd_sc_hd__mux4_1
X_28073_ _34372_/Q _27177_/X _28079_/S VGND VGND VPWR VPWR _28074_/A sky130_fd_sc_hd__mux2_1
X_22497_ _35209_/Q _35145_/Q _35081_/Q _32265_/Q _22316_/X _22317_/X VGND VGND VPWR
+ VPWR _22497_/X sky130_fd_sc_hd__mux4_1
X_25285_ _25285_/A VGND VGND VPWR VPWR _33116_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27024_ _27024_/A VGND VGND VPWR VPWR _33937_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24236_ _24236_/A VGND VGND VPWR VPWR _32653_/D sky130_fd_sc_hd__clkbuf_1
X_21448_ _22507_/A VGND VGND VPWR VPWR _21448_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_194_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24167_ _24167_/A VGND VGND VPWR VPWR _32620_/D sky130_fd_sc_hd__clkbuf_1
X_21379_ _22438_/A VGND VGND VPWR VPWR _21379_/X sky130_fd_sc_hd__buf_2
XFILLER_134_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23118_ _23118_/A VGND VGND VPWR VPWR _32098_/D sky130_fd_sc_hd__clkbuf_1
X_24098_ _24098_/A VGND VGND VPWR VPWR _32589_/D sky130_fd_sc_hd__clkbuf_1
X_28975_ _34798_/Q _27109_/X _28985_/S VGND VGND VPWR VPWR _28976_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27926_ _27766_/X _34302_/Q _27944_/S VGND VGND VPWR VPWR _27927_/A sky130_fd_sc_hd__mux2_1
XTAP_5210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23049_ input48/X VGND VGND VPWR VPWR _23049_/X sky130_fd_sc_hd__buf_2
XTAP_5221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_237_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27857_ _27857_/A VGND VGND VPWR VPWR _34269_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17610_ _33089_/Q _32065_/Q _35841_/Q _35777_/Q _17431_/X _17432_/X VGND VGND VPWR
+ VPWR _17610_/X sky130_fd_sc_hd__mux4_1
XTAP_4542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26808_ _26808_/A VGND VGND VPWR VPWR _33834_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18590_ _18330_/X _18586_/X _18589_/X _18341_/X VGND VGND VPWR VPWR _18590_/X sky130_fd_sc_hd__a22o_1
XTAP_4564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27788_ input42/X VGND VGND VPWR VPWR _27788_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29527_ _29797_/A _30607_/B VGND VGND VPWR VPWR _29660_/S sky130_fd_sc_hd__nor2_8
XTAP_4597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17541_ _17356_/X _17539_/X _17540_/X _17359_/X VGND VGND VPWR VPWR _17541_/X sky130_fd_sc_hd__a22o_1
XTAP_3852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26739_ _33802_/Q _23463_/X _26753_/S VGND VGND VPWR VPWR _26740_/A sky130_fd_sc_hd__mux2_1
XTAP_3863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29458_ _35007_/Q _29457_/X _29482_/S VGND VGND VPWR VPWR _29459_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17472_ _34941_/Q _34877_/Q _34813_/Q _34749_/Q _17160_/X _17161_/X VGND VGND VPWR
+ VPWR _17472_/X sky130_fd_sc_hd__mux4_1
XFILLER_205_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19211_ _34925_/Q _34861_/Q _34797_/Q _34733_/Q _19107_/X _19108_/X VGND VGND VPWR
+ VPWR _19211_/X sky130_fd_sc_hd__mux4_1
XFILLER_232_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16423_ _33376_/Q _33312_/Q _33248_/Q _33184_/Q _16421_/X _16422_/X VGND VGND VPWR
+ VPWR _16423_/X sky130_fd_sc_hd__mux4_1
X_28409_ _27683_/X _34531_/Q _28421_/S VGND VGND VPWR VPWR _28410_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29389_ _34985_/Q _29388_/X _29389_/S VGND VGND VPWR VPWR _29390_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_359_CLK clkbuf_6_46__f_CLK/X VGND VGND VPWR VPWR _35194_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_125_1220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31420_ _27639_/X _35926_/Q _31438_/S VGND VGND VPWR VPWR _31421_/A sky130_fd_sc_hd__mux2_1
X_19142_ _19105_/X _19140_/X _19141_/X _19110_/X VGND VGND VPWR VPWR _19142_/X sky130_fd_sc_hd__a22o_1
XFILLER_125_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16354_ _17766_/A VGND VGND VPWR VPWR _16354_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_81_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19073_ _18793_/X _19071_/X _19072_/X _18798_/X VGND VGND VPWR VPWR _19073_/X sky130_fd_sc_hd__a22o_1
X_31351_ _31351_/A VGND VGND VPWR VPWR _35893_/D sky130_fd_sc_hd__clkbuf_1
X_16285_ _16018_/X _16283_/X _16284_/X _16027_/X VGND VGND VPWR VPWR _16285_/X sky130_fd_sc_hd__a22o_1
XFILLER_8_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18024_ _35661_/Q _35021_/Q _34381_/Q _33741_/Q _17850_/X _17851_/X VGND VGND VPWR
+ VPWR _18024_/X sky130_fd_sc_hd__mux4_1
X_30302_ _35397_/Q _29475_/X _30306_/S VGND VGND VPWR VPWR _30303_/A sky130_fd_sc_hd__mux2_1
X_34070_ _34070_/CLK _34070_/D VGND VGND VPWR VPWR _34070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31282_ _31282_/A VGND VGND VPWR VPWR _35861_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33021_ _36029_/CLK _33021_/D VGND VGND VPWR VPWR _33021_/Q sky130_fd_sc_hd__dfxtp_1
X_30233_ _35364_/Q _29373_/X _30243_/S VGND VGND VPWR VPWR _30234_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30164_ _30164_/A VGND VGND VPWR VPWR _35331_/D sky130_fd_sc_hd__clkbuf_1
X_19975_ _35459_/Q _35395_/Q _35331_/Q _35267_/Q _19907_/X _19908_/X VGND VGND VPWR
+ VPWR _19975_/X sky130_fd_sc_hd__mux4_1
XFILLER_114_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18926_ _18922_/X _18925_/X _18759_/X VGND VGND VPWR VPWR _18927_/D sky130_fd_sc_hd__o21ba_1
XFILLER_68_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34972_ _36058_/CLK _34972_/D VGND VGND VPWR VPWR _34972_/Q sky130_fd_sc_hd__dfxtp_1
X_30095_ _30095_/A VGND VGND VPWR VPWR _35298_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33923_ _36101_/CLK _33923_/D VGND VGND VPWR VPWR _33923_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18857_ _34403_/Q _36131_/Q _34275_/Q _34211_/Q _18823_/X _18824_/X VGND VGND VPWR
+ VPWR _18857_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17808_ _33159_/Q _36039_/Q _33031_/Q _32967_/Q _17768_/X _17769_/X VGND VGND VPWR
+ VPWR _17808_/X sky130_fd_sc_hd__mux4_1
XFILLER_82_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33854_ _35456_/CLK _33854_/D VGND VGND VPWR VPWR _33854_/Q sky130_fd_sc_hd__dfxtp_1
X_18788_ _34913_/Q _34849_/Q _34785_/Q _34721_/Q _18754_/X _18755_/X VGND VGND VPWR
+ VPWR _18788_/X sky130_fd_sc_hd__mux4_1
XFILLER_48_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_243_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32805_ _32869_/CLK _32805_/D VGND VGND VPWR VPWR _32805_/Q sky130_fd_sc_hd__dfxtp_1
X_17739_ _32901_/Q _32837_/Q _32773_/Q _32709_/Q _17699_/X _17700_/X VGND VGND VPWR
+ VPWR _17739_/X sky130_fd_sc_hd__mux4_1
X_30997_ _30997_/A VGND VGND VPWR VPWR _35726_/D sky130_fd_sc_hd__clkbuf_1
X_33785_ _33850_/CLK _33785_/D VGND VGND VPWR VPWR _33785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35524_ _35843_/CLK _35524_/D VGND VGND VPWR VPWR _35524_/Q sky130_fd_sc_hd__dfxtp_1
X_20750_ _22469_/A VGND VGND VPWR VPWR _20750_/X sky130_fd_sc_hd__buf_6
X_32736_ _33119_/CLK _32736_/D VGND VGND VPWR VPWR _32736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19409_ _35635_/Q _34995_/Q _34355_/Q _33715_/Q _19091_/X _19092_/X VGND VGND VPWR
+ VPWR _19409_/X sky130_fd_sc_hd__mux4_1
X_20681_ _34646_/Q _34582_/Q _34518_/Q _34454_/Q _20679_/X _20680_/X VGND VGND VPWR
+ VPWR _20681_/X sky130_fd_sc_hd__mux4_1
X_32667_ _35669_/CLK _32667_/D VGND VGND VPWR VPWR _32667_/Q sky130_fd_sc_hd__dfxtp_1
X_35455_ _35456_/CLK _35455_/D VGND VGND VPWR VPWR _35455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22420_ _22416_/X _22419_/X _22104_/X VGND VGND VPWR VPWR _22428_/C sky130_fd_sc_hd__o21ba_1
XFILLER_17_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34406_ _34914_/CLK _34406_/D VGND VGND VPWR VPWR _34406_/Q sky130_fd_sc_hd__dfxtp_1
X_31618_ _27735_/X _36020_/Q _31636_/S VGND VGND VPWR VPWR _31619_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32598_ _35990_/CLK _32598_/D VGND VGND VPWR VPWR _32598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35386_ _35451_/CLK _35386_/D VGND VGND VPWR VPWR _35386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_906 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22351_ _22106_/X _22349_/X _22350_/X _22109_/X VGND VGND VPWR VPWR _22351_/X sky130_fd_sc_hd__a22o_1
XFILLER_149_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31549_ _27834_/X _35988_/Q _31551_/S VGND VGND VPWR VPWR _31550_/A sky130_fd_sc_hd__mux2_1
XFILLER_136_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34337_ _35618_/CLK _34337_/D VGND VGND VPWR VPWR _34337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21302_ _33384_/Q _33320_/Q _33256_/Q _33192_/Q _21021_/X _21022_/X VGND VGND VPWR
+ VPWR _21302_/X sky130_fd_sc_hd__mux4_1
XFILLER_148_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25070_ _24905_/X _33016_/Q _25080_/S VGND VGND VPWR VPWR _25071_/A sky130_fd_sc_hd__mux2_1
X_34268_ _36235_/CLK _34268_/D VGND VGND VPWR VPWR _34268_/Q sky130_fd_sc_hd__dfxtp_1
X_22282_ _34435_/Q _36163_/Q _34307_/Q _34243_/Q _22182_/X _22183_/X VGND VGND VPWR
+ VPWR _22282_/X sky130_fd_sc_hd__mux4_1
XFILLER_102_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24021_ _22946_/X _32553_/Q _24021_/S VGND VGND VPWR VPWR _24022_/A sky130_fd_sc_hd__mux2_1
XFILLER_219_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33219_ _33415_/CLK _33219_/D VGND VGND VPWR VPWR _33219_/Q sky130_fd_sc_hd__dfxtp_1
X_21233_ _33894_/Q _33830_/Q _33766_/Q _36070_/Q _20918_/X _20919_/X VGND VGND VPWR
+ VPWR _21233_/X sky130_fd_sc_hd__mux4_1
X_36007_ _36007_/CLK _36007_/D VGND VGND VPWR VPWR _36007_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1023 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34199_ _34773_/CLK _34199_/D VGND VGND VPWR VPWR _34199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21164_ _34148_/Q _34084_/Q _34020_/Q _33956_/Q _20987_/X _20988_/X VGND VGND VPWR
+ VPWR _21164_/X sky130_fd_sc_hd__mux4_1
XFILLER_236_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_1310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20115_ _35655_/Q _35015_/Q _34375_/Q _33735_/Q _19797_/X _19798_/X VGND VGND VPWR
+ VPWR _20115_/X sky130_fd_sc_hd__mux4_1
XFILLER_172_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28760_ _34697_/Q _27193_/X _28776_/S VGND VGND VPWR VPWR _28761_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_1332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21095_ _22507_/A VGND VGND VPWR VPWR _21095_/X sky130_fd_sc_hd__buf_4
X_25972_ _24834_/X _33441_/Q _25988_/S VGND VGND VPWR VPWR _25973_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_1302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27711_ input15/X VGND VGND VPWR VPWR _27711_/X sky130_fd_sc_hd__buf_2
XFILLER_246_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20046_ _33093_/Q _32069_/Q _35845_/Q _35781_/Q _19731_/X _19732_/X VGND VGND VPWR
+ VPWR _20046_/X sky130_fd_sc_hd__mux4_1
XFILLER_154_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24923_ input35/X VGND VGND VPWR VPWR _24923_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_115_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28691_ _28691_/A VGND VGND VPWR VPWR _34664_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27642_ _31283_/B _31823_/B VGND VGND VPWR VPWR _27838_/S sky130_fd_sc_hd__nand2_8
XFILLER_58_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24854_ _24854_/A VGND VGND VPWR VPWR _32935_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_206_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23805_ _23030_/X _32388_/Q _23811_/S VGND VGND VPWR VPWR _23806_/A sky130_fd_sc_hd__mux2_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27573_ _34166_/Q _27134_/X _27587_/S VGND VGND VPWR VPWR _27574_/A sky130_fd_sc_hd__mux2_1
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24785_ _24785_/A VGND VGND VPWR VPWR _32912_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21997_ _35195_/Q _35131_/Q _35067_/Q _32251_/Q _21963_/X _21964_/X VGND VGND VPWR
+ VPWR _21997_/X sky130_fd_sc_hd__mux4_1
X_29312_ _34958_/Q _27208_/X _29318_/S VGND VGND VPWR VPWR _29313_/A sky130_fd_sc_hd__mux2_1
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26524_ _24849_/X _33702_/Q _26530_/S VGND VGND VPWR VPWR _26525_/A sky130_fd_sc_hd__mux2_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23736_ _22928_/X _32355_/Q _23748_/S VGND VGND VPWR VPWR _23737_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20948_ _20740_/X _20946_/X _20947_/X _20745_/X VGND VGND VPWR VPWR _20948_/X sky130_fd_sc_hd__a22o_1
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29243_ _34925_/Q _27106_/X _29255_/S VGND VGND VPWR VPWR _29244_/A sky130_fd_sc_hd__mux2_1
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26455_ _33670_/Q _23447_/X _26457_/S VGND VGND VPWR VPWR _26456_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23667_ _23030_/X _32324_/Q _23673_/S VGND VGND VPWR VPWR _23668_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20879_ _33372_/Q _33308_/Q _33244_/Q _33180_/Q _20602_/X _20603_/X VGND VGND VPWR
+ VPWR _20879_/X sky130_fd_sc_hd__mux4_1
XFILLER_197_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25406_ _25406_/A VGND VGND VPWR VPWR _26352_/B sky130_fd_sc_hd__buf_12
X_29174_ _29174_/A VGND VGND VPWR VPWR _34892_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22618_ _22365_/X _22616_/X _22617_/X _22371_/X VGND VGND VPWR VPWR _22618_/X sky130_fd_sc_hd__a22o_1
XFILLER_41_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26386_ _33637_/Q _23277_/X _26394_/S VGND VGND VPWR VPWR _26387_/A sky130_fd_sc_hd__mux2_1
XFILLER_197_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23598_ _22928_/X _32291_/Q _23610_/S VGND VGND VPWR VPWR _23599_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28125_ _28125_/A VGND VGND VPWR VPWR _34396_/D sky130_fd_sc_hd__clkbuf_1
X_25337_ _33141_/Q _23393_/X _25353_/S VGND VGND VPWR VPWR _25338_/A sky130_fd_sc_hd__mux2_1
X_22549_ _22545_/X _22548_/X _22438_/X VGND VGND VPWR VPWR _22573_/A sky130_fd_sc_hd__o21ba_1
XFILLER_202_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16070_ _33046_/Q _32022_/Q _35798_/Q _35734_/Q _16067_/X _16069_/X VGND VGND VPWR
+ VPWR _16070_/X sky130_fd_sc_hd__mux4_1
XFILLER_127_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_1180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28056_ _34364_/Q _27152_/X _28058_/S VGND VGND VPWR VPWR _28057_/A sky130_fd_sc_hd__mux2_1
X_25268_ _25268_/A VGND VGND VPWR VPWR _33109_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27007_ _33929_/Q _23460_/X _27023_/S VGND VGND VPWR VPWR _27008_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_728 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24219_ _24219_/A VGND VGND VPWR VPWR _32645_/D sky130_fd_sc_hd__clkbuf_1
X_25199_ _33076_/Q _23387_/X _25217_/S VGND VGND VPWR VPWR _25200_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16972_ _16968_/X _16971_/X _16798_/X VGND VGND VPWR VPWR _16980_/C sky130_fd_sc_hd__o21ba_1
X_19760_ _19756_/X _19759_/X _19440_/X _19441_/X VGND VGND VPWR VPWR _19775_/B sky130_fd_sc_hd__o211a_1
X_28958_ _34790_/Q _27084_/X _28964_/S VGND VGND VPWR VPWR _28959_/A sky130_fd_sc_hd__mux2_1
XFILLER_231_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18711_ _18378_/X _18709_/X _18710_/X _18388_/X VGND VGND VPWR VPWR _18711_/X sky130_fd_sc_hd__a22o_1
XFILLER_231_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27909_ _27742_/X _34294_/Q _27923_/S VGND VGND VPWR VPWR _27910_/A sky130_fd_sc_hd__mux2_1
X_19691_ _19651_/X _19689_/X _19690_/X _19654_/X VGND VGND VPWR VPWR _19691_/X sky130_fd_sc_hd__a22o_1
X_28889_ _28889_/A VGND VGND VPWR VPWR _34757_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18642_ _18391_/X _18640_/X _18641_/X _18401_/X VGND VGND VPWR VPWR _18642_/X sky130_fd_sc_hd__a22o_1
XTAP_5084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30920_ _31010_/S VGND VGND VPWR VPWR _30939_/S sky130_fd_sc_hd__buf_6
XTAP_4350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18573_ _18569_/X _18572_/X _18404_/X VGND VGND VPWR VPWR _18574_/D sky130_fd_sc_hd__o21ba_1
X_30851_ _35657_/Q input47/X _30867_/S VGND VGND VPWR VPWR _30852_/A sky130_fd_sc_hd__mux2_1
XTAP_4394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17524_ _17199_/X _17522_/X _17523_/X _17204_/X VGND VGND VPWR VPWR _17524_/X sky130_fd_sc_hd__a22o_1
XFILLER_189_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33570_ _33573_/CLK _33570_/D VGND VGND VPWR VPWR _33570_/Q sky130_fd_sc_hd__dfxtp_1
X_30782_ _30782_/A VGND VGND VPWR VPWR _35624_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32521_ _35978_/CLK _32521_/D VGND VGND VPWR VPWR _32521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_935 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17455_ _33149_/Q _36029_/Q _33021_/Q _32957_/Q _17415_/X _17416_/X VGND VGND VPWR
+ VPWR _17455_/X sky130_fd_sc_hd__mux4_1
XFILLER_232_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16406_ _33055_/Q _32031_/Q _35807_/Q _35743_/Q _16372_/X _16373_/X VGND VGND VPWR
+ VPWR _16406_/X sky130_fd_sc_hd__mux4_1
X_32452_ _36085_/CLK _32452_/D VGND VGND VPWR VPWR _32452_/Q sky130_fd_sc_hd__dfxtp_1
X_35240_ _35685_/CLK _35240_/D VGND VGND VPWR VPWR _35240_/Q sky130_fd_sc_hd__dfxtp_1
X_17386_ _32891_/Q _32827_/Q _32763_/Q _32699_/Q _17346_/X _17347_/X VGND VGND VPWR
+ VPWR _17386_/X sky130_fd_sc_hd__mux4_1
XFILLER_125_1050 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31403_ _31403_/A VGND VGND VPWR VPWR _35918_/D sky130_fd_sc_hd__clkbuf_1
X_19125_ _19006_/X _19123_/X _19124_/X _19012_/X VGND VGND VPWR VPWR _19125_/X sky130_fd_sc_hd__a22o_1
X_16337_ _34653_/Q _34589_/Q _34525_/Q _34461_/Q _16233_/X _16234_/X VGND VGND VPWR
+ VPWR _16337_/X sky130_fd_sc_hd__mux4_1
X_35171_ _36210_/CLK _35171_/D VGND VGND VPWR VPWR _35171_/Q sky130_fd_sc_hd__dfxtp_1
X_32383_ _32896_/CLK _32383_/D VGND VGND VPWR VPWR _32383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34122_ _34186_/CLK _34122_/D VGND VGND VPWR VPWR _34122_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19056_ _35625_/Q _34985_/Q _34345_/Q _33705_/Q _18738_/X _18739_/X VGND VGND VPWR
+ VPWR _19056_/X sky130_fd_sc_hd__mux4_1
X_31334_ _31334_/A VGND VGND VPWR VPWR _35885_/D sky130_fd_sc_hd__clkbuf_1
X_16268_ _35163_/Q _35099_/Q _35035_/Q _32155_/Q _16083_/X _16085_/X VGND VGND VPWR
+ VPWR _16268_/X sky130_fd_sc_hd__mux4_1
X_18007_ _18007_/A _18007_/B _18007_/C _18007_/D VGND VGND VPWR VPWR _18008_/A sky130_fd_sc_hd__or4_2
XFILLER_161_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34053_ _34183_/CLK _34053_/D VGND VGND VPWR VPWR _34053_/Q sky130_fd_sc_hd__dfxtp_1
X_31265_ _27813_/X _35853_/Q _31273_/S VGND VGND VPWR VPWR _31266_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16199_ _16060_/X _16197_/X _16198_/X _16072_/X VGND VGND VPWR VPWR _16199_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_504_CLK clkbuf_leaf_2_CLK/A VGND VGND VPWR VPWR _36066_/CLK sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_60_CLK clkbuf_leaf_61_CLK/A VGND VGND VPWR VPWR _32914_/CLK sky130_fd_sc_hd__clkbuf_16
X_33004_ _36141_/CLK _33004_/D VGND VGND VPWR VPWR _33004_/Q sky130_fd_sc_hd__dfxtp_1
X_30216_ _35356_/Q _29348_/X _30222_/S VGND VGND VPWR VPWR _30217_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31196_ _27711_/X _35820_/Q _31210_/S VGND VGND VPWR VPWR _31197_/A sky130_fd_sc_hd__mux2_1
XFILLER_236_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30147_ _30147_/A VGND VGND VPWR VPWR _35323_/D sky130_fd_sc_hd__clkbuf_1
X_19958_ _19852_/X _19956_/X _19957_/X _19857_/X VGND VGND VPWR VPWR _19958_/X sky130_fd_sc_hd__a22o_1
XFILLER_45_1051 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18909_ _18661_/X _18907_/X _18908_/X _18665_/X VGND VGND VPWR VPWR _18909_/X sky130_fd_sc_hd__a22o_1
X_34955_ _34957_/CLK _34955_/D VGND VGND VPWR VPWR _34955_/Q sky130_fd_sc_hd__dfxtp_1
X_30078_ _30078_/A VGND VGND VPWR VPWR _35290_/D sky130_fd_sc_hd__clkbuf_1
X_19889_ _19889_/A VGND VGND VPWR VPWR _32448_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_142_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33906_ _34099_/CLK _33906_/D VGND VGND VPWR VPWR _33906_/Q sky130_fd_sc_hd__dfxtp_1
X_21920_ _35641_/Q _35001_/Q _34361_/Q _33721_/Q _21744_/X _21745_/X VGND VGND VPWR
+ VPWR _21920_/X sky130_fd_sc_hd__mux4_1
XFILLER_55_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34886_ _36165_/CLK _34886_/D VGND VGND VPWR VPWR _34886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_222_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33837_ _36076_/CLK _33837_/D VGND VGND VPWR VPWR _33837_/Q sky130_fd_sc_hd__dfxtp_1
X_21851_ _35703_/Q _32212_/Q _35575_/Q _35511_/Q _21564_/X _21565_/X VGND VGND VPWR
+ VPWR _21851_/X sky130_fd_sc_hd__mux4_1
XFILLER_71_918 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20802_ _35161_/Q _35097_/Q _35033_/Q _32153_/Q _20683_/X _20685_/X VGND VGND VPWR
+ VPWR _20802_/X sky130_fd_sc_hd__mux4_1
XFILLER_64_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24570_ _22949_/X _32810_/Q _24588_/S VGND VGND VPWR VPWR _24571_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21782_ _21778_/X _21781_/X _21740_/X _21741_/X VGND VGND VPWR VPWR _21797_/B sky130_fd_sc_hd__o211a_1
XFILLER_230_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33768_ _36073_/CLK _33768_/D VGND VGND VPWR VPWR _33768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23521_ _23521_/A VGND VGND VPWR VPWR _32255_/D sky130_fd_sc_hd__clkbuf_1
X_35507_ _35699_/CLK _35507_/D VGND VGND VPWR VPWR _35507_/Q sky130_fd_sc_hd__dfxtp_1
X_20733_ _20678_/X _20731_/X _20732_/X _20688_/X VGND VGND VPWR VPWR _20733_/X sky130_fd_sc_hd__a22o_1
XFILLER_180_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32719_ _32879_/CLK _32719_/D VGND VGND VPWR VPWR _32719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33699_ _35177_/CLK _33699_/D VGND VGND VPWR VPWR _33699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26240_ _24830_/X _33568_/Q _26258_/S VGND VGND VPWR VPWR _26241_/A sky130_fd_sc_hd__mux2_1
X_20664_ _22451_/A VGND VGND VPWR VPWR _20664_/X sky130_fd_sc_hd__buf_4
X_23452_ _23452_/A VGND VGND VPWR VPWR _32229_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35438_ _35438_/CLK _35438_/D VGND VGND VPWR VPWR _35438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22403_ _33415_/Q _33351_/Q _33287_/Q _33223_/Q _22080_/X _22081_/X VGND VGND VPWR
+ VPWR _22403_/X sky130_fd_sc_hd__mux4_1
XFILLER_13_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_1055 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26171_ _26171_/A VGND VGND VPWR VPWR _33535_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23383_ _23383_/A VGND VGND VPWR VPWR _32206_/D sky130_fd_sc_hd__clkbuf_1
X_20595_ _22400_/A VGND VGND VPWR VPWR _20595_/X sky130_fd_sc_hd__clkbuf_4
X_35369_ _35433_/CLK _35369_/D VGND VGND VPWR VPWR _35369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25122_ _24982_/X _33041_/Q _25122_/S VGND VGND VPWR VPWR _25123_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22334_ _22328_/X _22333_/X _22085_/X VGND VGND VPWR VPWR _22356_/A sky130_fd_sc_hd__o21ba_1
XFILLER_178_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29930_ _35221_/Q _29524_/X _29930_/S VGND VGND VPWR VPWR _29931_/A sky130_fd_sc_hd__mux2_1
X_22265_ _22012_/X _22263_/X _22264_/X _22018_/X VGND VGND VPWR VPWR _22265_/X sky130_fd_sc_hd__a22o_1
X_25053_ _24880_/X _33008_/Q _25059_/S VGND VGND VPWR VPWR _25054_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_51_CLK clkbuf_leaf_57_CLK/A VGND VGND VPWR VPWR _32552_/CLK sky130_fd_sc_hd__clkbuf_16
X_24004_ _24004_/A VGND VGND VPWR VPWR _32544_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21216_ _35429_/Q _35365_/Q _35301_/Q _35237_/Q _21148_/X _21149_/X VGND VGND VPWR
+ VPWR _21216_/X sky130_fd_sc_hd__mux4_1
XFILLER_183_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_1427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29861_ _29930_/S VGND VGND VPWR VPWR _29880_/S sky130_fd_sc_hd__buf_4
X_22196_ _22192_/X _22195_/X _22085_/X VGND VGND VPWR VPWR _22220_/A sky130_fd_sc_hd__o21ba_1
XFILLER_2_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28812_ _28812_/A VGND VGND VPWR VPWR _34720_/D sky130_fd_sc_hd__clkbuf_1
X_21147_ _20892_/X _21145_/X _21146_/X _20895_/X VGND VGND VPWR VPWR _21147_/X sky130_fd_sc_hd__a22o_1
X_29792_ _29792_/A VGND VGND VPWR VPWR _35155_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28743_ _34689_/Q _27168_/X _28755_/S VGND VGND VPWR VPWR _28744_/A sky130_fd_sc_hd__mux2_1
X_25955_ _24809_/X _33433_/Q _25967_/S VGND VGND VPWR VPWR _25956_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21078_ _35617_/Q _34977_/Q _34337_/Q _33697_/Q _21038_/X _21039_/X VGND VGND VPWR
+ VPWR _21078_/X sky130_fd_sc_hd__mux4_2
XFILLER_74_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20029_ _33413_/Q _33349_/Q _33285_/Q _33221_/Q _19780_/X _19781_/X VGND VGND VPWR
+ VPWR _20029_/X sky130_fd_sc_hd__mux4_1
X_24906_ _24905_/X _32952_/Q _24921_/S VGND VGND VPWR VPWR _24907_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_1165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28674_ _34656_/Q _27065_/X _28692_/S VGND VGND VPWR VPWR _28675_/A sky130_fd_sc_hd__mux2_1
X_25886_ _25886_/A VGND VGND VPWR VPWR _33400_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_246_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27625_ _34191_/Q _27211_/X _27629_/S VGND VGND VPWR VPWR _27626_/A sky130_fd_sc_hd__mux2_1
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24837_ input4/X VGND VGND VPWR VPWR _24837_/X sky130_fd_sc_hd__buf_4
XFILLER_62_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27556_ _34158_/Q _27109_/X _27566_/S VGND VGND VPWR VPWR _27557_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24768_ _23042_/X _32904_/Q _24786_/S VGND VGND VPWR VPWR _24769_/A sky130_fd_sc_hd__mux2_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26507_ _24824_/X _33694_/Q _26509_/S VGND VGND VPWR VPWR _26508_/A sky130_fd_sc_hd__mux2_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23719_ _22903_/X _32347_/Q _23727_/S VGND VGND VPWR VPWR _23720_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27487_ _27487_/A VGND VGND VPWR VPWR _34125_/D sky130_fd_sc_hd__clkbuf_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24699_ _24699_/A VGND VGND VPWR VPWR _32871_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17240_ _33399_/Q _33335_/Q _33271_/Q _33207_/Q _17127_/X _17128_/X VGND VGND VPWR
+ VPWR _17240_/X sky130_fd_sc_hd__mux4_1
X_29226_ _34917_/Q _27081_/X _29234_/S VGND VGND VPWR VPWR _29227_/A sky130_fd_sc_hd__mux2_1
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26438_ _26486_/S VGND VGND VPWR VPWR _26457_/S sky130_fd_sc_hd__buf_6
XFILLER_35_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29157_ _29157_/A VGND VGND VPWR VPWR _34884_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17171_ _16846_/X _17169_/X _17170_/X _16851_/X VGND VGND VPWR VPWR _17171_/X sky130_fd_sc_hd__a22o_1
XFILLER_167_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26369_ _33629_/Q _23252_/X _26373_/S VGND VGND VPWR VPWR _26370_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16122_ _16030_/X _16120_/X _16121_/X _16041_/X VGND VGND VPWR VPWR _16122_/X sky130_fd_sc_hd__a22o_1
X_28108_ _34389_/Q _27229_/X _28108_/S VGND VGND VPWR VPWR _28109_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29088_ _29088_/A VGND VGND VPWR VPWR _34851_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16053_ _17998_/A VGND VGND VPWR VPWR _16053_/X sky130_fd_sc_hd__buf_6
XFILLER_183_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28039_ _28108_/S VGND VGND VPWR VPWR _28058_/S sky130_fd_sc_hd__buf_4
XFILLER_196_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_42_CLK clkbuf_6_6__f_CLK/X VGND VGND VPWR VPWR _35810_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_108_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_6_48__f_CLK clkbuf_5_24_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_48__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_31050_ _31050_/A VGND VGND VPWR VPWR _35751_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_1046 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30001_ _35254_/Q _29429_/X _30015_/S VGND VGND VPWR VPWR _30002_/A sky130_fd_sc_hd__mux2_1
X_19812_ _34430_/Q _36158_/Q _34302_/Q _34238_/Q _19529_/X _19530_/X VGND VGND VPWR
+ VPWR _19812_/X sky130_fd_sc_hd__mux4_1
XFILLER_69_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19743_ _19743_/A _19743_/B _19743_/C _19743_/D VGND VGND VPWR VPWR _19744_/A sky130_fd_sc_hd__or4_2
X_16955_ _16853_/X _16953_/X _16954_/X _16856_/X VGND VGND VPWR VPWR _16955_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_238_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34740_ _35124_/CLK _34740_/D VGND VGND VPWR VPWR _34740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31952_ _23492_/X _36179_/Q _31956_/S VGND VGND VPWR VPWR _31953_/A sky130_fd_sc_hd__mux2_1
X_19674_ _34171_/Q _34107_/Q _34043_/Q _33979_/Q _19393_/X _19394_/X VGND VGND VPWR
+ VPWR _19674_/X sky130_fd_sc_hd__mux4_1
X_16886_ _16846_/X _16884_/X _16885_/X _16851_/X VGND VGND VPWR VPWR _16886_/X sky130_fd_sc_hd__a22o_1
XFILLER_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18625_ _18318_/X _18623_/X _18624_/X _18327_/X VGND VGND VPWR VPWR _18625_/X sky130_fd_sc_hd__a22o_1
X_30903_ _30903_/A VGND VGND VPWR VPWR _35681_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_237_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34671_ _34926_/CLK _34671_/D VGND VGND VPWR VPWR _34671_/Q sky130_fd_sc_hd__dfxtp_1
X_31883_ _23381_/X _36146_/Q _31885_/S VGND VGND VPWR VPWR _31884_/A sky130_fd_sc_hd__mux2_1
XTAP_4191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30834_ _35649_/Q input38/X _30846_/S VGND VGND VPWR VPWR _30835_/A sky130_fd_sc_hd__mux2_1
X_33622_ _35997_/CLK _33622_/D VGND VGND VPWR VPWR _33622_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18556_ _18330_/X _18554_/X _18555_/X _18341_/X VGND VGND VPWR VPWR _18556_/X sky130_fd_sc_hd__a22o_1
XFILLER_52_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17507_ _34686_/Q _34622_/Q _34558_/Q _34494_/Q _17292_/X _17293_/X VGND VGND VPWR
+ VPWR _17507_/X sky130_fd_sc_hd__mux4_1
X_33553_ _34441_/CLK _33553_/D VGND VGND VPWR VPWR _33553_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18487_ _18318_/X _18485_/X _18486_/X _18327_/X VGND VGND VPWR VPWR _18487_/X sky130_fd_sc_hd__a22o_1
X_30765_ _35616_/Q input2/X _30783_/S VGND VGND VPWR VPWR _30766_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17438_ _17153_/X _17436_/X _17437_/X _17156_/X VGND VGND VPWR VPWR _17438_/X sky130_fd_sc_hd__a22o_1
X_32504_ _35961_/CLK _32504_/D VGND VGND VPWR VPWR _32504_/Q sky130_fd_sc_hd__dfxtp_1
X_33484_ _33934_/CLK _33484_/D VGND VGND VPWR VPWR _33484_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30696_ _30696_/A VGND VGND VPWR VPWR _35583_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35223_ _35799_/CLK _35223_/D VGND VGND VPWR VPWR _35223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32435_ _33897_/CLK _32435_/D VGND VGND VPWR VPWR _32435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17369_ _17158_/X _17367_/X _17368_/X _17163_/X VGND VGND VPWR VPWR _17369_/X sky130_fd_sc_hd__a22o_1
XFILLER_105_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19108_ _19461_/A VGND VGND VPWR VPWR _19108_/X sky130_fd_sc_hd__clkbuf_4
X_35154_ _35730_/CLK _35154_/D VGND VGND VPWR VPWR _35154_/Q sky130_fd_sc_hd__dfxtp_1
X_20380_ _32911_/Q _32847_/Q _32783_/Q _32719_/Q _18284_/X _18287_/X VGND VGND VPWR
+ VPWR _20380_/X sky130_fd_sc_hd__mux4_1
X_32366_ _35951_/CLK _32366_/D VGND VGND VPWR VPWR _32366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34105_ _35641_/CLK _34105_/D VGND VGND VPWR VPWR _34105_/Q sky130_fd_sc_hd__dfxtp_1
X_19039_ _33641_/Q _33577_/Q _33513_/Q _33449_/Q _18794_/X _18795_/X VGND VGND VPWR
+ VPWR _19039_/X sky130_fd_sc_hd__mux4_1
X_31317_ _31317_/A VGND VGND VPWR VPWR _35877_/D sky130_fd_sc_hd__clkbuf_1
X_35085_ _35663_/CLK _35085_/D VGND VGND VPWR VPWR _35085_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput100 _31977_/Q VGND VGND VPWR VPWR D1[19] sky130_fd_sc_hd__buf_2
X_32297_ _35947_/CLK _32297_/D VGND VGND VPWR VPWR _32297_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput111 _31987_/Q VGND VGND VPWR VPWR D1[29] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_33_CLK clkbuf_6_5__f_CLK/X VGND VGND VPWR VPWR _34593_/CLK sky130_fd_sc_hd__clkbuf_16
Xoutput122 _31997_/Q VGND VGND VPWR VPWR D1[39] sky130_fd_sc_hd__buf_2
X_22050_ _33405_/Q _33341_/Q _33277_/Q _33213_/Q _21727_/X _21728_/X VGND VGND VPWR
+ VPWR _22050_/X sky130_fd_sc_hd__mux4_1
Xoutput133 _32007_/Q VGND VGND VPWR VPWR D1[49] sky130_fd_sc_hd__buf_2
XFILLER_217_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31248_ _27788_/X _35845_/Q _31252_/S VGND VGND VPWR VPWR _31249_/A sky130_fd_sc_hd__mux2_1
X_34036_ _34166_/CLK _34036_/D VGND VGND VPWR VPWR _34036_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput144 _32017_/Q VGND VGND VPWR VPWR D1[59] sky130_fd_sc_hd__buf_2
Xoutput155 _36192_/Q VGND VGND VPWR VPWR D2[10] sky130_fd_sc_hd__buf_2
XFILLER_138_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput166 _36202_/Q VGND VGND VPWR VPWR D2[20] sky130_fd_sc_hd__buf_2
X_21001_ _20997_/X _21000_/X _20644_/X _20646_/X VGND VGND VPWR VPWR _21016_/B sky130_fd_sc_hd__o211a_1
Xoutput177 _36212_/Q VGND VGND VPWR VPWR D2[30] sky130_fd_sc_hd__buf_2
XFILLER_82_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput188 _36222_/Q VGND VGND VPWR VPWR D2[40] sky130_fd_sc_hd__buf_2
XTAP_5809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31179_ _27686_/X _35812_/Q _31189_/S VGND VGND VPWR VPWR _31180_/A sky130_fd_sc_hd__mux2_1
Xoutput199 _36232_/Q VGND VGND VPWR VPWR D2[50] sky130_fd_sc_hd__buf_2
XFILLER_141_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35987_ _36051_/CLK _35987_/D VGND VGND VPWR VPWR _35987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25740_ _25740_/A VGND VGND VPWR VPWR _33331_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_214_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34938_ _36154_/CLK _34938_/D VGND VGND VPWR VPWR _34938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22952_ _22952_/A VGND VGND VPWR VPWR _32042_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21903_ _33657_/Q _33593_/Q _33529_/Q _33465_/Q _21800_/X _21801_/X VGND VGND VPWR
+ VPWR _21903_/X sky130_fd_sc_hd__mux4_1
XFILLER_244_846 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25671_ _24988_/X _33299_/Q _25675_/S VGND VGND VPWR VPWR _25672_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22883_ input83/X input89/X VGND VGND VPWR VPWR _28786_/A sky130_fd_sc_hd__nand2_4
X_34869_ _35126_/CLK _34869_/D VGND VGND VPWR VPWR _34869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_216_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27410_ _34089_/Q _27093_/X _27410_/S VGND VGND VPWR VPWR _27411_/A sky130_fd_sc_hd__mux2_1
X_24622_ _23027_/X _32835_/Q _24630_/S VGND VGND VPWR VPWR _24623_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28390_ _27655_/X _34522_/Q _28400_/S VGND VGND VPWR VPWR _28391_/A sky130_fd_sc_hd__mux2_1
X_21834_ _21828_/X _21833_/X _21765_/X VGND VGND VPWR VPWR _21835_/D sky130_fd_sc_hd__o21ba_1
XFILLER_243_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27341_ _34056_/Q _27189_/X _27359_/S VGND VGND VPWR VPWR _27342_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24553_ _22925_/X _32802_/Q _24567_/S VGND VGND VPWR VPWR _24554_/A sky130_fd_sc_hd__mux2_1
X_21765_ _22471_/A VGND VGND VPWR VPWR _21765_/X sky130_fd_sc_hd__buf_2
XFILLER_51_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23504_ _23504_/A VGND VGND VPWR VPWR _32247_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20716_ _20710_/X _20715_/X _20615_/X VGND VGND VPWR VPWR _20738_/A sky130_fd_sc_hd__o21ba_1
XFILLER_180_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27272_ _27272_/A VGND VGND VPWR VPWR _34023_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24484_ _24484_/A VGND VGND VPWR VPWR _32769_/D sky130_fd_sc_hd__clkbuf_1
X_21696_ _21446_/X _21692_/X _21695_/X _21451_/X VGND VGND VPWR VPWR _21696_/X sky130_fd_sc_hd__a22o_1
X_29011_ _34815_/Q _27162_/X _29027_/S VGND VGND VPWR VPWR _29012_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26223_ _24806_/X _33560_/Q _26237_/S VGND VGND VPWR VPWR _26224_/A sky130_fd_sc_hd__mux2_1
X_23435_ input39/X VGND VGND VPWR VPWR _23435_/X sky130_fd_sc_hd__buf_4
X_20647_ _20628_/X _20642_/X _20644_/X _20646_/X VGND VGND VPWR VPWR _20706_/B sky130_fd_sc_hd__o211a_1
XFILLER_109_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26154_ _26154_/A VGND VGND VPWR VPWR _33527_/D sky130_fd_sc_hd__clkbuf_1
X_20578_ _20578_/A VGND VGND VPWR VPWR _32469_/D sky130_fd_sc_hd__clkbuf_4
X_23366_ _23366_/A VGND VGND VPWR VPWR _32198_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_3_0_CLK clkbuf_0_CLK/X VGND VGND VPWR VPWR clkbuf_2_3_0_CLK/X sky130_fd_sc_hd__clkbuf_8
X_25105_ _25105_/A VGND VGND VPWR VPWR _33032_/D sky130_fd_sc_hd__clkbuf_1
X_22317_ _22317_/A VGND VGND VPWR VPWR _22317_/X sky130_fd_sc_hd__buf_4
XFILLER_165_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26085_ _26085_/A VGND VGND VPWR VPWR _33494_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23297_ _32171_/Q _23296_/X _23424_/S VGND VGND VPWR VPWR _23298_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_24_CLK clkbuf_6_5__f_CLK/X VGND VGND VPWR VPWR _36197_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_124_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29913_ _29913_/A VGND VGND VPWR VPWR _35212_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25036_ _24855_/X _33000_/Q _25038_/S VGND VGND VPWR VPWR _25037_/A sky130_fd_sc_hd__mux2_1
X_22248_ _35202_/Q _35138_/Q _35074_/Q _32258_/Q _21963_/X _21964_/X VGND VGND VPWR
+ VPWR _22248_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1051 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22179_ _34688_/Q _34624_/Q _34560_/Q _34496_/Q _21892_/X _21893_/X VGND VGND VPWR
+ VPWR _22179_/X sky130_fd_sc_hd__mux4_1
X_29844_ _29844_/A VGND VGND VPWR VPWR _35179_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29775_ _35147_/Q _29494_/X _29787_/S VGND VGND VPWR VPWR _29776_/A sky130_fd_sc_hd__mux2_1
X_26987_ _26987_/A VGND VGND VPWR VPWR _33919_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16740_ _17960_/A VGND VGND VPWR VPWR _16740_/X sky130_fd_sc_hd__buf_4
X_25938_ _25938_/A VGND VGND VPWR VPWR _33425_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28726_ _34681_/Q _27143_/X _28734_/S VGND VGND VPWR VPWR _28727_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28657_ _34648_/Q _27041_/X _28671_/S VGND VGND VPWR VPWR _28658_/A sky130_fd_sc_hd__mux2_1
X_16671_ _17850_/A VGND VGND VPWR VPWR _16671_/X sky130_fd_sc_hd__buf_4
X_25869_ _25869_/A VGND VGND VPWR VPWR _33392_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18410_ _18281_/X _18408_/X _18409_/X _18291_/X VGND VGND VPWR VPWR _18410_/X sky130_fd_sc_hd__a22o_1
XFILLER_28_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27608_ _34183_/Q _27186_/X _27608_/S VGND VGND VPWR VPWR _27609_/A sky130_fd_sc_hd__mux2_1
X_19390_ _19390_/A _19390_/B _19390_/C _19390_/D VGND VGND VPWR VPWR _19391_/A sky130_fd_sc_hd__or4_4
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28588_ _27748_/X _34616_/Q _28598_/S VGND VGND VPWR VPWR _28589_/A sky130_fd_sc_hd__mux2_1
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_912 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18341_ _20215_/A VGND VGND VPWR VPWR _18341_/X sky130_fd_sc_hd__buf_4
XFILLER_43_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27539_ _34150_/Q _27084_/X _27545_/S VGND VGND VPWR VPWR _27540_/A sky130_fd_sc_hd__mux2_1
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_995 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18272_ _16048_/X _18270_/X _18271_/X _16058_/X VGND VGND VPWR VPWR _18272_/X sky130_fd_sc_hd__a22o_1
XFILLER_202_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_967 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30550_ _30550_/A VGND VGND VPWR VPWR _35514_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_203_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17223_ _33078_/Q _32054_/Q _35830_/Q _35766_/Q _17078_/X _17079_/X VGND VGND VPWR
+ VPWR _17223_/X sky130_fd_sc_hd__mux4_1
X_29209_ _34909_/Q _27056_/X _29213_/S VGND VGND VPWR VPWR _29210_/A sky130_fd_sc_hd__mux2_1
X_30481_ _30481_/A VGND VGND VPWR VPWR _35481_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput13 DW[20] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__buf_6
X_32220_ _35187_/CLK _32220_/D VGND VGND VPWR VPWR _32220_/Q sky130_fd_sc_hd__dfxtp_1
Xinput24 DW[30] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__clkbuf_4
X_17154_ _34676_/Q _34612_/Q _34548_/Q _34484_/Q _16939_/X _16940_/X VGND VGND VPWR
+ VPWR _17154_/X sky130_fd_sc_hd__mux4_1
XFILLER_7_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput35 DW[40] VGND VGND VPWR VPWR input35/X sky130_fd_sc_hd__buf_6
Xinput46 DW[50] VGND VGND VPWR VPWR input46/X sky130_fd_sc_hd__buf_8
XFILLER_200_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput57 DW[60] VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__buf_8
Xinput68 R1[3] VGND VGND VPWR VPWR input68/X sky130_fd_sc_hd__clkbuf_8
X_16105_ _16089_/X _16102_/X _16104_/X VGND VGND VPWR VPWR _16106_/D sky130_fd_sc_hd__o21ba_1
XFILLER_7_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32151_ _35160_/CLK _32151_/D VGND VGND VPWR VPWR _32151_/Q sky130_fd_sc_hd__dfxtp_1
Xinput79 R3[2] VGND VGND VPWR VPWR input79/X sky130_fd_sc_hd__buf_4
X_17085_ _16800_/X _17083_/X _17084_/X _16803_/X VGND VGND VPWR VPWR _17085_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_15_CLK clkbuf_6_6__f_CLK/X VGND VGND VPWR VPWR _35684_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_170_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31102_ _35776_/Q input37/X _31116_/S VGND VGND VPWR VPWR _31103_/A sky130_fd_sc_hd__mux2_1
X_16036_ _16061_/A VGND VGND VPWR VPWR _17833_/A sky130_fd_sc_hd__buf_12
XFILLER_48_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32082_ _35858_/CLK _32082_/D VGND VGND VPWR VPWR _32082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31033_ _31033_/A VGND VGND VPWR VPWR _35743_/D sky130_fd_sc_hd__clkbuf_1
X_35910_ _35973_/CLK _35910_/D VGND VGND VPWR VPWR _35910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35841_ _35841_/CLK _35841_/D VGND VGND VPWR VPWR _35841_/Q sky130_fd_sc_hd__dfxtp_1
X_17987_ _32140_/Q _32332_/Q _32396_/Q _35916_/Q _17986_/X _17774_/X VGND VGND VPWR
+ VPWR _17987_/X sky130_fd_sc_hd__mux4_1
XFILLER_42_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19726_ _19719_/X _19725_/X _19440_/X _19441_/X VGND VGND VPWR VPWR _19743_/B sky130_fd_sc_hd__o211a_1
XFILLER_111_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16938_ _16934_/X _16937_/X _16798_/X VGND VGND VPWR VPWR _16948_/C sky130_fd_sc_hd__o21ba_1
X_35772_ _36029_/CLK _35772_/D VGND VGND VPWR VPWR _35772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32984_ _35992_/CLK _32984_/D VGND VGND VPWR VPWR _32984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1076 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34723_ _34914_/CLK _34723_/D VGND VGND VPWR VPWR _34723_/Q sky130_fd_sc_hd__dfxtp_1
X_31935_ _31935_/A VGND VGND VPWR VPWR _36170_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_1106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19657_ _35450_/Q _35386_/Q _35322_/Q _35258_/Q _19554_/X _19555_/X VGND VGND VPWR
+ VPWR _19657_/X sky130_fd_sc_hd__mux4_1
X_16869_ _35436_/Q _35372_/Q _35308_/Q _35244_/Q _16548_/X _16549_/X VGND VGND VPWR
+ VPWR _16869_/X sky130_fd_sc_hd__mux4_1
XFILLER_246_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18608_ _34396_/Q _36124_/Q _34268_/Q _34204_/Q _18470_/X _18471_/X VGND VGND VPWR
+ VPWR _18608_/X sky130_fd_sc_hd__mux4_1
XFILLER_168_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34654_ _34654_/CLK _34654_/D VGND VGND VPWR VPWR _34654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19588_ _35448_/Q _35384_/Q _35320_/Q _35256_/Q _19554_/X _19555_/X VGND VGND VPWR
+ VPWR _19588_/X sky130_fd_sc_hd__mux4_1
X_31866_ _31956_/S VGND VGND VPWR VPWR _31885_/S sky130_fd_sc_hd__buf_4
XFILLER_241_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33605_ _34179_/CLK _33605_/D VGND VGND VPWR VPWR _33605_/Q sky130_fd_sc_hd__dfxtp_1
X_18539_ _34906_/Q _34842_/Q _34778_/Q _34714_/Q _18396_/X _18398_/X VGND VGND VPWR
+ VPWR _18539_/X sky130_fd_sc_hd__mux4_1
X_30817_ _35641_/Q input29/X _30825_/S VGND VGND VPWR VPWR _30818_/A sky130_fd_sc_hd__mux2_1
X_34585_ _34585_/CLK _34585_/D VGND VGND VPWR VPWR _34585_/Q sky130_fd_sc_hd__dfxtp_1
X_31797_ _36105_/Q input47/X _31813_/S VGND VGND VPWR VPWR _31798_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33536_ _33984_/CLK _33536_/D VGND VGND VPWR VPWR _33536_/Q sky130_fd_sc_hd__dfxtp_1
X_21550_ _33647_/Q _33583_/Q _33519_/Q _33455_/Q _21447_/X _21448_/X VGND VGND VPWR
+ VPWR _21550_/X sky130_fd_sc_hd__mux4_1
X_30748_ _35608_/Q input23/X _30762_/S VGND VGND VPWR VPWR _30749_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20501_ _19458_/A _20499_/X _20500_/X _19463_/A VGND VGND VPWR VPWR _20501_/X sky130_fd_sc_hd__a22o_1
X_21481_ _21475_/X _21480_/X _21412_/X VGND VGND VPWR VPWR _21482_/D sky130_fd_sc_hd__o21ba_1
X_33467_ _34172_/CLK _33467_/D VGND VGND VPWR VPWR _33467_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30679_ _30679_/A VGND VGND VPWR VPWR _35575_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20432_ _33425_/Q _33361_/Q _33297_/Q _33233_/Q _20133_/X _20134_/X VGND VGND VPWR
+ VPWR _20432_/X sky130_fd_sc_hd__mux4_2
X_35206_ _35718_/CLK _35206_/D VGND VGND VPWR VPWR _35206_/Q sky130_fd_sc_hd__dfxtp_1
X_23220_ _23220_/A VGND VGND VPWR VPWR _32147_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32418_ _33573_/CLK _32418_/D VGND VGND VPWR VPWR _32418_/Q sky130_fd_sc_hd__dfxtp_1
X_36186_ _36191_/CLK _36186_/D VGND VGND VPWR VPWR _36186_/Q sky130_fd_sc_hd__dfxtp_1
X_33398_ _36087_/CLK _33398_/D VGND VGND VPWR VPWR _33398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20363_ _34446_/Q _36174_/Q _34318_/Q _34254_/Q _20235_/X _20236_/X VGND VGND VPWR
+ VPWR _20363_/X sky130_fd_sc_hd__mux4_1
X_35137_ _35715_/CLK _35137_/D VGND VGND VPWR VPWR _35137_/Q sky130_fd_sc_hd__dfxtp_1
X_23151_ _23151_/A VGND VGND VPWR VPWR _32114_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_834 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32349_ _32797_/CLK _32349_/D VGND VGND VPWR VPWR _32349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22102_ _33086_/Q _32062_/Q _35838_/Q _35774_/Q _22031_/X _22032_/X VGND VGND VPWR
+ VPWR _22102_/X sky130_fd_sc_hd__mux4_1
XTAP_7019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23082_ input60/X VGND VGND VPWR VPWR _23082_/X sky130_fd_sc_hd__buf_2
X_20294_ _35468_/Q _35404_/Q _35340_/Q _35276_/Q _20260_/X _20261_/X VGND VGND VPWR
+ VPWR _20294_/X sky130_fd_sc_hd__mux4_1
XFILLER_162_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35068_ _35581_/CLK _35068_/D VGND VGND VPWR VPWR _35068_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_6_31__f_CLK clkbuf_5_15_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_31__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XTAP_6318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26910_ _33883_/Q _23246_/X _26918_/S VGND VGND VPWR VPWR _26911_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22033_ _33084_/Q _32060_/Q _35836_/Q _35772_/Q _22031_/X _22032_/X VGND VGND VPWR
+ VPWR _22033_/X sky130_fd_sc_hd__mux4_1
XTAP_6329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34019_ _34148_/CLK _34019_/D VGND VGND VPWR VPWR _34019_/Q sky130_fd_sc_hd__dfxtp_1
X_27890_ _27714_/X _34285_/Q _27902_/S VGND VGND VPWR VPWR _27891_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26841_ _26841_/A VGND VGND VPWR VPWR _33850_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29560_ _35045_/Q _29376_/X _29568_/S VGND VGND VPWR VPWR _29561_/A sky130_fd_sc_hd__mux2_1
XFILLER_229_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26772_ _26772_/A VGND VGND VPWR VPWR _33817_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23984_ _22891_/X _32535_/Q _24000_/S VGND VGND VPWR VPWR _23985_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28511_ _27834_/X _34580_/Q _28513_/S VGND VGND VPWR VPWR _28512_/A sky130_fd_sc_hd__mux2_1
X_25723_ _24865_/X _33323_/Q _25739_/S VGND VGND VPWR VPWR _25724_/A sky130_fd_sc_hd__mux2_1
X_29491_ input48/X VGND VGND VPWR VPWR _29491_/X sky130_fd_sc_hd__buf_2
X_22935_ _22934_/X _32037_/Q _22947_/S VGND VGND VPWR VPWR _22936_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28442_ _27732_/X _34547_/Q _28442_/S VGND VGND VPWR VPWR _28443_/A sky130_fd_sc_hd__mux2_1
X_25654_ _25654_/A VGND VGND VPWR VPWR _33290_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_204_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22866_ _35477_/Q _35413_/Q _35349_/Q _35285_/Q _20609_/X _20611_/X VGND VGND VPWR
+ VPWR _22866_/X sky130_fd_sc_hd__mux4_1
XFILLER_232_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_231_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24605_ _23002_/X _32827_/Q _24609_/S VGND VGND VPWR VPWR _24606_/A sky130_fd_sc_hd__mux2_1
XFILLER_231_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28373_ _28373_/A VGND VGND VPWR VPWR _34514_/D sky130_fd_sc_hd__clkbuf_1
XPHY_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21817_ _21667_/X _21815_/X _21816_/X _21671_/X VGND VGND VPWR VPWR _21817_/X sky130_fd_sc_hd__a22o_1
XPHY_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25585_ _25675_/S VGND VGND VPWR VPWR _25604_/S sky130_fd_sc_hd__buf_4
X_22797_ _33171_/Q _36051_/Q _33043_/Q _32979_/Q _20632_/X _21761_/A VGND VGND VPWR
+ VPWR _22797_/X sky130_fd_sc_hd__mux4_1
XPHY_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27324_ _34048_/Q _27165_/X _27338_/S VGND VGND VPWR VPWR _27325_/A sky130_fd_sc_hd__mux2_1
XPHY_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24536_ _22900_/X _32794_/Q _24546_/S VGND VGND VPWR VPWR _24537_/A sky130_fd_sc_hd__mux2_1
XPHY_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21748_ _35444_/Q _35380_/Q _35316_/Q _35252_/Q _21501_/X _21502_/X VGND VGND VPWR
+ VPWR _21748_/X sky130_fd_sc_hd__mux4_1
XPHY_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27255_ _27255_/A VGND VGND VPWR VPWR _34015_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24467_ _24467_/A VGND VGND VPWR VPWR _32761_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21679_ _22536_/A VGND VGND VPWR VPWR _21679_/X sky130_fd_sc_hd__clkbuf_8
X_26206_ _26206_/A VGND VGND VPWR VPWR _33552_/D sky130_fd_sc_hd__clkbuf_1
X_23418_ _32218_/Q _23417_/X _23418_/S VGND VGND VPWR VPWR _23419_/A sky130_fd_sc_hd__mux2_1
X_27186_ input44/X VGND VGND VPWR VPWR _27186_/X sky130_fd_sc_hd__buf_4
XFILLER_149_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24398_ _24398_/A VGND VGND VPWR VPWR _32728_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26137_ _26137_/A VGND VGND VPWR VPWR _33519_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23349_ _32191_/Q _23274_/X _23359_/S VGND VGND VPWR VPWR _23350_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26068_ _24976_/X _33487_/Q _26072_/S VGND VGND VPWR VPWR _26069_/A sky130_fd_sc_hd__mux2_1
XFILLER_238_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17910_ _17910_/A VGND VGND VPWR VPWR _17910_/X sky130_fd_sc_hd__buf_4
XFILLER_180_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25019_ _25130_/S VGND VGND VPWR VPWR _25038_/S sky130_fd_sc_hd__buf_4
XFILLER_238_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_1324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18890_ _18747_/X _18888_/X _18889_/X _18750_/X VGND VGND VPWR VPWR _18890_/X sky130_fd_sc_hd__a22o_1
XTAP_6830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17841_ _33160_/Q _36040_/Q _33032_/Q _32968_/Q _17768_/X _17769_/X VGND VGND VPWR
+ VPWR _17841_/X sky130_fd_sc_hd__mux4_1
X_29827_ _29827_/A VGND VGND VPWR VPWR _35171_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_226_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29758_ _35139_/Q _29469_/X _29766_/S VGND VGND VPWR VPWR _29759_/A sky130_fd_sc_hd__mux2_1
X_17772_ _17765_/X _17767_/X _17770_/X _17771_/X VGND VGND VPWR VPWR _17772_/X sky130_fd_sc_hd__a22o_1
XFILLER_93_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19511_ _19505_/X _19510_/X _19432_/X VGND VGND VPWR VPWR _19535_/A sky130_fd_sc_hd__o21ba_1
X_16723_ _16645_/X _16721_/X _16722_/X _16648_/X VGND VGND VPWR VPWR _16723_/X sky130_fd_sc_hd__a22o_1
X_28709_ _34673_/Q _27118_/X _28713_/S VGND VGND VPWR VPWR _28710_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29689_ _35106_/Q _29367_/X _29703_/S VGND VGND VPWR VPWR _29690_/A sky130_fd_sc_hd__mux2_1
XFILLER_207_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_223_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31720_ _31720_/A VGND VGND VPWR VPWR _36068_/D sky130_fd_sc_hd__clkbuf_1
X_16654_ _16650_/X _16651_/X _16652_/X _16653_/X VGND VGND VPWR VPWR _16654_/X sky130_fd_sc_hd__a22o_1
X_19442_ _19436_/X _19439_/X _19440_/X _19441_/X VGND VGND VPWR VPWR _19467_/B sky130_fd_sc_hd__o211a_1
XFILLER_207_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_4_CLK clkbuf_leaf_9_CLK/A VGND VGND VPWR VPWR _34790_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_234_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31651_ _27785_/X _36036_/Q _31657_/S VGND VGND VPWR VPWR _31652_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16585_ _16581_/X _16584_/X _16445_/X VGND VGND VPWR VPWR _16595_/C sky130_fd_sc_hd__o21ba_1
X_19373_ _19366_/X _19372_/X _19087_/X _19088_/X VGND VGND VPWR VPWR _19390_/B sky130_fd_sc_hd__o211a_1
XFILLER_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_1475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18324_ _20206_/A VGND VGND VPWR VPWR _18324_/X sky130_fd_sc_hd__clkbuf_8
X_30602_ _30602_/A VGND VGND VPWR VPWR _35539_/D sky130_fd_sc_hd__clkbuf_1
X_34370_ _35715_/CLK _34370_/D VGND VGND VPWR VPWR _34370_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31582_ _27683_/X _36003_/Q _31594_/S VGND VGND VPWR VPWR _31583_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18255_ _18251_/X _18254_/X _17838_/A VGND VGND VPWR VPWR _18277_/A sky130_fd_sc_hd__o21ba_1
XFILLER_188_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33321_ _35622_/CLK _33321_/D VGND VGND VPWR VPWR _33321_/Q sky130_fd_sc_hd__dfxtp_1
X_30533_ _30533_/A VGND VGND VPWR VPWR _35506_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17206_ _17912_/A VGND VGND VPWR VPWR _17206_/X sky130_fd_sc_hd__buf_6
X_36040_ _36040_/CLK _36040_/D VGND VGND VPWR VPWR _36040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18186_ _18182_/X _18185_/X _17871_/A VGND VGND VPWR VPWR _18187_/D sky130_fd_sc_hd__o21ba_1
X_30464_ _35474_/Q _29515_/X _30470_/S VGND VGND VPWR VPWR _30465_/A sky130_fd_sc_hd__mux2_1
X_33252_ _33828_/CLK _33252_/D VGND VGND VPWR VPWR _33252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32203_ _35439_/CLK _32203_/D VGND VGND VPWR VPWR _32203_/Q sky130_fd_sc_hd__dfxtp_1
X_17137_ _32116_/Q _32308_/Q _32372_/Q _35892_/Q _16927_/X _17068_/X VGND VGND VPWR
+ VPWR _17137_/X sky130_fd_sc_hd__mux4_1
X_33183_ _35551_/CLK _33183_/D VGND VGND VPWR VPWR _33183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30395_ _35441_/Q _29413_/X _30399_/S VGND VGND VPWR VPWR _30396_/A sky130_fd_sc_hd__mux2_1
X_32134_ _35974_/CLK _32134_/D VGND VGND VPWR VPWR _32134_/Q sky130_fd_sc_hd__dfxtp_1
X_17068_ _17774_/A VGND VGND VPWR VPWR _17068_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_170_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16019_ _16061_/A VGND VGND VPWR VPWR _17982_/A sky130_fd_sc_hd__buf_12
X_32065_ _36034_/CLK _32065_/D VGND VGND VPWR VPWR _32065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31016_ _35735_/Q input12/X _31032_/S VGND VGND VPWR VPWR _31017_/A sky130_fd_sc_hd__mux2_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35824_ _36144_/CLK _35824_/D VGND VGND VPWR VPWR _35824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19709_ _33916_/Q _33852_/Q _33788_/Q _36092_/Q _19677_/X _19678_/X VGND VGND VPWR
+ VPWR _19709_/X sky130_fd_sc_hd__mux4_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35755_ _35755_/CLK _35755_/D VGND VGND VPWR VPWR _35755_/Q sky130_fd_sc_hd__dfxtp_1
X_20981_ _34910_/Q _34846_/Q _34782_/Q _34718_/Q _20696_/X _20698_/X VGND VGND VPWR
+ VPWR _20981_/X sky130_fd_sc_hd__mux4_1
X_32967_ _33160_/CLK _32967_/D VGND VGND VPWR VPWR _32967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22720_ _34704_/Q _34640_/Q _34576_/Q _34512_/Q _22598_/X _22599_/X VGND VGND VPWR
+ VPWR _22720_/X sky130_fd_sc_hd__mux4_1
X_34706_ _36115_/CLK _34706_/D VGND VGND VPWR VPWR _34706_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31918_ _31918_/A VGND VGND VPWR VPWR _36162_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_225_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35686_ _35687_/CLK _35686_/D VGND VGND VPWR VPWR _35686_/Q sky130_fd_sc_hd__dfxtp_1
X_32898_ _35970_/CLK _32898_/D VGND VGND VPWR VPWR _32898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34637_ _35663_/CLK _34637_/D VGND VGND VPWR VPWR _34637_/Q sky130_fd_sc_hd__dfxtp_1
X_22651_ _22373_/X _22649_/X _22650_/X _22377_/X VGND VGND VPWR VPWR _22651_/X sky130_fd_sc_hd__a22o_1
XFILLER_213_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31849_ _31849_/A VGND VGND VPWR VPWR _36129_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21602_ _21598_/X _21599_/X _21600_/X _21601_/X VGND VGND VPWR VPWR _21602_/X sky130_fd_sc_hd__a22o_1
X_25370_ _33157_/Q _23444_/X _25374_/S VGND VGND VPWR VPWR _25371_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34568_ _35208_/CLK _34568_/D VGND VGND VPWR VPWR _34568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22582_ _22582_/A VGND VGND VPWR VPWR _22582_/X sky130_fd_sc_hd__buf_6
XFILLER_55_1256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24321_ _22980_/X _32692_/Q _24339_/S VGND VGND VPWR VPWR _24322_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33519_ _33902_/CLK _33519_/D VGND VGND VPWR VPWR _33519_/Q sky130_fd_sc_hd__dfxtp_1
X_21533_ _35630_/Q _34990_/Q _34350_/Q _33710_/Q _21391_/X _21392_/X VGND VGND VPWR
+ VPWR _21533_/X sky130_fd_sc_hd__mux4_1
XFILLER_107_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34499_ _34693_/CLK _34499_/D VGND VGND VPWR VPWR _34499_/Q sky130_fd_sc_hd__dfxtp_1
X_27040_ _27040_/A VGND VGND VPWR VPWR _33943_/D sky130_fd_sc_hd__clkbuf_1
X_36238_ _36242_/CLK _36238_/D VGND VGND VPWR VPWR _36238_/Q sky130_fd_sc_hd__dfxtp_1
X_24252_ _24252_/A VGND VGND VPWR VPWR _32661_/D sky130_fd_sc_hd__clkbuf_1
X_21464_ _21314_/X _21462_/X _21463_/X _21318_/X VGND VGND VPWR VPWR _21464_/X sky130_fd_sc_hd__a22o_1
XFILLER_135_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23203_ _23052_/X _32139_/Q _23215_/S VGND VGND VPWR VPWR _23204_/A sky130_fd_sc_hd__mux2_1
X_20415_ _18281_/X _20413_/X _20414_/X _18291_/X VGND VGND VPWR VPWR _20415_/X sky130_fd_sc_hd__a22o_1
X_36169_ _36169_/CLK _36169_/D VGND VGND VPWR VPWR _36169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21395_ _35434_/Q _35370_/Q _35306_/Q _35242_/Q _21148_/X _21149_/X VGND VGND VPWR
+ VPWR _21395_/X sky130_fd_sc_hd__mux4_1
X_24183_ _32628_/Q _23387_/X _24201_/S VGND VGND VPWR VPWR _24184_/A sky130_fd_sc_hd__mux2_1
XFILLER_209_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23134_ _22949_/X _32106_/Q _23152_/S VGND VGND VPWR VPWR _23135_/A sky130_fd_sc_hd__mux2_1
X_20346_ _32654_/Q _32590_/Q _32526_/Q _35982_/Q _20282_/X _20066_/X VGND VGND VPWR
+ VPWR _20346_/X sky130_fd_sc_hd__mux4_1
X_28991_ _28991_/A VGND VGND VPWR VPWR _34805_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20277_ _20205_/X _20275_/X _20276_/X _20210_/X VGND VGND VPWR VPWR _20277_/X sky130_fd_sc_hd__a22o_1
XTAP_6115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27942_ _27791_/X _34310_/Q _27944_/S VGND VGND VPWR VPWR _27943_/A sky130_fd_sc_hd__mux2_1
X_23065_ _23064_/X _32079_/Q _23071_/S VGND VGND VPWR VPWR _23066_/A sky130_fd_sc_hd__mux2_1
XTAP_6126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_248_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22016_ _22374_/A VGND VGND VPWR VPWR _22016_/X sky130_fd_sc_hd__buf_4
XTAP_6159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27873_ _27689_/X _34277_/Q _27881_/S VGND VGND VPWR VPWR _27874_/A sky130_fd_sc_hd__mux2_1
XTAP_5425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29612_ _29660_/S VGND VGND VPWR VPWR _29631_/S sky130_fd_sc_hd__buf_4
XTAP_4713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26824_ _26824_/A VGND VGND VPWR VPWR _33842_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_208_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26755_ _33810_/Q _23487_/X _26761_/S VGND VGND VPWR VPWR _26756_/A sky130_fd_sc_hd__mux2_1
X_29543_ _35037_/Q _29351_/X _29547_/S VGND VGND VPWR VPWR _29544_/A sky130_fd_sc_hd__mux2_1
XTAP_4768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23967_ _23067_/X _32528_/Q _23969_/S VGND VGND VPWR VPWR _23968_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25706_ _24840_/X _33315_/Q _25718_/S VGND VGND VPWR VPWR _25707_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22918_ input2/X VGND VGND VPWR VPWR _22918_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_244_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29474_ _29474_/A VGND VGND VPWR VPWR _35012_/D sky130_fd_sc_hd__clkbuf_1
X_26686_ _33777_/Q _23364_/X _26690_/S VGND VGND VPWR VPWR _26687_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23898_ _22965_/X _32495_/Q _23906_/S VGND VGND VPWR VPWR _23899_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25637_ _25637_/A VGND VGND VPWR VPWR _33282_/D sky130_fd_sc_hd__clkbuf_1
X_28425_ _28425_/A VGND VGND VPWR VPWR _34538_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22849_ _33685_/Q _33621_/Q _33557_/Q _33493_/Q _20624_/X _20625_/X VGND VGND VPWR
+ VPWR _22849_/X sky130_fd_sc_hd__mux4_1
XFILLER_44_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28356_ _27804_/X _34506_/Q _28370_/S VGND VGND VPWR VPWR _28357_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_1451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16370_ _16292_/X _16368_/X _16369_/X _16295_/X VGND VGND VPWR VPWR _16370_/X sky130_fd_sc_hd__a22o_1
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25568_ _25568_/A VGND VGND VPWR VPWR _33249_/D sky130_fd_sc_hd__clkbuf_1
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27307_ _34040_/Q _27140_/X _27317_/S VGND VGND VPWR VPWR _27308_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24519_ _24519_/A VGND VGND VPWR VPWR _32786_/D sky130_fd_sc_hd__clkbuf_1
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28287_ _28287_/A VGND VGND VPWR VPWR _34473_/D sky130_fd_sc_hd__clkbuf_1
X_25499_ _24933_/X _33217_/Q _25511_/S VGND VGND VPWR VPWR _25500_/A sky130_fd_sc_hd__mux2_1
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18040_ _34190_/Q _34126_/Q _34062_/Q _33998_/Q _17799_/X _17800_/X VGND VGND VPWR
+ VPWR _18040_/X sky130_fd_sc_hd__mux4_1
X_27238_ _34007_/Q _27038_/X _27254_/S VGND VGND VPWR VPWR _27239_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27169_ _33985_/Q _27168_/X _27187_/S VGND VGND VPWR VPWR _27170_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30180_ _35339_/Q _29494_/X _30192_/S VGND VGND VPWR VPWR _30181_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19991_ _33412_/Q _33348_/Q _33284_/Q _33220_/Q _19780_/X _19781_/X VGND VGND VPWR
+ VPWR _19991_/X sky130_fd_sc_hd__mux4_1
XFILLER_99_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18942_ _32870_/Q _32806_/Q _32742_/Q _32678_/Q _18940_/X _18941_/X VGND VGND VPWR
+ VPWR _18942_/X sky130_fd_sc_hd__mux4_1
XFILLER_45_1414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_1132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18873_ _18653_/X _18871_/X _18872_/X _18659_/X VGND VGND VPWR VPWR _18873_/X sky130_fd_sc_hd__a22o_1
XTAP_6660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17824_ _34439_/Q _36167_/Q _34311_/Q _34247_/Q _17582_/X _17583_/X VGND VGND VPWR
+ VPWR _17824_/X sky130_fd_sc_hd__mux4_1
X_33870_ _33934_/CLK _33870_/D VGND VGND VPWR VPWR _33870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_212_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32821_ _32903_/CLK _32821_/D VGND VGND VPWR VPWR _32821_/Q sky130_fd_sc_hd__dfxtp_1
X_17755_ _17751_/X _17754_/X _17518_/X VGND VGND VPWR VPWR _17756_/D sky130_fd_sc_hd__o21ba_1
XFILLER_78_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35540_ _35733_/CLK _35540_/D VGND VGND VPWR VPWR _35540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16706_ _17905_/A VGND VGND VPWR VPWR _16706_/X sky130_fd_sc_hd__clkbuf_4
X_32752_ _32879_/CLK _32752_/D VGND VGND VPWR VPWR _32752_/Q sky130_fd_sc_hd__dfxtp_1
X_17686_ _17686_/A _17686_/B _17686_/C _17686_/D VGND VGND VPWR VPWR _17687_/A sky130_fd_sc_hd__or4_1
XFILLER_208_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31703_ _31703_/A VGND VGND VPWR VPWR _36060_/D sky130_fd_sc_hd__clkbuf_1
X_19425_ _34164_/Q _34100_/Q _34036_/Q _33972_/Q _19393_/X _19394_/X VGND VGND VPWR
+ VPWR _19425_/X sky130_fd_sc_hd__mux4_1
X_35471_ _35471_/CLK _35471_/D VGND VGND VPWR VPWR _35471_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16637_ _33126_/Q _36006_/Q _32998_/Q _32934_/Q _16356_/X _16357_/X VGND VGND VPWR
+ VPWR _16637_/X sky130_fd_sc_hd__mux4_1
XFILLER_165_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32683_ _32875_/CLK _32683_/D VGND VGND VPWR VPWR _32683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34422_ _35126_/CLK _34422_/D VGND VGND VPWR VPWR _34422_/Q sky130_fd_sc_hd__dfxtp_1
X_19356_ _33906_/Q _33842_/Q _33778_/Q _36082_/Q _19324_/X _19325_/X VGND VGND VPWR
+ VPWR _19356_/X sky130_fd_sc_hd__mux4_1
X_31634_ _27760_/X _36028_/Q _31636_/S VGND VGND VPWR VPWR _31635_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16568_ _16500_/X _16566_/X _16567_/X _16503_/X VGND VGND VPWR VPWR _16568_/X sky130_fd_sc_hd__a22o_1
XFILLER_222_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18307_ _20215_/A VGND VGND VPWR VPWR _18307_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_52_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34353_ _35439_/CLK _34353_/D VGND VGND VPWR VPWR _34353_/Q sky130_fd_sc_hd__dfxtp_1
X_31565_ _27658_/X _35995_/Q _31573_/S VGND VGND VPWR VPWR _31566_/A sky130_fd_sc_hd__mux2_1
X_16499_ _16493_/X _16496_/X _16497_/X _16498_/X VGND VGND VPWR VPWR _16499_/X sky130_fd_sc_hd__a22o_1
X_19287_ _19153_/X _19285_/X _19286_/X _19156_/X VGND VGND VPWR VPWR _19287_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33304_ _36057_/CLK _33304_/D VGND VGND VPWR VPWR _33304_/Q sky130_fd_sc_hd__dfxtp_1
X_18238_ _16001_/X _18236_/X _18237_/X _16007_/X VGND VGND VPWR VPWR _18238_/X sky130_fd_sc_hd__a22o_1
XFILLER_30_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30516_ _35498_/Q _29391_/X _30534_/S VGND VGND VPWR VPWR _30517_/A sky130_fd_sc_hd__mux2_1
XFILLER_176_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34284_ _36140_/CLK _34284_/D VGND VGND VPWR VPWR _34284_/Q sky130_fd_sc_hd__dfxtp_1
X_31496_ _31496_/A VGND VGND VPWR VPWR _35962_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36023_ _36023_/CLK _36023_/D VGND VGND VPWR VPWR _36023_/Q sky130_fd_sc_hd__dfxtp_1
X_33235_ _36180_/CLK _33235_/D VGND VGND VPWR VPWR _33235_/Q sky130_fd_sc_hd__dfxtp_1
X_30447_ _30447_/A VGND VGND VPWR VPWR _35465_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18169_ _32146_/Q _32338_/Q _32402_/Q _35922_/Q _17986_/X _17011_/A VGND VGND VPWR
+ VPWR _18169_/X sky130_fd_sc_hd__mux4_1
XFILLER_11_1137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20200_ _34953_/Q _34889_/Q _34825_/Q _34761_/Q _20166_/X _20167_/X VGND VGND VPWR
+ VPWR _20200_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21180_ _35620_/Q _34980_/Q _34340_/Q _33700_/Q _21038_/X _21039_/X VGND VGND VPWR
+ VPWR _21180_/X sky130_fd_sc_hd__mux4_1
XFILLER_239_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33166_ _36045_/CLK _33166_/D VGND VGND VPWR VPWR _33166_/Q sky130_fd_sc_hd__dfxtp_1
X_30378_ _35433_/Q _29388_/X _30378_/S VGND VGND VPWR VPWR _30379_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_1298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20131_ _34184_/Q _34120_/Q _34056_/Q _33992_/Q _20099_/X _20100_/X VGND VGND VPWR
+ VPWR _20131_/X sky130_fd_sc_hd__mux4_1
XFILLER_143_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32117_ _32885_/CLK _32117_/D VGND VGND VPWR VPWR _32117_/Q sky130_fd_sc_hd__dfxtp_1
X_33097_ _35849_/CLK _33097_/D VGND VGND VPWR VPWR _33097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_217_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20062_ _33926_/Q _33862_/Q _33798_/Q _36102_/Q _20030_/X _20031_/X VGND VGND VPWR
+ VPWR _20062_/X sky130_fd_sc_hd__mux4_1
X_32048_ _36017_/CLK _32048_/D VGND VGND VPWR VPWR _32048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_217_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24870_ _24870_/A VGND VGND VPWR VPWR _32940_/D sky130_fd_sc_hd__clkbuf_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35807_ _35807_/CLK _35807_/D VGND VGND VPWR VPWR _35807_/Q sky130_fd_sc_hd__dfxtp_1
X_23821_ _23821_/A VGND VGND VPWR VPWR _32395_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33999_ _34192_/CLK _33999_/D VGND VGND VPWR VPWR _33999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26540_ _26540_/A VGND VGND VPWR VPWR _33709_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35738_ _35801_/CLK _35738_/D VGND VGND VPWR VPWR _35738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23752_ _23752_/A VGND VGND VPWR VPWR _32362_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_241_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20964_ _32862_/Q _32798_/Q _32734_/Q _32670_/Q _20887_/X _20888_/X VGND VGND VPWR
+ VPWR _20964_/X sky130_fd_sc_hd__mux4_1
XFILLER_26_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22703_ _33936_/Q _33872_/Q _33808_/Q _36112_/Q _20662_/X _20664_/X VGND VGND VPWR
+ VPWR _22703_/X sky130_fd_sc_hd__mux4_1
XFILLER_214_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26471_ _26471_/A VGND VGND VPWR VPWR _33677_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35669_ _35669_/CLK _35669_/D VGND VGND VPWR VPWR _35669_/Q sky130_fd_sc_hd__dfxtp_1
X_23683_ _23683_/A VGND VGND VPWR VPWR _32331_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20895_ _22462_/A VGND VGND VPWR VPWR _20895_/X sky130_fd_sc_hd__buf_4
XFILLER_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_246_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28210_ _27788_/X _34437_/Q _28214_/S VGND VGND VPWR VPWR _28211_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_1359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25422_ _25422_/A VGND VGND VPWR VPWR _33180_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29190_ _29190_/A VGND VGND VPWR VPWR _34900_/D sky130_fd_sc_hd__clkbuf_1
X_22634_ _34957_/Q _34893_/Q _34829_/Q _34765_/Q _22466_/X _22467_/X VGND VGND VPWR
+ VPWR _22634_/X sky130_fd_sc_hd__mux4_1
XFILLER_179_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28141_ _27686_/X _34404_/Q _28151_/S VGND VGND VPWR VPWR _28142_/A sky130_fd_sc_hd__mux2_1
X_25353_ _33149_/Q _23417_/X _25353_/S VGND VGND VPWR VPWR _25354_/A sky130_fd_sc_hd__mux2_1
X_22565_ _22559_/X _22564_/X _22457_/X VGND VGND VPWR VPWR _22573_/C sky130_fd_sc_hd__o21ba_1
XFILLER_16_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24304_ _22956_/X _32684_/Q _24318_/S VGND VGND VPWR VPWR _24305_/A sky130_fd_sc_hd__mux2_1
X_28072_ _28072_/A VGND VGND VPWR VPWR _34371_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21516_ _33646_/Q _33582_/Q _33518_/Q _33454_/Q _21447_/X _21448_/X VGND VGND VPWR
+ VPWR _21516_/X sky130_fd_sc_hd__mux4_1
X_25284_ _33116_/Q _23249_/X _25290_/S VGND VGND VPWR VPWR _25285_/A sky130_fd_sc_hd__mux2_1
X_22496_ _34697_/Q _34633_/Q _34569_/Q _34505_/Q _22245_/X _22246_/X VGND VGND VPWR
+ VPWR _22496_/X sky130_fd_sc_hd__mux4_1
XFILLER_222_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27023_ _33937_/Q _23484_/X _27023_/S VGND VGND VPWR VPWR _27024_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24235_ _32653_/Q _23472_/X _24243_/S VGND VGND VPWR VPWR _24236_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21447_ _22506_/A VGND VGND VPWR VPWR _21447_/X sky130_fd_sc_hd__buf_4
XFILLER_163_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24166_ _32620_/Q _23299_/X _24180_/S VGND VGND VPWR VPWR _24167_/A sky130_fd_sc_hd__mux2_1
X_21378_ _21100_/X _21376_/X _21377_/X _21103_/X VGND VGND VPWR VPWR _21378_/X sky130_fd_sc_hd__a22o_1
XFILLER_162_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23117_ _22925_/X _32098_/Q _23131_/S VGND VGND VPWR VPWR _23118_/A sky130_fd_sc_hd__mux2_1
XFILLER_218_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20329_ _20325_/X _20328_/X _20157_/X VGND VGND VPWR VPWR _20337_/C sky130_fd_sc_hd__o21ba_1
XFILLER_235_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24097_ _23058_/X _32589_/Q _24105_/S VGND VGND VPWR VPWR _24098_/A sky130_fd_sc_hd__mux2_1
X_28974_ _28974_/A VGND VGND VPWR VPWR _34797_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27925_ _27973_/S VGND VGND VPWR VPWR _27944_/S sky130_fd_sc_hd__buf_4
XTAP_5200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23048_ _23048_/A VGND VGND VPWR VPWR _32073_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27856_ _27664_/X _34269_/Q _27860_/S VGND VGND VPWR VPWR _27857_/A sky130_fd_sc_hd__mux2_1
XTAP_5255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26807_ _33834_/Q _23292_/X _26825_/S VGND VGND VPWR VPWR _26808_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_618 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27787_ _27787_/A VGND VGND VPWR VPWR _34244_/D sky130_fd_sc_hd__clkbuf_1
X_24999_ _24796_/X _32982_/Q _25017_/S VGND VGND VPWR VPWR _25000_/A sky130_fd_sc_hd__mux2_1
XTAP_4565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29526_ _29526_/A VGND VGND VPWR VPWR _35029_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17540_ _33087_/Q _32063_/Q _35839_/Q _35775_/Q _17431_/X _17432_/X VGND VGND VPWR
+ VPWR _17540_/X sky130_fd_sc_hd__mux4_1
XTAP_3853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26738_ _26738_/A VGND VGND VPWR VPWR _33801_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17471_ _34429_/Q _36157_/Q _34301_/Q _34237_/Q _17229_/X _17230_/X VGND VGND VPWR
+ VPWR _17471_/X sky130_fd_sc_hd__mux4_1
XFILLER_204_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29457_ input36/X VGND VGND VPWR VPWR _29457_/X sky130_fd_sc_hd__clkbuf_4
X_26669_ _33769_/Q _23289_/X _26669_/S VGND VGND VPWR VPWR _26670_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19210_ _34413_/Q _36141_/Q _34285_/Q _34221_/Q _19176_/X _19177_/X VGND VGND VPWR
+ VPWR _19210_/X sky130_fd_sc_hd__mux4_1
X_16422_ _17800_/A VGND VGND VPWR VPWR _16422_/X sky130_fd_sc_hd__buf_4
X_28408_ _28408_/A VGND VGND VPWR VPWR _34530_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29388_ input11/X VGND VGND VPWR VPWR _29388_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_220_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16353_ _17905_/A VGND VGND VPWR VPWR _16353_/X sky130_fd_sc_hd__buf_2
X_19141_ _34923_/Q _34859_/Q _34795_/Q _34731_/Q _19107_/X _19108_/X VGND VGND VPWR
+ VPWR _19141_/X sky130_fd_sc_hd__mux4_1
XFILLER_201_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28339_ _27779_/X _34498_/Q _28349_/S VGND VGND VPWR VPWR _28340_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19072_ _34154_/Q _34090_/Q _34026_/Q _33962_/Q _19040_/X _19041_/X VGND VGND VPWR
+ VPWR _19072_/X sky130_fd_sc_hd__mux4_1
X_31350_ _27739_/X _35893_/Q _31366_/S VGND VGND VPWR VPWR _31351_/A sky130_fd_sc_hd__mux2_1
X_16284_ _33116_/Q _35996_/Q _32988_/Q _32924_/Q _16024_/X _16025_/X VGND VGND VPWR
+ VPWR _16284_/X sky130_fd_sc_hd__mux4_1
XFILLER_125_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30301_ _30301_/A VGND VGND VPWR VPWR _35396_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_1191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18023_ _35725_/Q _32236_/Q _35597_/Q _35533_/Q _15993_/X _15995_/X VGND VGND VPWR
+ VPWR _18023_/X sky130_fd_sc_hd__mux4_1
XFILLER_199_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31281_ _27837_/X _35861_/Q _31281_/S VGND VGND VPWR VPWR _31282_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30232_ _30232_/A VGND VGND VPWR VPWR _35363_/D sky130_fd_sc_hd__clkbuf_1
X_33020_ _35451_/CLK _33020_/D VGND VGND VPWR VPWR _33020_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_236_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30163_ _35331_/Q _29469_/X _30171_/S VGND VGND VPWR VPWR _30164_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19974_ _19651_/X _19972_/X _19973_/X _19654_/X VGND VGND VPWR VPWR _19974_/X sky130_fd_sc_hd__a22o_1
XFILLER_125_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18925_ _18752_/X _18923_/X _18924_/X _18757_/X VGND VGND VPWR VPWR _18925_/X sky130_fd_sc_hd__a22o_1
XFILLER_84_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34971_ _35802_/CLK _34971_/D VGND VGND VPWR VPWR _34971_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30094_ _35298_/Q _29367_/X _30108_/S VGND VGND VPWR VPWR _30095_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_295_CLK clkbuf_6_56__f_CLK/X VGND VGND VPWR VPWR _36037_/CLK sky130_fd_sc_hd__clkbuf_16
X_33922_ _36099_/CLK _33922_/D VGND VGND VPWR VPWR _33922_/Q sky130_fd_sc_hd__dfxtp_1
X_18856_ _18747_/X _18854_/X _18855_/X _18750_/X VGND VGND VPWR VPWR _18856_/X sky130_fd_sc_hd__a22o_1
XFILLER_94_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17807_ _32647_/Q _32583_/Q _32519_/Q _35975_/Q _17629_/X _17766_/X VGND VGND VPWR
+ VPWR _17807_/X sky130_fd_sc_hd__mux4_1
XFILLER_209_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33853_ _36093_/CLK _33853_/D VGND VGND VPWR VPWR _33853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_927 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18787_ _34401_/Q _36129_/Q _34273_/Q _34209_/Q _18470_/X _18471_/X VGND VGND VPWR
+ VPWR _18787_/X sky130_fd_sc_hd__mux4_2
X_15999_ _15999_/A VGND VGND VPWR VPWR _17773_/A sky130_fd_sc_hd__buf_2
XFILLER_54_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32804_ _32804_/CLK _32804_/D VGND VGND VPWR VPWR _32804_/Q sky130_fd_sc_hd__dfxtp_1
X_17738_ _32133_/Q _32325_/Q _32389_/Q _35909_/Q _17633_/X _17421_/X VGND VGND VPWR
+ VPWR _17738_/X sky130_fd_sc_hd__mux4_1
X_33784_ _33911_/CLK _33784_/D VGND VGND VPWR VPWR _33784_/Q sky130_fd_sc_hd__dfxtp_1
X_30996_ _35726_/Q input52/X _31002_/S VGND VGND VPWR VPWR _30997_/A sky130_fd_sc_hd__mux2_1
XFILLER_235_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_247_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35523_ _35655_/CLK _35523_/D VGND VGND VPWR VPWR _35523_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32735_ _35870_/CLK _32735_/D VGND VGND VPWR VPWR _32735_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17669_ _17665_/X _17668_/X _17493_/X _17494_/X VGND VGND VPWR VPWR _17686_/B sky130_fd_sc_hd__o211a_1
X_19408_ _35699_/Q _32207_/Q _35571_/Q _35507_/Q _19264_/X _19265_/X VGND VGND VPWR
+ VPWR _19408_/X sky130_fd_sc_hd__mux4_1
X_35454_ _35454_/CLK _35454_/D VGND VGND VPWR VPWR _35454_/Q sky130_fd_sc_hd__dfxtp_1
X_20680_ _22536_/A VGND VGND VPWR VPWR _20680_/X sky130_fd_sc_hd__buf_6
X_32666_ _34070_/CLK _32666_/D VGND VGND VPWR VPWR _32666_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34405_ _34405_/CLK _34405_/D VGND VGND VPWR VPWR _34405_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19339_ _35441_/Q _35377_/Q _35313_/Q _35249_/Q _19201_/X _19202_/X VGND VGND VPWR
+ VPWR _19339_/X sky130_fd_sc_hd__mux4_1
X_31617_ _31686_/S VGND VGND VPWR VPWR _31636_/S sky130_fd_sc_hd__buf_4
XFILLER_143_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35385_ _35449_/CLK _35385_/D VGND VGND VPWR VPWR _35385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32597_ _35988_/CLK _32597_/D VGND VGND VPWR VPWR _32597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22350_ _35205_/Q _35141_/Q _35077_/Q _32261_/Q _22316_/X _22317_/X VGND VGND VPWR
+ VPWR _22350_/X sky130_fd_sc_hd__mux4_1
XFILLER_137_918 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34336_ _34913_/CLK _34336_/D VGND VGND VPWR VPWR _34336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31548_ _31548_/A VGND VGND VPWR VPWR _35987_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21301_ _21093_/X _21299_/X _21300_/X _21098_/X VGND VGND VPWR VPWR _21301_/X sky130_fd_sc_hd__a22o_1
XFILLER_108_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34267_ _36127_/CLK _34267_/D VGND VGND VPWR VPWR _34267_/Q sky130_fd_sc_hd__dfxtp_1
X_22281_ _22106_/X _22279_/X _22280_/X _22109_/X VGND VGND VPWR VPWR _22281_/X sky130_fd_sc_hd__a22o_1
XFILLER_163_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31479_ _31479_/A VGND VGND VPWR VPWR _35954_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24020_ _24020_/A VGND VGND VPWR VPWR _32552_/D sky130_fd_sc_hd__clkbuf_1
X_36006_ _36007_/CLK _36006_/D VGND VGND VPWR VPWR _36006_/Q sky130_fd_sc_hd__dfxtp_1
X_33218_ _36099_/CLK _33218_/D VGND VGND VPWR VPWR _33218_/Q sky130_fd_sc_hd__dfxtp_1
X_21232_ _33382_/Q _33318_/Q _33254_/Q _33190_/Q _21021_/X _21022_/X VGND VGND VPWR
+ VPWR _21232_/X sky130_fd_sc_hd__mux4_1
XFILLER_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34198_ _34647_/CLK _34198_/D VGND VGND VPWR VPWR _34198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_219_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21163_ _33636_/Q _33572_/Q _33508_/Q _33444_/Q _21094_/X _21095_/X VGND VGND VPWR
+ VPWR _21163_/X sky130_fd_sc_hd__mux4_1
XFILLER_46_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33149_ _35965_/CLK _33149_/D VGND VGND VPWR VPWR _33149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20114_ _35719_/Q _32229_/Q _35591_/Q _35527_/Q _19970_/X _19971_/X VGND VGND VPWR
+ VPWR _20114_/X sky130_fd_sc_hd__mux4_1
XFILLER_172_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25971_ _25971_/A VGND VGND VPWR VPWR _33440_/D sky130_fd_sc_hd__clkbuf_1
X_21094_ _22506_/A VGND VGND VPWR VPWR _21094_/X sky130_fd_sc_hd__buf_6
XFILLER_213_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_286_CLK clkbuf_6_58__f_CLK/X VGND VGND VPWR VPWR _35456_/CLK sky130_fd_sc_hd__clkbuf_16
X_20045_ _35461_/Q _35397_/Q _35333_/Q _35269_/Q _19907_/X _19908_/X VGND VGND VPWR
+ VPWR _20045_/X sky130_fd_sc_hd__mux4_1
XFILLER_150_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27710_ _27710_/A VGND VGND VPWR VPWR _34219_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24922_ _24922_/A VGND VGND VPWR VPWR _32957_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28690_ _34664_/Q _27090_/X _28692_/S VGND VGND VPWR VPWR _28691_/A sky130_fd_sc_hd__mux2_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27641_ _27641_/A VGND VGND VPWR VPWR _31823_/B sky130_fd_sc_hd__buf_12
XFILLER_150_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24853_ _24852_/X _32935_/Q _24859_/S VGND VGND VPWR VPWR _24854_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23804_ _23804_/A VGND VGND VPWR VPWR _32387_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27572_ _27572_/A VGND VGND VPWR VPWR _34165_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24784_ _23067_/X _32912_/Q _24786_/S VGND VGND VPWR VPWR _24785_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_1191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21996_ _34683_/Q _34619_/Q _34555_/Q _34491_/Q _21892_/X _21893_/X VGND VGND VPWR
+ VPWR _21996_/X sky130_fd_sc_hd__mux4_1
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29311_ _29311_/A VGND VGND VPWR VPWR _34957_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_214_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26523_ _26523_/A VGND VGND VPWR VPWR _33701_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23735_ _23735_/A VGND VGND VPWR VPWR _32354_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20947_ _34142_/Q _34078_/Q _34014_/Q _33950_/Q _20609_/X _20611_/X VGND VGND VPWR
+ VPWR _20947_/X sky130_fd_sc_hd__mux4_1
XFILLER_42_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26454_ _26454_/A VGND VGND VPWR VPWR _33669_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_230_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29242_ _29242_/A VGND VGND VPWR VPWR _34924_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23666_ _23666_/A VGND VGND VPWR VPWR _32323_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_947 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20878_ _20740_/X _20876_/X _20877_/X _20745_/X VGND VGND VPWR VPWR _20878_/X sky130_fd_sc_hd__a22o_1
XFILLER_202_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25405_ input87/X input86/X input88/X VGND VGND VPWR VPWR _25406_/A sky130_fd_sc_hd__and3b_1
X_29173_ _34892_/Q _27202_/X _29183_/S VGND VGND VPWR VPWR _29174_/A sky130_fd_sc_hd__mux2_1
X_22617_ _33165_/Q _36045_/Q _33037_/Q _32973_/Q _22368_/X _22369_/X VGND VGND VPWR
+ VPWR _22617_/X sky130_fd_sc_hd__mux4_1
X_26385_ _26385_/A VGND VGND VPWR VPWR _33636_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23597_ _23597_/A VGND VGND VPWR VPWR _32290_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28124_ _27661_/X _34396_/Q _28130_/S VGND VGND VPWR VPWR _28125_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_210_CLK clkbuf_6_52__f_CLK/X VGND VGND VPWR VPWR _35208_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_161_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25336_ _25336_/A VGND VGND VPWR VPWR _33140_/D sky130_fd_sc_hd__clkbuf_1
X_22548_ _22512_/X _22546_/X _22547_/X _22515_/X VGND VGND VPWR VPWR _22548_/X sky130_fd_sc_hd__a22o_1
XFILLER_224_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_9_0_CLK clkbuf_5_9_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_9_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_5_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28055_ _28055_/A VGND VGND VPWR VPWR _34363_/D sky130_fd_sc_hd__clkbuf_1
X_25267_ _33109_/Q _23498_/X _25267_/S VGND VGND VPWR VPWR _25268_/A sky130_fd_sc_hd__mux2_1
X_22479_ _33929_/Q _33865_/Q _33801_/Q _36105_/Q _22330_/X _22331_/X VGND VGND VPWR
+ VPWR _22479_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27006_ _27006_/A VGND VGND VPWR VPWR _33928_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24218_ _32645_/Q _23444_/X _24222_/S VGND VGND VPWR VPWR _24219_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25198_ _25267_/S VGND VGND VPWR VPWR _25217_/S sky130_fd_sc_hd__buf_8
XFILLER_108_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24149_ _32612_/Q _23274_/X _24159_/S VGND VGND VPWR VPWR _24150_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28957_ _28957_/A VGND VGND VPWR VPWR _34789_/D sky130_fd_sc_hd__clkbuf_1
X_16971_ _16650_/X _16969_/X _16970_/X _16653_/X VGND VGND VPWR VPWR _16971_/X sky130_fd_sc_hd__a22o_1
XFILLER_96_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_277_CLK clkbuf_6_59__f_CLK/X VGND VGND VPWR VPWR _36097_/CLK sky130_fd_sc_hd__clkbuf_16
X_18710_ _35167_/Q _35103_/Q _35039_/Q _32159_/Q _18604_/X _18605_/X VGND VGND VPWR
+ VPWR _18710_/X sky130_fd_sc_hd__mux4_1
XFILLER_81_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27908_ _27908_/A VGND VGND VPWR VPWR _34293_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19690_ _35643_/Q _35003_/Q _34363_/Q _33723_/Q _19444_/X _19445_/X VGND VGND VPWR
+ VPWR _19690_/X sky130_fd_sc_hd__mux4_1
XFILLER_103_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28888_ _34757_/Q _27180_/X _28892_/S VGND VGND VPWR VPWR _28889_/A sky130_fd_sc_hd__mux2_1
XTAP_5052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18641_ _34909_/Q _34845_/Q _34781_/Q _34717_/Q _18396_/X _18398_/X VGND VGND VPWR
+ VPWR _18641_/X sky130_fd_sc_hd__mux4_1
XTAP_5074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27839_ _27839_/A VGND VGND VPWR VPWR _34261_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18572_ _18391_/X _18570_/X _18571_/X _18401_/X VGND VGND VPWR VPWR _18572_/X sky130_fd_sc_hd__a22o_1
XFILLER_206_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30850_ _30850_/A VGND VGND VPWR VPWR _35656_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29509_ input54/X VGND VGND VPWR VPWR _29509_/X sky130_fd_sc_hd__buf_2
XTAP_3683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17523_ _34175_/Q _34111_/Q _34047_/Q _33983_/Q _17446_/X _17447_/X VGND VGND VPWR
+ VPWR _17523_/X sky130_fd_sc_hd__mux4_1
XFILLER_17_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30781_ _35624_/Q input10/X _30783_/S VGND VGND VPWR VPWR _30782_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32520_ _35975_/CLK _32520_/D VGND VGND VPWR VPWR _32520_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17454_ _32637_/Q _32573_/Q _32509_/Q _35965_/Q _17276_/X _17413_/X VGND VGND VPWR
+ VPWR _17454_/X sky130_fd_sc_hd__mux4_1
XFILLER_33_868 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_969 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16405_ _35423_/Q _35359_/Q _35295_/Q _35231_/Q _16195_/X _16196_/X VGND VGND VPWR
+ VPWR _16405_/X sky130_fd_sc_hd__mux4_1
X_32451_ _36076_/CLK _32451_/D VGND VGND VPWR VPWR _32451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17385_ _32123_/Q _32315_/Q _32379_/Q _35899_/Q _17280_/X _17068_/X VGND VGND VPWR
+ VPWR _17385_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_201_CLK clkbuf_6_49__f_CLK/X VGND VGND VPWR VPWR _35785_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_13_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31402_ _27816_/X _35918_/Q _31408_/S VGND VGND VPWR VPWR _31403_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19124_ _33131_/Q _36011_/Q _33003_/Q _32939_/Q _19009_/X _19010_/X VGND VGND VPWR
+ VPWR _19124_/X sky130_fd_sc_hd__mux4_1
XFILLER_158_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16336_ _16332_/X _16335_/X _16075_/X VGND VGND VPWR VPWR _16344_/C sky130_fd_sc_hd__o21ba_1
X_35170_ _36197_/CLK _35170_/D VGND VGND VPWR VPWR _35170_/Q sky130_fd_sc_hd__dfxtp_1
X_32382_ _32895_/CLK _32382_/D VGND VGND VPWR VPWR _32382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34121_ _34121_/CLK _34121_/D VGND VGND VPWR VPWR _34121_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16267_ _34651_/Q _34587_/Q _34523_/Q _34459_/Q _16233_/X _16234_/X VGND VGND VPWR
+ VPWR _16267_/X sky130_fd_sc_hd__mux4_1
X_19055_ _35689_/Q _32196_/Q _35561_/Q _35497_/Q _18911_/X _18912_/X VGND VGND VPWR
+ VPWR _19055_/X sky130_fd_sc_hd__mux4_1
X_31333_ _27714_/X _35885_/Q _31345_/S VGND VGND VPWR VPWR _31334_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18006_ _18002_/X _18005_/X _17871_/X VGND VGND VPWR VPWR _18007_/D sky130_fd_sc_hd__o21ba_1
XFILLER_195_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34052_ _34180_/CLK _34052_/D VGND VGND VPWR VPWR _34052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16198_ _33049_/Q _32025_/Q _35801_/Q _35737_/Q _16067_/X _16069_/X VGND VGND VPWR
+ VPWR _16198_/X sky130_fd_sc_hd__mux4_1
XFILLER_160_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31264_ _31264_/A VGND VGND VPWR VPWR _35852_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33003_ _35820_/CLK _33003_/D VGND VGND VPWR VPWR _33003_/Q sky130_fd_sc_hd__dfxtp_1
X_30215_ _30215_/A VGND VGND VPWR VPWR _35355_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_236_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31195_ _31195_/A VGND VGND VPWR VPWR _35819_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30146_ _35323_/Q _29444_/X _30150_/S VGND VGND VPWR VPWR _30147_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19957_ _34179_/Q _34115_/Q _34051_/Q _33987_/Q _19746_/X _19747_/X VGND VGND VPWR
+ VPWR _19957_/X sky130_fd_sc_hd__mux4_1
XFILLER_214_1300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_268_CLK clkbuf_6_60__f_CLK/X VGND VGND VPWR VPWR _34626_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_113_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18908_ _32869_/Q _32805_/Q _32741_/Q _32677_/Q _18587_/X _18588_/X VGND VGND VPWR
+ VPWR _18908_/X sky130_fd_sc_hd__mux4_1
X_34954_ _34954_/CLK _34954_/D VGND VGND VPWR VPWR _34954_/Q sky130_fd_sc_hd__dfxtp_1
X_30077_ _35290_/Q _29342_/X _30087_/S VGND VGND VPWR VPWR _30078_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19888_ _19888_/A _19888_/B _19888_/C _19888_/D VGND VGND VPWR VPWR _19889_/A sky130_fd_sc_hd__or4_4
XFILLER_132_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33905_ _36082_/CLK _33905_/D VGND VGND VPWR VPWR _33905_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18839_ _33123_/Q _36003_/Q _32995_/Q _32931_/Q _18656_/X _18657_/X VGND VGND VPWR
+ VPWR _18839_/X sky130_fd_sc_hd__mux4_1
XFILLER_110_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34885_ _34949_/CLK _34885_/D VGND VGND VPWR VPWR _34885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33836_ _36076_/CLK _33836_/D VGND VGND VPWR VPWR _33836_/Q sky130_fd_sc_hd__dfxtp_1
X_21850_ _21846_/X _21849_/X _21740_/X _21741_/X VGND VGND VPWR VPWR _21867_/B sky130_fd_sc_hd__o211a_1
XFILLER_167_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20801_ _34649_/Q _34585_/Q _34521_/Q _34457_/Q _20679_/X _20680_/X VGND VGND VPWR
+ VPWR _20801_/X sky130_fd_sc_hd__mux4_1
X_33767_ _36072_/CLK _33767_/D VGND VGND VPWR VPWR _33767_/Q sky130_fd_sc_hd__dfxtp_1
X_21781_ _21667_/X _21779_/X _21780_/X _21671_/X VGND VGND VPWR VPWR _21781_/X sky130_fd_sc_hd__a22o_1
XFILLER_247_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30979_ _35718_/Q input43/X _30981_/S VGND VGND VPWR VPWR _30980_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23520_ _32255_/Q _23426_/X _23536_/S VGND VGND VPWR VPWR _23521_/A sky130_fd_sc_hd__mux2_1
X_35506_ _35698_/CLK _35506_/D VGND VGND VPWR VPWR _35506_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_440_CLK clkbuf_6_37__f_CLK/X VGND VGND VPWR VPWR _35955_/CLK sky130_fd_sc_hd__clkbuf_16
X_20732_ _35159_/Q _35095_/Q _35031_/Q _32151_/Q _20683_/X _20685_/X VGND VGND VPWR
+ VPWR _20732_/X sky130_fd_sc_hd__mux4_1
XFILLER_208_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32718_ _32911_/CLK _32718_/D VGND VGND VPWR VPWR _32718_/Q sky130_fd_sc_hd__dfxtp_1
X_33698_ _35618_/CLK _33698_/D VGND VGND VPWR VPWR _33698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23451_ _32229_/Q _23450_/X _23451_/S VGND VGND VPWR VPWR _23452_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35437_ _35694_/CLK _35437_/D VGND VGND VPWR VPWR _35437_/Q sky130_fd_sc_hd__dfxtp_1
X_20663_ _20663_/A VGND VGND VPWR VPWR _22451_/A sky130_fd_sc_hd__buf_12
X_32649_ _36040_/CLK _32649_/D VGND VGND VPWR VPWR _32649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22402_ _22152_/X _22398_/X _22401_/X _22157_/X VGND VGND VPWR VPWR _22402_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26170_ _24927_/X _33535_/Q _26186_/S VGND VGND VPWR VPWR _26171_/A sky130_fd_sc_hd__mux2_1
X_23382_ _32206_/Q _23381_/X _23385_/S VGND VGND VPWR VPWR _23383_/A sky130_fd_sc_hd__mux2_1
X_35368_ _35685_/CLK _35368_/D VGND VGND VPWR VPWR _35368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20594_ _20663_/A VGND VGND VPWR VPWR _22400_/A sky130_fd_sc_hd__buf_12
XFILLER_149_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25121_ _25121_/A VGND VGND VPWR VPWR _33040_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34319_ _36175_/CLK _34319_/D VGND VGND VPWR VPWR _34319_/Q sky130_fd_sc_hd__dfxtp_1
X_22333_ _22159_/X _22329_/X _22332_/X _22162_/X VGND VGND VPWR VPWR _22333_/X sky130_fd_sc_hd__a22o_1
XFILLER_104_1168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35299_ _35814_/CLK _35299_/D VGND VGND VPWR VPWR _35299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25052_ _25052_/A VGND VGND VPWR VPWR _33007_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22264_ _33155_/Q _36035_/Q _33027_/Q _32963_/Q _22015_/X _22016_/X VGND VGND VPWR
+ VPWR _22264_/X sky130_fd_sc_hd__mux4_1
XFILLER_219_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24003_ _22918_/X _32544_/Q _24021_/S VGND VGND VPWR VPWR _24004_/A sky130_fd_sc_hd__mux2_1
X_21215_ _20892_/X _21213_/X _21214_/X _20895_/X VGND VGND VPWR VPWR _21215_/X sky130_fd_sc_hd__a22o_1
X_29860_ _29860_/A VGND VGND VPWR VPWR _35187_/D sky130_fd_sc_hd__clkbuf_1
X_22195_ _22159_/X _22193_/X _22194_/X _22162_/X VGND VGND VPWR VPWR _22195_/X sky130_fd_sc_hd__a22o_1
XFILLER_183_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28811_ _34720_/Q _27065_/X _28829_/S VGND VGND VPWR VPWR _28812_/A sky130_fd_sc_hd__mux2_1
X_21146_ _35619_/Q _34979_/Q _34339_/Q _33699_/Q _21038_/X _21039_/X VGND VGND VPWR
+ VPWR _21146_/X sky130_fd_sc_hd__mux4_1
X_29791_ _35155_/Q _29518_/X _29795_/S VGND VGND VPWR VPWR _29792_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_259_CLK clkbuf_6_62__f_CLK/X VGND VGND VPWR VPWR _36159_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_28_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28742_ _28742_/A VGND VGND VPWR VPWR _34688_/D sky130_fd_sc_hd__clkbuf_1
X_25954_ _25954_/A VGND VGND VPWR VPWR _33432_/D sky130_fd_sc_hd__clkbuf_1
X_21077_ _35681_/Q _32188_/Q _35553_/Q _35489_/Q _20858_/X _20859_/X VGND VGND VPWR
+ VPWR _21077_/X sky130_fd_sc_hd__mux4_1
XFILLER_115_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_1125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20028_ _19852_/X _20026_/X _20027_/X _19857_/X VGND VGND VPWR VPWR _20028_/X sky130_fd_sc_hd__a22o_1
XFILLER_232_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24905_ input28/X VGND VGND VPWR VPWR _24905_/X sky130_fd_sc_hd__clkbuf_4
X_25885_ _24905_/X _33400_/Q _25895_/S VGND VGND VPWR VPWR _25886_/A sky130_fd_sc_hd__mux2_1
X_28673_ _28784_/S VGND VGND VPWR VPWR _28692_/S sky130_fd_sc_hd__buf_4
XFILLER_246_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_246_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27624_ _27624_/A VGND VGND VPWR VPWR _34190_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_246_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24836_ _24836_/A VGND VGND VPWR VPWR _32929_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24767_ _24794_/S VGND VGND VPWR VPWR _24786_/S sky130_fd_sc_hd__buf_4
XFILLER_27_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27555_ _27555_/A VGND VGND VPWR VPWR _34157_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21979_ _33915_/Q _33851_/Q _33787_/Q _36091_/Q _21977_/X _21978_/X VGND VGND VPWR
+ VPWR _21979_/X sky130_fd_sc_hd__mux4_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_431_CLK clkbuf_6_38__f_CLK/X VGND VGND VPWR VPWR _36020_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_215_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23718_ _23718_/A VGND VGND VPWR VPWR _32346_/D sky130_fd_sc_hd__clkbuf_1
X_26506_ _26506_/A VGND VGND VPWR VPWR _33693_/D sky130_fd_sc_hd__clkbuf_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27486_ _34125_/Q _27205_/X _27494_/S VGND VGND VPWR VPWR _27487_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24698_ _22940_/X _32871_/Q _24702_/S VGND VGND VPWR VPWR _24699_/A sky130_fd_sc_hd__mux2_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29225_ _29225_/A VGND VGND VPWR VPWR _34916_/D sky130_fd_sc_hd__clkbuf_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26437_ _26437_/A VGND VGND VPWR VPWR _33661_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23649_ _23649_/A VGND VGND VPWR VPWR _32315_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17170_ _34165_/Q _34101_/Q _34037_/Q _33973_/Q _17093_/X _17094_/X VGND VGND VPWR
+ VPWR _17170_/X sky130_fd_sc_hd__mux4_1
X_29156_ _34884_/Q _27177_/X _29162_/S VGND VGND VPWR VPWR _29157_/A sky130_fd_sc_hd__mux2_1
X_26368_ _26368_/A VGND VGND VPWR VPWR _33628_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16121_ _32855_/Q _32791_/Q _32727_/Q _32663_/Q _16037_/X _16039_/X VGND VGND VPWR
+ VPWR _16121_/X sky130_fd_sc_hd__mux4_1
XFILLER_35_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28107_ _28107_/A VGND VGND VPWR VPWR _34388_/D sky130_fd_sc_hd__clkbuf_1
X_25319_ _25319_/A VGND VGND VPWR VPWR _33132_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26299_ _26299_/A VGND VGND VPWR VPWR _33596_/D sky130_fd_sc_hd__clkbuf_1
X_29087_ _34851_/Q _27075_/X _29099_/S VGND VGND VPWR VPWR _29088_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16052_ _17982_/A VGND VGND VPWR VPWR _17998_/A sky130_fd_sc_hd__buf_12
X_28038_ _28038_/A VGND VGND VPWR VPWR _34355_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_237_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_498_CLK clkbuf_6_2__f_CLK/X VGND VGND VPWR VPWR _35624_/CLK sky130_fd_sc_hd__clkbuf_16
Xclkbuf_0_CLK CLK VGND VGND VPWR VPWR clkbuf_0_CLK/X sky130_fd_sc_hd__clkbuf_16
X_30000_ _30000_/A VGND VGND VPWR VPWR _35253_/D sky130_fd_sc_hd__clkbuf_1
X_19811_ _20164_/A VGND VGND VPWR VPWR _19811_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_237_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29989_ _29989_/A VGND VGND VPWR VPWR _35248_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19742_ _19738_/X _19741_/X _19465_/X VGND VGND VPWR VPWR _19743_/D sky130_fd_sc_hd__o21ba_1
X_16954_ _33903_/Q _33839_/Q _33775_/Q _36079_/Q _16671_/X _16672_/X VGND VGND VPWR
+ VPWR _16954_/X sky130_fd_sc_hd__mux4_1
X_31951_ _31951_/A VGND VGND VPWR VPWR _36178_/D sky130_fd_sc_hd__clkbuf_1
X_19673_ _33659_/Q _33595_/Q _33531_/Q _33467_/Q _19500_/X _19501_/X VGND VGND VPWR
+ VPWR _19673_/X sky130_fd_sc_hd__mux4_1
X_16885_ _34157_/Q _34093_/Q _34029_/Q _33965_/Q _16740_/X _16741_/X VGND VGND VPWR
+ VPWR _16885_/X sky130_fd_sc_hd__mux4_1
X_18624_ _33117_/Q _35997_/Q _32989_/Q _32925_/Q _18324_/X _18325_/X VGND VGND VPWR
+ VPWR _18624_/X sky130_fd_sc_hd__mux4_1
XFILLER_49_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30902_ _35681_/Q input3/X _30918_/S VGND VGND VPWR VPWR _30903_/A sky130_fd_sc_hd__mux2_1
XTAP_4170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34670_ _34926_/CLK _34670_/D VGND VGND VPWR VPWR _34670_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31882_ _31882_/A VGND VGND VPWR VPWR _36145_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33621_ _33685_/CLK _33621_/D VGND VGND VPWR VPWR _33621_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18555_ _32859_/Q _32795_/Q _32731_/Q _32667_/Q _18337_/X _18339_/X VGND VGND VPWR
+ VPWR _18555_/X sky130_fd_sc_hd__mux4_1
X_30833_ _30833_/A VGND VGND VPWR VPWR _35648_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_422_CLK clkbuf_6_33__f_CLK/X VGND VGND VPWR VPWR _35377_/CLK sky130_fd_sc_hd__clkbuf_16
X_17506_ _17859_/A VGND VGND VPWR VPWR _17506_/X sky130_fd_sc_hd__clkbuf_4
X_33552_ _34064_/CLK _33552_/D VGND VGND VPWR VPWR _33552_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18486_ _33113_/Q _35993_/Q _32985_/Q _32921_/Q _18324_/X _18325_/X VGND VGND VPWR
+ VPWR _18486_/X sky130_fd_sc_hd__mux4_1
X_30764_ _30875_/S VGND VGND VPWR VPWR _30783_/S sky130_fd_sc_hd__buf_4
XFILLER_166_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32503_ _36023_/CLK _32503_/D VGND VGND VPWR VPWR _32503_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17437_ _35196_/Q _35132_/Q _35068_/Q _32252_/Q _17363_/X _17364_/X VGND VGND VPWR
+ VPWR _17437_/X sky130_fd_sc_hd__mux4_1
X_33483_ _34188_/CLK _33483_/D VGND VGND VPWR VPWR _33483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30695_ _35583_/Q _29457_/X _30711_/S VGND VGND VPWR VPWR _30696_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_1460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35222_ _36118_/CLK _35222_/D VGND VGND VPWR VPWR _35222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32434_ _33895_/CLK _32434_/D VGND VGND VPWR VPWR _32434_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17368_ _34938_/Q _34874_/Q _34810_/Q _34746_/Q _17160_/X _17161_/X VGND VGND VPWR
+ VPWR _17368_/X sky130_fd_sc_hd__mux4_1
XFILLER_186_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19107_ _20166_/A VGND VGND VPWR VPWR _19107_/X sky130_fd_sc_hd__buf_4
X_35153_ _36115_/CLK _35153_/D VGND VGND VPWR VPWR _35153_/Q sky130_fd_sc_hd__dfxtp_1
X_16319_ _17851_/A VGND VGND VPWR VPWR _16319_/X sky130_fd_sc_hd__buf_4
X_32365_ _35951_/CLK _32365_/D VGND VGND VPWR VPWR _32365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17299_ _17158_/X _17297_/X _17298_/X _17163_/X VGND VGND VPWR VPWR _17299_/X sky130_fd_sc_hd__a22o_1
X_34104_ _35320_/CLK _34104_/D VGND VGND VPWR VPWR _34104_/Q sky130_fd_sc_hd__dfxtp_1
X_19038_ _19038_/A VGND VGND VPWR VPWR _32424_/D sky130_fd_sc_hd__clkbuf_1
X_31316_ _27689_/X _35877_/Q _31324_/S VGND VGND VPWR VPWR _31317_/A sky130_fd_sc_hd__mux2_1
X_35084_ _35147_/CLK _35084_/D VGND VGND VPWR VPWR _35084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput101 _31959_/Q VGND VGND VPWR VPWR D1[1] sky130_fd_sc_hd__buf_2
X_32296_ _32873_/CLK _32296_/D VGND VGND VPWR VPWR _32296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput112 _31960_/Q VGND VGND VPWR VPWR D1[2] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_489_CLK clkbuf_6_9__f_CLK/X VGND VGND VPWR VPWR _35691_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_138_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34035_ _34035_/CLK _34035_/D VGND VGND VPWR VPWR _34035_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput123 _31961_/Q VGND VGND VPWR VPWR D1[3] sky130_fd_sc_hd__buf_2
X_31247_ _31247_/A VGND VGND VPWR VPWR _35844_/D sky130_fd_sc_hd__clkbuf_1
Xoutput134 _31962_/Q VGND VGND VPWR VPWR D1[4] sky130_fd_sc_hd__buf_2
Xoutput145 _31963_/Q VGND VGND VPWR VPWR D1[5] sky130_fd_sc_hd__buf_2
Xoutput156 _36193_/Q VGND VGND VPWR VPWR D2[11] sky130_fd_sc_hd__buf_2
XFILLER_114_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21000_ _20961_/X _20998_/X _20999_/X _20965_/X VGND VGND VPWR VPWR _21000_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_902 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput167 _36203_/Q VGND VGND VPWR VPWR D2[21] sky130_fd_sc_hd__buf_2
XFILLER_82_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput178 _36213_/Q VGND VGND VPWR VPWR D2[31] sky130_fd_sc_hd__buf_2
Xoutput189 _36223_/Q VGND VGND VPWR VPWR D2[41] sky130_fd_sc_hd__buf_2
XFILLER_153_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31178_ _31178_/A VGND VGND VPWR VPWR _35811_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30129_ _35315_/Q _29419_/X _30129_/S VGND VGND VPWR VPWR _30130_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_1303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35986_ _35986_/CLK _35986_/D VGND VGND VPWR VPWR _35986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34937_ _36153_/CLK _34937_/D VGND VGND VPWR VPWR _34937_/Q sky130_fd_sc_hd__dfxtp_1
X_22951_ _22949_/X _32042_/Q _22978_/S VGND VGND VPWR VPWR _22952_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21902_ _21902_/A VGND VGND VPWR VPWR _36216_/D sky130_fd_sc_hd__buf_6
XFILLER_243_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25670_ _25670_/A VGND VGND VPWR VPWR _33298_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_216_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22882_ input84/X VGND VGND VPWR VPWR _25132_/A sky130_fd_sc_hd__buf_2
XFILLER_3_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34868_ _35828_/CLK _34868_/D VGND VGND VPWR VPWR _34868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24621_ _24621_/A VGND VGND VPWR VPWR _32834_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33819_ _36059_/CLK _33819_/D VGND VGND VPWR VPWR _33819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21833_ _21758_/X _21831_/X _21832_/X _21763_/X VGND VGND VPWR VPWR _21833_/X sky130_fd_sc_hd__a22o_1
XFILLER_71_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34799_ _34926_/CLK _34799_/D VGND VGND VPWR VPWR _34799_/Q sky130_fd_sc_hd__dfxtp_1
X_27340_ _27367_/S VGND VGND VPWR VPWR _27359_/S sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_413_CLK clkbuf_6_32__f_CLK/X VGND VGND VPWR VPWR _36080_/CLK sky130_fd_sc_hd__clkbuf_16
X_24552_ _24552_/A VGND VGND VPWR VPWR _32801_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21764_ _21758_/X _21759_/X _21762_/X _21763_/X VGND VGND VPWR VPWR _21764_/X sky130_fd_sc_hd__a22o_1
XFILLER_19_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_816 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23503_ _32247_/Q _23399_/X _23515_/S VGND VGND VPWR VPWR _23504_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_6_54__f_CLK clkbuf_5_27_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_54__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_20715_ _20601_/X _20711_/X _20714_/X _20607_/X VGND VGND VPWR VPWR _20715_/X sky130_fd_sc_hd__a22o_1
X_27271_ _34023_/Q _27087_/X _27275_/S VGND VGND VPWR VPWR _27272_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24483_ _23021_/X _32769_/Q _24495_/S VGND VGND VPWR VPWR _24484_/A sky130_fd_sc_hd__mux2_1
X_21695_ _34163_/Q _34099_/Q _34035_/Q _33971_/Q _21693_/X _21694_/X VGND VGND VPWR
+ VPWR _21695_/X sky130_fd_sc_hd__mux4_1
XFILLER_239_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29010_ _29010_/A VGND VGND VPWR VPWR _34814_/D sky130_fd_sc_hd__clkbuf_1
X_26222_ _26222_/A VGND VGND VPWR VPWR _33559_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23434_ _23434_/A VGND VGND VPWR VPWR _32223_/D sky130_fd_sc_hd__clkbuf_1
X_20646_ _22447_/A VGND VGND VPWR VPWR _20646_/X sky130_fd_sc_hd__buf_4
XFILLER_165_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26153_ _24902_/X _33527_/Q _26165_/S VGND VGND VPWR VPWR _26154_/A sky130_fd_sc_hd__mux2_1
X_23365_ _32198_/Q _23364_/X _23424_/S VGND VGND VPWR VPWR _23366_/A sky130_fd_sc_hd__mux2_1
X_20577_ _20577_/A _20577_/B _20577_/C _20577_/D VGND VGND VPWR VPWR _20578_/A sky130_fd_sc_hd__or4_1
X_25104_ _24954_/X _33032_/Q _25122_/S VGND VGND VPWR VPWR _25105_/A sky130_fd_sc_hd__mux2_1
X_22316_ _22316_/A VGND VGND VPWR VPWR _22316_/X sky130_fd_sc_hd__buf_6
XFILLER_180_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26084_ _24796_/X _33494_/Q _26102_/S VGND VGND VPWR VPWR _26085_/A sky130_fd_sc_hd__mux2_1
X_23296_ input14/X VGND VGND VPWR VPWR _23296_/X sky130_fd_sc_hd__buf_4
XFILLER_127_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29912_ _35212_/Q _29497_/X _29922_/S VGND VGND VPWR VPWR _29913_/A sky130_fd_sc_hd__mux2_1
X_25035_ _25035_/A VGND VGND VPWR VPWR _32999_/D sky130_fd_sc_hd__clkbuf_1
X_22247_ _34690_/Q _34626_/Q _34562_/Q _34498_/Q _22245_/X _22246_/X VGND VGND VPWR
+ VPWR _22247_/X sky130_fd_sc_hd__mux4_1
XFILLER_219_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29843_ _35179_/Q _29395_/X _29859_/S VGND VGND VPWR VPWR _29844_/A sky130_fd_sc_hd__mux2_1
X_22178_ _22174_/X _22177_/X _22104_/X VGND VGND VPWR VPWR _22188_/C sky130_fd_sc_hd__o21ba_1
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21129_ _21129_/A _21129_/B _21129_/C _21129_/D VGND VGND VPWR VPWR _21130_/A sky130_fd_sc_hd__or4_1
X_29774_ _29774_/A VGND VGND VPWR VPWR _35146_/D sky130_fd_sc_hd__clkbuf_1
X_26986_ _33919_/Q _23426_/X _27002_/S VGND VGND VPWR VPWR _26987_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28725_ _28725_/A VGND VGND VPWR VPWR _34680_/D sky130_fd_sc_hd__clkbuf_1
X_25937_ _24982_/X _33425_/Q _25937_/S VGND VGND VPWR VPWR _25938_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_219_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28656_ _28656_/A VGND VGND VPWR VPWR _34647_/D sky130_fd_sc_hd__clkbuf_1
X_16670_ _33383_/Q _33319_/Q _33255_/Q _33191_/Q _16421_/X _16422_/X VGND VGND VPWR
+ VPWR _16670_/X sky130_fd_sc_hd__mux4_1
X_25868_ _24880_/X _33392_/Q _25874_/S VGND VGND VPWR VPWR _25869_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27607_ _27607_/A VGND VGND VPWR VPWR _34182_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24819_ _24818_/X _32924_/Q _24828_/S VGND VGND VPWR VPWR _24820_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28587_ _28587_/A VGND VGND VPWR VPWR _34615_/D sky130_fd_sc_hd__clkbuf_1
X_25799_ _25799_/A VGND VGND VPWR VPWR _33359_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_222_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_404_CLK clkbuf_6_34__f_CLK/X VGND VGND VPWR VPWR _34101_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18340_ _32854_/Q _32790_/Q _32726_/Q _32662_/Q _18337_/X _18339_/X VGND VGND VPWR
+ VPWR _18340_/X sky130_fd_sc_hd__mux4_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27538_ _27538_/A VGND VGND VPWR VPWR _34149_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18271_ _35221_/Q _35157_/Q _35093_/Q _32277_/Q _16092_/X _16094_/X VGND VGND VPWR
+ VPWR _18271_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27469_ _34117_/Q _27180_/X _27473_/S VGND VGND VPWR VPWR _27470_/A sky130_fd_sc_hd__mux2_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29208_ _29208_/A VGND VGND VPWR VPWR _34908_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17222_ _35446_/Q _35382_/Q _35318_/Q _35254_/Q _16901_/X _16902_/X VGND VGND VPWR
+ VPWR _17222_/X sky130_fd_sc_hd__mux4_1
X_30480_ _35481_/Q _29339_/X _30492_/S VGND VGND VPWR VPWR _30481_/A sky130_fd_sc_hd__mux2_1
Xinput14 DW[21] VGND VGND VPWR VPWR input14/X sky130_fd_sc_hd__clkbuf_8
Xinput25 DW[31] VGND VGND VPWR VPWR input25/X sky130_fd_sc_hd__clkbuf_4
X_29139_ _34876_/Q _27152_/X _29141_/S VGND VGND VPWR VPWR _29140_/A sky130_fd_sc_hd__mux2_1
X_17153_ _17153_/A VGND VGND VPWR VPWR _17153_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_196_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput36 DW[41] VGND VGND VPWR VPWR input36/X sky130_fd_sc_hd__buf_6
XFILLER_200_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput47 DW[51] VGND VGND VPWR VPWR input47/X sky130_fd_sc_hd__buf_8
X_16104_ _17871_/A VGND VGND VPWR VPWR _16104_/X sky130_fd_sc_hd__clkbuf_4
Xinput58 DW[61] VGND VGND VPWR VPWR input58/X sky130_fd_sc_hd__buf_8
Xinput69 R1[4] VGND VGND VPWR VPWR input69/X sky130_fd_sc_hd__clkbuf_4
X_32150_ _34585_/CLK _32150_/D VGND VGND VPWR VPWR _32150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17084_ _35186_/Q _35122_/Q _35058_/Q _32209_/Q _17010_/X _17011_/X VGND VGND VPWR
+ VPWR _17084_/X sky130_fd_sc_hd__mux4_1
XFILLER_128_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31101_ _31101_/A VGND VGND VPWR VPWR _35775_/D sky130_fd_sc_hd__clkbuf_1
X_16035_ _32086_/Q _32278_/Q _32342_/Q _35862_/Q _16032_/X _17867_/A VGND VGND VPWR
+ VPWR _16035_/X sky130_fd_sc_hd__mux4_1
XFILLER_237_1130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32081_ _35857_/CLK _32081_/D VGND VGND VPWR VPWR _32081_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31032_ _35743_/Q input64/X _31032_/S VGND VGND VPWR VPWR _31033_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35840_ _36030_/CLK _35840_/D VGND VGND VPWR VPWR _35840_/Q sky130_fd_sc_hd__dfxtp_1
X_17986_ _17986_/A VGND VGND VPWR VPWR _17986_/X sky130_fd_sc_hd__buf_6
X_19725_ _19720_/X _19722_/X _19723_/X _19724_/X VGND VGND VPWR VPWR _19725_/X sky130_fd_sc_hd__a22o_1
X_16937_ _16650_/X _16935_/X _16936_/X _16653_/X VGND VGND VPWR VPWR _16937_/X sky130_fd_sc_hd__a22o_1
X_35771_ _35835_/CLK _35771_/D VGND VGND VPWR VPWR _35771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32983_ _34135_/CLK _32983_/D VGND VGND VPWR VPWR _32983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34722_ _34914_/CLK _34722_/D VGND VGND VPWR VPWR _34722_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31934_ _23463_/X _36170_/Q _31948_/S VGND VGND VPWR VPWR _31935_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19656_ _20164_/A VGND VGND VPWR VPWR _19656_/X sky130_fd_sc_hd__clkbuf_8
X_16868_ _16645_/X _16866_/X _16867_/X _16648_/X VGND VGND VPWR VPWR _16868_/X sky130_fd_sc_hd__a22o_1
XFILLER_77_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18607_ _18378_/X _18603_/X _18606_/X _18388_/X VGND VGND VPWR VPWR _18607_/X sky130_fd_sc_hd__a22o_1
X_34653_ _36229_/CLK _34653_/D VGND VGND VPWR VPWR _34653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19587_ _19298_/X _19585_/X _19586_/X _19301_/X VGND VGND VPWR VPWR _19587_/X sky130_fd_sc_hd__a22o_1
X_31865_ _31865_/A VGND VGND VPWR VPWR _36137_/D sky130_fd_sc_hd__clkbuf_1
X_16799_ _16794_/X _16797_/X _16798_/X VGND VGND VPWR VPWR _16814_/C sky130_fd_sc_hd__o21ba_1
XFILLER_240_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33604_ _34182_/CLK _33604_/D VGND VGND VPWR VPWR _33604_/Q sky130_fd_sc_hd__dfxtp_1
X_18538_ _34394_/Q _36122_/Q _34266_/Q _34202_/Q _18470_/X _18471_/X VGND VGND VPWR
+ VPWR _18538_/X sky130_fd_sc_hd__mux4_1
XFILLER_206_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30816_ _30816_/A VGND VGND VPWR VPWR _35640_/D sky130_fd_sc_hd__clkbuf_1
X_34584_ _34903_/CLK _34584_/D VGND VGND VPWR VPWR _34584_/Q sky130_fd_sc_hd__dfxtp_1
X_31796_ _31796_/A VGND VGND VPWR VPWR _36104_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_1427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33535_ _35453_/CLK _33535_/D VGND VGND VPWR VPWR _33535_/Q sky130_fd_sc_hd__dfxtp_1
X_18469_ _18378_/X _18467_/X _18468_/X _18388_/X VGND VGND VPWR VPWR _18469_/X sky130_fd_sc_hd__a22o_1
X_30747_ _30747_/A VGND VGND VPWR VPWR _35607_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20500_ _32915_/Q _32851_/Q _32787_/Q _32723_/Q _18284_/X _18287_/X VGND VGND VPWR
+ VPWR _20500_/X sky130_fd_sc_hd__mux4_1
XFILLER_32_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33466_ _33913_/CLK _33466_/D VGND VGND VPWR VPWR _33466_/Q sky130_fd_sc_hd__dfxtp_1
X_21480_ _21405_/X _21478_/X _21479_/X _21410_/X VGND VGND VPWR VPWR _21480_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30678_ _35575_/Q _29432_/X _30690_/S VGND VGND VPWR VPWR _30679_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35205_ _35718_/CLK _35205_/D VGND VGND VPWR VPWR _35205_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_523 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20431_ _20205_/X _20429_/X _20430_/X _20210_/X VGND VGND VPWR VPWR _20431_/X sky130_fd_sc_hd__a22o_1
X_32417_ _33573_/CLK _32417_/D VGND VGND VPWR VPWR _32417_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36185_ _36191_/CLK _36185_/D VGND VGND VPWR VPWR _36185_/Q sky130_fd_sc_hd__dfxtp_1
X_33397_ _34100_/CLK _33397_/D VGND VGND VPWR VPWR _33397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35136_ _35715_/CLK _35136_/D VGND VGND VPWR VPWR _35136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23150_ _22974_/X _32114_/Q _23152_/S VGND VGND VPWR VPWR _23151_/A sky130_fd_sc_hd__mux2_1
X_20362_ _20159_/X _20360_/X _20361_/X _20162_/X VGND VGND VPWR VPWR _20362_/X sky130_fd_sc_hd__a22o_1
X_32348_ _35861_/CLK _32348_/D VGND VGND VPWR VPWR _32348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22101_ _35454_/Q _35390_/Q _35326_/Q _35262_/Q _21854_/X _21855_/X VGND VGND VPWR
+ VPWR _22101_/X sky130_fd_sc_hd__mux4_1
XFILLER_31_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23081_ _23081_/A VGND VGND VPWR VPWR _32084_/D sky130_fd_sc_hd__clkbuf_1
X_35067_ _35197_/CLK _35067_/D VGND VGND VPWR VPWR _35067_/Q sky130_fd_sc_hd__dfxtp_1
X_32279_ _35221_/CLK _32279_/D VGND VGND VPWR VPWR _32279_/Q sky130_fd_sc_hd__dfxtp_1
X_20293_ _20004_/X _20291_/X _20292_/X _20007_/X VGND VGND VPWR VPWR _20293_/X sky130_fd_sc_hd__a22o_1
XTAP_6308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22032_ _22536_/A VGND VGND VPWR VPWR _22032_/X sky130_fd_sc_hd__buf_4
X_34018_ _34085_/CLK _34018_/D VGND VGND VPWR VPWR _34018_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26840_ _33850_/Q _23408_/X _26846_/S VGND VGND VPWR VPWR _26841_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23983_ _23983_/A VGND VGND VPWR VPWR _32534_/D sky130_fd_sc_hd__clkbuf_1
X_26771_ _33817_/Q _23240_/X _26783_/S VGND VGND VPWR VPWR _26772_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_217_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35969_ _35969_/CLK _35969_/D VGND VGND VPWR VPWR _35969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28510_ _28510_/A VGND VGND VPWR VPWR _34579_/D sky130_fd_sc_hd__clkbuf_1
X_25722_ _25722_/A VGND VGND VPWR VPWR _33322_/D sky130_fd_sc_hd__clkbuf_1
X_22934_ input7/X VGND VGND VPWR VPWR _22934_/X sky130_fd_sc_hd__buf_4
X_29490_ _29490_/A VGND VGND VPWR VPWR _35017_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28441_ _28441_/A VGND VGND VPWR VPWR _34546_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25653_ _24961_/X _33290_/Q _25667_/S VGND VGND VPWR VPWR _25654_/A sky130_fd_sc_hd__mux2_1
X_22865_ _20581_/X _22863_/X _22864_/X _20591_/X VGND VGND VPWR VPWR _22865_/X sky130_fd_sc_hd__a22o_1
XFILLER_204_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24604_ _24604_/A VGND VGND VPWR VPWR _32826_/D sky130_fd_sc_hd__clkbuf_1
X_21816_ _32886_/Q _32822_/Q _32758_/Q _32694_/Q _21593_/X _21594_/X VGND VGND VPWR
+ VPWR _21816_/X sky130_fd_sc_hd__mux4_1
XFILLER_225_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28372_ _27828_/X _34514_/Q _28378_/S VGND VGND VPWR VPWR _28373_/A sky130_fd_sc_hd__mux2_1
X_25584_ _25584_/A VGND VGND VPWR VPWR _33257_/D sky130_fd_sc_hd__clkbuf_1
XPHY_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22796_ _32659_/Q _32595_/Q _32531_/Q _35987_/Q _22582_/X _21477_/A VGND VGND VPWR
+ VPWR _22796_/X sky130_fd_sc_hd__mux4_1
XFILLER_58_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_911 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24535_ _24535_/A VGND VGND VPWR VPWR _32793_/D sky130_fd_sc_hd__clkbuf_1
X_27323_ _27323_/A VGND VGND VPWR VPWR _34047_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_996 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21747_ _21598_/X _21743_/X _21746_/X _21601_/X VGND VGND VPWR VPWR _21747_/X sky130_fd_sc_hd__a22o_1
XPHY_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27254_ _34015_/Q _27062_/X _27254_/S VGND VGND VPWR VPWR _27255_/A sky130_fd_sc_hd__mux2_1
X_24466_ _22996_/X _32761_/Q _24474_/S VGND VGND VPWR VPWR _24467_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21678_ _22535_/A VGND VGND VPWR VPWR _21678_/X sky130_fd_sc_hd__buf_6
XFILLER_200_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26205_ _24979_/X _33552_/Q _26207_/S VGND VGND VPWR VPWR _26206_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23417_ input33/X VGND VGND VPWR VPWR _23417_/X sky130_fd_sc_hd__buf_4
X_27185_ _27185_/A VGND VGND VPWR VPWR _33990_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20629_ _22373_/A VGND VGND VPWR VPWR _22512_/A sky130_fd_sc_hd__buf_12
X_24397_ _22894_/X _32728_/Q _24411_/S VGND VGND VPWR VPWR _24398_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26136_ _24877_/X _33519_/Q _26144_/S VGND VGND VPWR VPWR _26137_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23348_ _23348_/A VGND VGND VPWR VPWR _32190_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26067_ _26067_/A VGND VGND VPWR VPWR _33486_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23279_ _23279_/A VGND VGND VPWR VPWR _32165_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_238_1450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25018_ _25018_/A VGND VGND VPWR VPWR _32991_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17840_ _32648_/Q _32584_/Q _32520_/Q _35976_/Q _17629_/X _17766_/X VGND VGND VPWR
+ VPWR _17840_/X sky130_fd_sc_hd__mux4_1
X_29826_ _35171_/Q _29370_/X _29838_/S VGND VGND VPWR VPWR _29827_/A sky130_fd_sc_hd__mux2_1
XTAP_6853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29757_ _29757_/A VGND VGND VPWR VPWR _35138_/D sky130_fd_sc_hd__clkbuf_1
X_17771_ _17771_/A VGND VGND VPWR VPWR _17771_/X sky130_fd_sc_hd__clkbuf_4
X_26969_ _33911_/Q _23399_/X _26981_/S VGND VGND VPWR VPWR _26970_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19510_ _19506_/X _19507_/X _19508_/X _19509_/X VGND VGND VPWR VPWR _19510_/X sky130_fd_sc_hd__a22o_1
XFILLER_75_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16722_ _35624_/Q _34984_/Q _34344_/Q _33704_/Q _16438_/X _16439_/X VGND VGND VPWR
+ VPWR _16722_/X sky130_fd_sc_hd__mux4_1
XFILLER_47_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28708_ _28708_/A VGND VGND VPWR VPWR _34672_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29688_ _29688_/A VGND VGND VPWR VPWR _35105_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_208_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19441_ _20147_/A VGND VGND VPWR VPWR _19441_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_228_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28639_ _28639_/A VGND VGND VPWR VPWR _34640_/D sky130_fd_sc_hd__clkbuf_1
X_16653_ _17869_/A VGND VGND VPWR VPWR _16653_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_234_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31650_ _31650_/A VGND VGND VPWR VPWR _36035_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19372_ _19367_/X _19369_/X _19370_/X _19371_/X VGND VGND VPWR VPWR _19372_/X sky130_fd_sc_hd__a22o_1
X_16584_ _16297_/X _16582_/X _16583_/X _16300_/X VGND VGND VPWR VPWR _16584_/X sky130_fd_sc_hd__a22o_1
XFILLER_76_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18323_ _32598_/Q _32534_/Q _32470_/Q _35926_/Q _20166_/A _20017_/A VGND VGND VPWR
+ VPWR _18323_/X sky130_fd_sc_hd__mux4_1
X_30601_ _35539_/Q _29518_/X _30605_/S VGND VGND VPWR VPWR _30602_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31581_ _31581_/A VGND VGND VPWR VPWR _36002_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33320_ _36072_/CLK _33320_/D VGND VGND VPWR VPWR _33320_/Q sky130_fd_sc_hd__dfxtp_1
X_18254_ _16030_/X _18252_/X _18253_/X _16041_/X VGND VGND VPWR VPWR _18254_/X sky130_fd_sc_hd__a22o_1
X_30532_ _35506_/Q _29416_/X _30534_/S VGND VGND VPWR VPWR _30533_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17205_ _17199_/X _17202_/X _17203_/X _17204_/X VGND VGND VPWR VPWR _17205_/X sky130_fd_sc_hd__a22o_1
X_33251_ _33573_/CLK _33251_/D VGND VGND VPWR VPWR _33251_/Q sky130_fd_sc_hd__dfxtp_1
X_18185_ _16060_/X _18183_/X _18184_/X _16072_/X VGND VGND VPWR VPWR _18185_/X sky130_fd_sc_hd__a22o_1
X_30463_ _30463_/A VGND VGND VPWR VPWR _35473_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32202_ _35566_/CLK _32202_/D VGND VGND VPWR VPWR _32202_/Q sky130_fd_sc_hd__dfxtp_1
X_17136_ _17059_/X _17134_/X _17135_/X _17065_/X VGND VGND VPWR VPWR _17136_/X sky130_fd_sc_hd__a22o_1
X_33182_ _36191_/CLK _33182_/D VGND VGND VPWR VPWR _33182_/Q sky130_fd_sc_hd__dfxtp_1
X_30394_ _30394_/A VGND VGND VPWR VPWR _35440_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32133_ _32894_/CLK _32133_/D VGND VGND VPWR VPWR _32133_/Q sky130_fd_sc_hd__dfxtp_1
X_17067_ _17912_/A VGND VGND VPWR VPWR _17067_/X sky130_fd_sc_hd__clkbuf_4
X_16018_ _17905_/A VGND VGND VPWR VPWR _16018_/X sky130_fd_sc_hd__buf_4
XFILLER_131_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32064_ _36030_/CLK _32064_/D VGND VGND VPWR VPWR _32064_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31015_ _31015_/A VGND VGND VPWR VPWR _35734_/D sky130_fd_sc_hd__clkbuf_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35823_ _36015_/CLK _35823_/D VGND VGND VPWR VPWR _35823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17969_ _34443_/Q _36171_/Q _34315_/Q _34251_/Q _17935_/X _17936_/X VGND VGND VPWR
+ VPWR _17969_/X sky130_fd_sc_hd__mux4_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19708_ _33404_/Q _33340_/Q _33276_/Q _33212_/Q _19427_/X _19428_/X VGND VGND VPWR
+ VPWR _19708_/X sky130_fd_sc_hd__mux4_1
X_35754_ _35754_/CLK _35754_/D VGND VGND VPWR VPWR _35754_/Q sky130_fd_sc_hd__dfxtp_1
X_20980_ _34398_/Q _36126_/Q _34270_/Q _34206_/Q _20770_/X _20771_/X VGND VGND VPWR
+ VPWR _20980_/X sky130_fd_sc_hd__mux4_1
X_32966_ _36039_/CLK _32966_/D VGND VGND VPWR VPWR _32966_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34705_ _34705_/CLK _34705_/D VGND VGND VPWR VPWR _34705_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_1199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31917_ _23435_/X _36162_/Q _31927_/S VGND VGND VPWR VPWR _31918_/A sky130_fd_sc_hd__mux2_1
X_19639_ _33914_/Q _33850_/Q _33786_/Q _36090_/Q _19324_/X _19325_/X VGND VGND VPWR
+ VPWR _19639_/X sky130_fd_sc_hd__mux4_1
XFILLER_226_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35685_ _35685_/CLK _35685_/D VGND VGND VPWR VPWR _35685_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_2_2_0_CLK clkbuf_0_CLK/X VGND VGND VPWR VPWR clkbuf_2_2_0_CLK/X sky130_fd_sc_hd__clkbuf_8
X_32897_ _35902_/CLK _32897_/D VGND VGND VPWR VPWR _32897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34636_ _36173_/CLK _34636_/D VGND VGND VPWR VPWR _34636_/Q sky130_fd_sc_hd__dfxtp_1
X_22650_ _32910_/Q _32846_/Q _32782_/Q _32718_/Q _20584_/X _20587_/X VGND VGND VPWR
+ VPWR _22650_/X sky130_fd_sc_hd__mux4_1
XFILLER_129_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31848_ _23265_/X _36129_/Q _31864_/S VGND VGND VPWR VPWR _31849_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_1051 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21601_ _22462_/A VGND VGND VPWR VPWR _21601_/X sky130_fd_sc_hd__clkbuf_4
X_22581_ _22577_/X _22580_/X _22438_/X VGND VGND VPWR VPWR _22607_/A sky130_fd_sc_hd__o21ba_1
X_34567_ _35657_/CLK _34567_/D VGND VGND VPWR VPWR _34567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31779_ _31779_/A VGND VGND VPWR VPWR _36096_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24320_ _24389_/S VGND VGND VPWR VPWR _24339_/S sky130_fd_sc_hd__buf_4
XFILLER_55_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33518_ _33902_/CLK _33518_/D VGND VGND VPWR VPWR _33518_/Q sky130_fd_sc_hd__dfxtp_1
X_21532_ _35694_/Q _32202_/Q _35566_/Q _35502_/Q _21211_/X _21212_/X VGND VGND VPWR
+ VPWR _21532_/X sky130_fd_sc_hd__mux4_1
XFILLER_181_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34498_ _34691_/CLK _34498_/D VGND VGND VPWR VPWR _34498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36237_ _36242_/CLK _36237_/D VGND VGND VPWR VPWR _36237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24251_ _32661_/Q _23498_/X _24251_/S VGND VGND VPWR VPWR _24252_/A sky130_fd_sc_hd__mux2_1
X_21463_ _32876_/Q _32812_/Q _32748_/Q _32684_/Q _21240_/X _21241_/X VGND VGND VPWR
+ VPWR _21463_/X sky130_fd_sc_hd__mux4_1
X_33449_ _33895_/CLK _33449_/D VGND VGND VPWR VPWR _33449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23202_ _23202_/A VGND VGND VPWR VPWR _32138_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_239_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20414_ _35664_/Q _35024_/Q _34384_/Q _33744_/Q _20150_/X _20151_/X VGND VGND VPWR
+ VPWR _20414_/X sky130_fd_sc_hd__mux4_1
XFILLER_193_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36168_ _36171_/CLK _36168_/D VGND VGND VPWR VPWR _36168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24182_ _24251_/S VGND VGND VPWR VPWR _24201_/S sky130_fd_sc_hd__buf_4
X_21394_ _21245_/X _21390_/X _21393_/X _21248_/X VGND VGND VPWR VPWR _21394_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35119_ _35183_/CLK _35119_/D VGND VGND VPWR VPWR _35119_/Q sky130_fd_sc_hd__dfxtp_1
X_23133_ _23223_/S VGND VGND VPWR VPWR _23152_/S sky130_fd_sc_hd__buf_4
X_20345_ _20341_/X _20344_/X _20138_/X VGND VGND VPWR VPWR _20367_/A sky130_fd_sc_hd__o21ba_2
XFILLER_107_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36099_ _36099_/CLK _36099_/D VGND VGND VPWR VPWR _36099_/Q sky130_fd_sc_hd__dfxtp_1
X_28990_ _34805_/Q _27131_/X _29006_/S VGND VGND VPWR VPWR _28991_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27941_ _27941_/A VGND VGND VPWR VPWR _34309_/D sky130_fd_sc_hd__clkbuf_1
X_23064_ input53/X VGND VGND VPWR VPWR _23064_/X sky130_fd_sc_hd__buf_2
X_20276_ _34188_/Q _34124_/Q _34060_/Q _33996_/Q _20099_/X _20100_/X VGND VGND VPWR
+ VPWR _20276_/X sky130_fd_sc_hd__mux4_1
XTAP_6116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22015_ _22586_/A VGND VGND VPWR VPWR _22015_/X sky130_fd_sc_hd__buf_6
XTAP_6149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27872_ _27872_/A VGND VGND VPWR VPWR _34276_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29611_ _29611_/A VGND VGND VPWR VPWR _35069_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26823_ _33842_/Q _23381_/X _26825_/S VGND VGND VPWR VPWR _26824_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29542_ _29542_/A VGND VGND VPWR VPWR _35036_/D sky130_fd_sc_hd__clkbuf_1
X_26754_ _26754_/A VGND VGND VPWR VPWR _33809_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23966_ _23966_/A VGND VGND VPWR VPWR _32527_/D sky130_fd_sc_hd__clkbuf_1
X_25705_ _25705_/A VGND VGND VPWR VPWR _33314_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29473_ _35012_/Q _29472_/X _29482_/S VGND VGND VPWR VPWR _29474_/A sky130_fd_sc_hd__mux2_1
X_22917_ _22917_/A VGND VGND VPWR VPWR _32031_/D sky130_fd_sc_hd__clkbuf_1
X_26685_ _26685_/A VGND VGND VPWR VPWR _33776_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23897_ _23897_/A VGND VGND VPWR VPWR _32494_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_1007 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28424_ _27704_/X _34538_/Q _28442_/S VGND VGND VPWR VPWR _28425_/A sky130_fd_sc_hd__mux2_1
X_22848_ _22848_/A VGND VGND VPWR VPWR _36244_/D sky130_fd_sc_hd__clkbuf_1
X_25636_ _24936_/X _33282_/Q _25646_/S VGND VGND VPWR VPWR _25637_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28355_ _28355_/A VGND VGND VPWR VPWR _34505_/D sky130_fd_sc_hd__clkbuf_1
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22779_ _22775_/X _22778_/X _22457_/A VGND VGND VPWR VPWR _22787_/C sky130_fd_sc_hd__o21ba_1
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25567_ _24834_/X _33249_/Q _25583_/S VGND VGND VPWR VPWR _25568_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27306_ _27306_/A VGND VGND VPWR VPWR _34039_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_966 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24518_ _23073_/X _32786_/Q _24524_/S VGND VGND VPWR VPWR _24519_/A sky130_fd_sc_hd__mux2_1
XFILLER_200_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25498_ _25498_/A VGND VGND VPWR VPWR _33216_/D sky130_fd_sc_hd__clkbuf_1
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28286_ _27701_/X _34473_/Q _28286_/S VGND VGND VPWR VPWR _28287_/A sky130_fd_sc_hd__mux2_1
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_1010 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27237_ _27237_/A VGND VGND VPWR VPWR _34006_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24449_ _22971_/X _32753_/Q _24453_/S VGND VGND VPWR VPWR _24450_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27168_ input38/X VGND VGND VPWR VPWR _27168_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_137_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26119_ _24852_/X _33511_/Q _26123_/S VGND VGND VPWR VPWR _26120_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19990_ _19852_/X _19988_/X _19989_/X _19857_/X VGND VGND VPWR VPWR _19990_/X sky130_fd_sc_hd__a22o_1
X_27099_ _27099_/A VGND VGND VPWR VPWR _33962_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18941_ _20134_/A VGND VGND VPWR VPWR _18941_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_152_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18872_ _33124_/Q _36004_/Q _32996_/Q _32932_/Q _18656_/X _18657_/X VGND VGND VPWR
+ VPWR _18872_/X sky130_fd_sc_hd__mux4_1
XTAP_6650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29809_ _35163_/Q _29345_/X _29817_/S VGND VGND VPWR VPWR _29810_/A sky130_fd_sc_hd__mux2_1
X_17823_ _17506_/X _17821_/X _17822_/X _17509_/X VGND VGND VPWR VPWR _17823_/X sky130_fd_sc_hd__a22o_1
XFILLER_132_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32820_ _32904_/CLK _32820_/D VGND VGND VPWR VPWR _32820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_212_1464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17754_ _17511_/X _17752_/X _17753_/X _17516_/X VGND VGND VPWR VPWR _17754_/X sky130_fd_sc_hd__a22o_1
XTAP_5993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16705_ _16701_/X _16704_/X _16426_/X VGND VGND VPWR VPWR _16737_/A sky130_fd_sc_hd__o21ba_1
XFILLER_48_896 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32751_ _32877_/CLK _32751_/D VGND VGND VPWR VPWR _32751_/Q sky130_fd_sc_hd__dfxtp_1
X_17685_ _17681_/X _17684_/X _17518_/X VGND VGND VPWR VPWR _17686_/D sky130_fd_sc_hd__o21ba_1
XFILLER_74_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31702_ _36060_/Q input61/X _31708_/S VGND VGND VPWR VPWR _31703_/A sky130_fd_sc_hd__mux2_1
X_19424_ _33652_/Q _33588_/Q _33524_/Q _33460_/Q _19147_/X _19148_/X VGND VGND VPWR
+ VPWR _19424_/X sky130_fd_sc_hd__mux4_1
XFILLER_222_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35470_ _35599_/CLK _35470_/D VGND VGND VPWR VPWR _35470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16636_ _32614_/Q _32550_/Q _32486_/Q _35942_/Q _16570_/X _16354_/X VGND VGND VPWR
+ VPWR _16636_/X sky130_fd_sc_hd__mux4_1
X_32682_ _32914_/CLK _32682_/D VGND VGND VPWR VPWR _32682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34421_ _34612_/CLK _34421_/D VGND VGND VPWR VPWR _34421_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_245_1251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19355_ _33394_/Q _33330_/Q _33266_/Q _33202_/Q _19074_/X _19075_/X VGND VGND VPWR
+ VPWR _19355_/X sky130_fd_sc_hd__mux4_1
X_31633_ _31633_/A VGND VGND VPWR VPWR _36027_/D sky130_fd_sc_hd__clkbuf_1
X_16567_ _33892_/Q _33828_/Q _33764_/Q _36068_/Q _16318_/X _16319_/X VGND VGND VPWR
+ VPWR _16567_/X sky130_fd_sc_hd__mux4_1
XFILLER_91_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18306_ _20077_/A VGND VGND VPWR VPWR _20215_/A sky130_fd_sc_hd__buf_12
XFILLER_176_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34352_ _35439_/CLK _34352_/D VGND VGND VPWR VPWR _34352_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31564_ _31564_/A VGND VGND VPWR VPWR _35994_/D sky130_fd_sc_hd__clkbuf_1
X_19286_ _33904_/Q _33840_/Q _33776_/Q _36080_/Q _18971_/X _18972_/X VGND VGND VPWR
+ VPWR _19286_/X sky130_fd_sc_hd__mux4_1
XFILLER_206_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16498_ _17862_/A VGND VGND VPWR VPWR _16498_/X sky130_fd_sc_hd__buf_4
X_33303_ _36059_/CLK _33303_/D VGND VGND VPWR VPWR _33303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18237_ _33108_/Q _32084_/Q _35860_/Q _35796_/Q _16079_/X _16080_/X VGND VGND VPWR
+ VPWR _18237_/X sky130_fd_sc_hd__mux4_1
X_30515_ _30605_/S VGND VGND VPWR VPWR _30534_/S sky130_fd_sc_hd__buf_6
XFILLER_54_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34283_ _36141_/CLK _34283_/D VGND VGND VPWR VPWR _34283_/Q sky130_fd_sc_hd__dfxtp_1
X_31495_ _27754_/X _35962_/Q _31501_/S VGND VGND VPWR VPWR _31496_/A sky130_fd_sc_hd__mux2_1
XFILLER_191_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36022_ _36023_/CLK _36022_/D VGND VGND VPWR VPWR _36022_/Q sky130_fd_sc_hd__dfxtp_1
X_33234_ _36179_/CLK _33234_/D VGND VGND VPWR VPWR _33234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30446_ _35465_/Q _29488_/X _30462_/S VGND VGND VPWR VPWR _30447_/A sky130_fd_sc_hd__mux2_1
X_18168_ _17153_/A _18166_/X _18167_/X _17156_/A VGND VGND VPWR VPWR _18168_/X sky130_fd_sc_hd__a22o_1
XFILLER_129_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17119_ _34931_/Q _34867_/Q _34803_/Q _34739_/Q _16807_/X _16808_/X VGND VGND VPWR
+ VPWR _17119_/X sky130_fd_sc_hd__mux4_1
X_33165_ _36045_/CLK _33165_/D VGND VGND VPWR VPWR _33165_/Q sky130_fd_sc_hd__dfxtp_1
X_18099_ _33680_/Q _33616_/Q _33552_/Q _33488_/Q _17906_/X _17907_/X VGND VGND VPWR
+ VPWR _18099_/X sky130_fd_sc_hd__mux4_1
X_30377_ _30377_/A VGND VGND VPWR VPWR _35432_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_176_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20130_ _33672_/Q _33608_/Q _33544_/Q _33480_/Q _19853_/X _19854_/X VGND VGND VPWR
+ VPWR _20130_/X sky130_fd_sc_hd__mux4_1
X_32116_ _32882_/CLK _32116_/D VGND VGND VPWR VPWR _32116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33096_ _35849_/CLK _33096_/D VGND VGND VPWR VPWR _33096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20061_ _33414_/Q _33350_/Q _33286_/Q _33222_/Q _19780_/X _19781_/X VGND VGND VPWR
+ VPWR _20061_/X sky130_fd_sc_hd__mux4_1
X_32047_ _36144_/CLK _32047_/D VGND VGND VPWR VPWR _32047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_920 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35806_ _35807_/CLK _35806_/D VGND VGND VPWR VPWR _35806_/Q sky130_fd_sc_hd__dfxtp_1
X_23820_ _23052_/X _32395_/Q _23832_/S VGND VGND VPWR VPWR _23821_/A sky130_fd_sc_hd__mux2_1
XTAP_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33998_ _34192_/CLK _33998_/D VGND VGND VPWR VPWR _33998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23751_ _22949_/X _32362_/Q _23769_/S VGND VGND VPWR VPWR _23752_/A sky130_fd_sc_hd__mux2_1
X_35737_ _35801_/CLK _35737_/D VGND VGND VPWR VPWR _35737_/Q sky130_fd_sc_hd__dfxtp_1
X_20963_ _32094_/Q _32286_/Q _32350_/Q _35870_/Q _20821_/X _20962_/X VGND VGND VPWR
+ VPWR _20963_/X sky130_fd_sc_hd__mux4_1
XFILLER_113_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32949_ _34485_/CLK _32949_/D VGND VGND VPWR VPWR _32949_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22702_ _33424_/Q _33360_/Q _33296_/Q _33232_/Q _22433_/X _22434_/X VGND VGND VPWR
+ VPWR _22702_/X sky130_fd_sc_hd__mux4_2
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26470_ _33677_/Q _23472_/X _26478_/S VGND VGND VPWR VPWR _26471_/A sky130_fd_sc_hd__mux2_1
XFILLER_199_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23682_ _23052_/X _32331_/Q _23694_/S VGND VGND VPWR VPWR _23683_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35668_ _35668_/CLK _35668_/D VGND VGND VPWR VPWR _35668_/Q sky130_fd_sc_hd__dfxtp_1
X_20894_ _35612_/Q _34972_/Q _34332_/Q _33692_/Q _20653_/X _20655_/X VGND VGND VPWR
+ VPWR _20894_/X sky130_fd_sc_hd__mux4_1
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22633_ _34445_/Q _36173_/Q _34317_/Q _34253_/Q _22535_/X _22536_/X VGND VGND VPWR
+ VPWR _22633_/X sky130_fd_sc_hd__mux4_1
XFILLER_213_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25421_ _24818_/X _33180_/Q _25427_/S VGND VGND VPWR VPWR _25422_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34619_ _34685_/CLK _34619_/D VGND VGND VPWR VPWR _34619_/Q sky130_fd_sc_hd__dfxtp_1
X_35599_ _35599_/CLK _35599_/D VGND VGND VPWR VPWR _35599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28140_ _28140_/A VGND VGND VPWR VPWR _34403_/D sky130_fd_sc_hd__clkbuf_1
X_25352_ _25352_/A VGND VGND VPWR VPWR _33148_/D sky130_fd_sc_hd__clkbuf_1
X_22564_ _22309_/X _22562_/X _22563_/X _22312_/X VGND VGND VPWR VPWR _22564_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21515_ _21515_/A VGND VGND VPWR VPWR _36205_/D sky130_fd_sc_hd__clkbuf_1
X_24303_ _24303_/A VGND VGND VPWR VPWR _32683_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_221_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28071_ _34371_/Q _27174_/X _28079_/S VGND VGND VPWR VPWR _28072_/A sky130_fd_sc_hd__mux2_1
X_25283_ _25283_/A VGND VGND VPWR VPWR _33115_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22495_ _22491_/X _22494_/X _22457_/X VGND VGND VPWR VPWR _22503_/C sky130_fd_sc_hd__o21ba_1
XFILLER_10_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27022_ _27022_/A VGND VGND VPWR VPWR _33936_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24234_ _24234_/A VGND VGND VPWR VPWR _32652_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21446_ _22505_/A VGND VGND VPWR VPWR _21446_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_119_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24165_ _24165_/A VGND VGND VPWR VPWR _32619_/D sky130_fd_sc_hd__clkbuf_1
X_21377_ _33898_/Q _33834_/Q _33770_/Q _36074_/Q _21271_/X _21272_/X VGND VGND VPWR
+ VPWR _21377_/X sky130_fd_sc_hd__mux4_1
XFILLER_163_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23116_ _23116_/A VGND VGND VPWR VPWR _32097_/D sky130_fd_sc_hd__clkbuf_1
X_20328_ _20009_/X _20326_/X _20327_/X _20012_/X VGND VGND VPWR VPWR _20328_/X sky130_fd_sc_hd__a22o_1
X_24096_ _24096_/A VGND VGND VPWR VPWR _32588_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28973_ _34797_/Q _27106_/X _28985_/S VGND VGND VPWR VPWR _28974_/A sky130_fd_sc_hd__mux2_1
XFILLER_134_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23047_ _23046_/X _32073_/Q _23071_/S VGND VGND VPWR VPWR _23048_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27924_ _27924_/A VGND VGND VPWR VPWR _34301_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20259_ _20004_/X _20257_/X _20258_/X _20007_/X VGND VGND VPWR VPWR _20259_/X sky130_fd_sc_hd__a22o_1
XFILLER_77_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27855_ _27855_/A VGND VGND VPWR VPWR _34268_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_6_1__f_CLK clkbuf_5_0_0_CLK/X VGND VGND VPWR VPWR clkbuf_leaf_9_CLK/A sky130_fd_sc_hd__clkbuf_16
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26806_ _26896_/S VGND VGND VPWR VPWR _26825_/S sky130_fd_sc_hd__clkbuf_8
XTAP_5289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27786_ _27785_/X _34244_/Q _27795_/S VGND VGND VPWR VPWR _27787_/A sky130_fd_sc_hd__mux2_1
XTAP_4555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24998_ _25130_/S VGND VGND VPWR VPWR _25017_/S sky130_fd_sc_hd__buf_6
XTAP_3821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29525_ _35029_/Q _29524_/X _29525_/S VGND VGND VPWR VPWR _29526_/A sky130_fd_sc_hd__mux2_1
XTAP_4577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26737_ _33801_/Q _23460_/X _26753_/S VGND VGND VPWR VPWR _26738_/A sky130_fd_sc_hd__mux2_1
XTAP_4588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23949_ _23949_/A VGND VGND VPWR VPWR _32519_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29456_ _29456_/A VGND VGND VPWR VPWR _35006_/D sky130_fd_sc_hd__clkbuf_1
X_17470_ _17153_/X _17468_/X _17469_/X _17156_/X VGND VGND VPWR VPWR _17470_/X sky130_fd_sc_hd__a22o_1
XTAP_3898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26668_ _26668_/A VGND VGND VPWR VPWR _33768_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_204_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16421_ _17799_/A VGND VGND VPWR VPWR _16421_/X sky130_fd_sc_hd__buf_4
X_28407_ _27680_/X _34530_/Q _28421_/S VGND VGND VPWR VPWR _28408_/A sky130_fd_sc_hd__mux2_1
X_25619_ _24911_/X _33274_/Q _25625_/S VGND VGND VPWR VPWR _25620_/A sky130_fd_sc_hd__mux2_1
XFILLER_232_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29387_ _29387_/A VGND VGND VPWR VPWR _34984_/D sky130_fd_sc_hd__clkbuf_1
X_26599_ _26599_/A VGND VGND VPWR VPWR _33737_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19140_ _34411_/Q _36139_/Q _34283_/Q _34219_/Q _18823_/X _18824_/X VGND VGND VPWR
+ VPWR _19140_/X sky130_fd_sc_hd__mux4_1
X_28338_ _28338_/A VGND VGND VPWR VPWR _34497_/D sky130_fd_sc_hd__clkbuf_1
X_16352_ _16348_/X _16351_/X _16015_/X VGND VGND VPWR VPWR _16384_/A sky130_fd_sc_hd__o21ba_1
XFILLER_9_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19071_ _33642_/Q _33578_/Q _33514_/Q _33450_/Q _18794_/X _18795_/X VGND VGND VPWR
+ VPWR _19071_/X sky130_fd_sc_hd__mux4_1
XFILLER_40_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16283_ _32604_/Q _32540_/Q _32476_/Q _35932_/Q _16217_/X _17717_/A VGND VGND VPWR
+ VPWR _16283_/X sky130_fd_sc_hd__mux4_1
XFILLER_121_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28269_ _28269_/A VGND VGND VPWR VPWR _34464_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30300_ _35396_/Q _29472_/X _30306_/S VGND VGND VPWR VPWR _30301_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18022_ _18018_/X _18021_/X _17846_/X _17847_/X VGND VGND VPWR VPWR _18037_/B sky130_fd_sc_hd__o211a_1
XFILLER_172_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31280_ _31280_/A VGND VGND VPWR VPWR _35860_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30231_ _35363_/Q _29370_/X _30243_/S VGND VGND VPWR VPWR _30232_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_962 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30162_ _30162_/A VGND VGND VPWR VPWR _35330_/D sky130_fd_sc_hd__clkbuf_1
X_19973_ _35651_/Q _35011_/Q _34371_/Q _33731_/Q _19797_/X _19798_/X VGND VGND VPWR
+ VPWR _19973_/X sky130_fd_sc_hd__mux4_1
XFILLER_49_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18924_ _34917_/Q _34853_/Q _34789_/Q _34725_/Q _18754_/X _18755_/X VGND VGND VPWR
+ VPWR _18924_/X sky130_fd_sc_hd__mux4_1
X_34970_ _35610_/CLK _34970_/D VGND VGND VPWR VPWR _34970_/Q sky130_fd_sc_hd__dfxtp_1
X_30093_ _30093_/A VGND VGND VPWR VPWR _35297_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33921_ _33921_/CLK _33921_/D VGND VGND VPWR VPWR _33921_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18855_ _35171_/Q _35107_/Q _35043_/Q _32163_/Q _18604_/X _18605_/X VGND VGND VPWR
+ VPWR _18855_/X sky130_fd_sc_hd__mux4_1
XTAP_6480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17806_ _17802_/X _17805_/X _17485_/X VGND VGND VPWR VPWR _17828_/A sky130_fd_sc_hd__o21ba_2
X_33852_ _36092_/CLK _33852_/D VGND VGND VPWR VPWR _33852_/Q sky130_fd_sc_hd__dfxtp_1
X_18786_ _18747_/X _18784_/X _18785_/X _18750_/X VGND VGND VPWR VPWR _18786_/X sky130_fd_sc_hd__a22o_1
XFILLER_212_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15998_ input67/X input68/X VGND VGND VPWR VPWR _15999_/A sky130_fd_sc_hd__and2_1
XFILLER_243_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_939 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32803_ _32871_/CLK _32803_/D VGND VGND VPWR VPWR _32803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17737_ _17412_/X _17735_/X _17736_/X _17418_/X VGND VGND VPWR VPWR _17737_/X sky130_fd_sc_hd__a22o_1
X_33783_ _33910_/CLK _33783_/D VGND VGND VPWR VPWR _33783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30995_ _30995_/A VGND VGND VPWR VPWR _35725_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_844 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35522_ _36033_/CLK _35522_/D VGND VGND VPWR VPWR _35522_/Q sky130_fd_sc_hd__dfxtp_1
X_32734_ _35870_/CLK _32734_/D VGND VGND VPWR VPWR _32734_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17668_ _17420_/X _17666_/X _17667_/X _17424_/X VGND VGND VPWR VPWR _17668_/X sky130_fd_sc_hd__a22o_1
XFILLER_247_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19407_ _19403_/X _19406_/X _19087_/X _19088_/X VGND VGND VPWR VPWR _19422_/B sky130_fd_sc_hd__o211a_1
X_16619_ _16615_/X _16618_/X _16445_/X VGND VGND VPWR VPWR _16627_/C sky130_fd_sc_hd__o21ba_1
X_35453_ _35453_/CLK _35453_/D VGND VGND VPWR VPWR _35453_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32665_ _34070_/CLK _32665_/D VGND VGND VPWR VPWR _32665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17599_ _17412_/X _17597_/X _17598_/X _17418_/X VGND VGND VPWR VPWR _17599_/X sky130_fd_sc_hd__a22o_1
XFILLER_195_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34404_ _34405_/CLK _34404_/D VGND VGND VPWR VPWR _34404_/Q sky130_fd_sc_hd__dfxtp_1
X_19338_ _19298_/X _19336_/X _19337_/X _19301_/X VGND VGND VPWR VPWR _19338_/X sky130_fd_sc_hd__a22o_1
X_31616_ _31616_/A VGND VGND VPWR VPWR _36019_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35384_ _35448_/CLK _35384_/D VGND VGND VPWR VPWR _35384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32596_ _35988_/CLK _32596_/D VGND VGND VPWR VPWR _32596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34335_ _35615_/CLK _34335_/D VGND VGND VPWR VPWR _34335_/Q sky130_fd_sc_hd__dfxtp_1
X_31547_ _27831_/X _35987_/Q _31551_/S VGND VGND VPWR VPWR _31548_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19269_ _35439_/Q _35375_/Q _35311_/Q _35247_/Q _19201_/X _19202_/X VGND VGND VPWR
+ VPWR _19269_/X sky130_fd_sc_hd__mux4_1
X_21300_ _34152_/Q _34088_/Q _34024_/Q _33960_/Q _20987_/X _20988_/X VGND VGND VPWR
+ VPWR _21300_/X sky130_fd_sc_hd__mux4_1
XFILLER_108_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34266_ _36235_/CLK _34266_/D VGND VGND VPWR VPWR _34266_/Q sky130_fd_sc_hd__dfxtp_1
X_22280_ _35203_/Q _35139_/Q _35075_/Q _32259_/Q _21963_/X _21964_/X VGND VGND VPWR
+ VPWR _22280_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31478_ _27729_/X _35954_/Q _31480_/S VGND VGND VPWR VPWR _31479_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36005_ _36005_/CLK _36005_/D VGND VGND VPWR VPWR _36005_/Q sky130_fd_sc_hd__dfxtp_1
X_33217_ _33924_/CLK _33217_/D VGND VGND VPWR VPWR _33217_/Q sky130_fd_sc_hd__dfxtp_1
X_21231_ _21093_/X _21229_/X _21230_/X _21098_/X VGND VGND VPWR VPWR _21231_/X sky130_fd_sc_hd__a22o_1
X_30429_ _35457_/Q _29463_/X _30441_/S VGND VGND VPWR VPWR _30430_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34197_ _34773_/CLK _34197_/D VGND VGND VPWR VPWR _34197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_1104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21162_ _21162_/A VGND VGND VPWR VPWR _36195_/D sky130_fd_sc_hd__clkbuf_1
X_33148_ _35965_/CLK _33148_/D VGND VGND VPWR VPWR _33148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20113_ _20109_/X _20112_/X _19793_/X _19794_/X VGND VGND VPWR VPWR _20128_/B sky130_fd_sc_hd__o211a_1
XFILLER_154_1440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25970_ _24830_/X _33440_/Q _25988_/S VGND VGND VPWR VPWR _25971_/A sky130_fd_sc_hd__mux2_1
X_21093_ _22505_/A VGND VGND VPWR VPWR _21093_/X sky130_fd_sc_hd__buf_4
X_33079_ _35768_/CLK _33079_/D VGND VGND VPWR VPWR _33079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20044_ _20004_/X _20042_/X _20043_/X _20007_/X VGND VGND VPWR VPWR _20044_/X sky130_fd_sc_hd__a22o_1
X_24921_ _24920_/X _32957_/Q _24921_/S VGND VGND VPWR VPWR _24922_/A sky130_fd_sc_hd__mux2_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27640_ input88/X input87/X input86/X VGND VGND VPWR VPWR _27641_/A sky130_fd_sc_hd__and3b_1
X_24852_ input9/X VGND VGND VPWR VPWR _24852_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_58_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23803_ _23027_/X _32387_/Q _23811_/S VGND VGND VPWR VPWR _23804_/A sky130_fd_sc_hd__mux2_1
XTAP_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27571_ _34165_/Q _27131_/X _27587_/S VGND VGND VPWR VPWR _27572_/A sky130_fd_sc_hd__mux2_1
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24783_ _24783_/A VGND VGND VPWR VPWR _32911_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21995_ _21991_/X _21994_/X _21751_/X VGND VGND VPWR VPWR _22003_/C sky130_fd_sc_hd__o21ba_1
XFILLER_227_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29310_ _34957_/Q _27205_/X _29318_/S VGND VGND VPWR VPWR _29311_/A sky130_fd_sc_hd__mux2_1
X_26522_ _24846_/X _33701_/Q _26530_/S VGND VGND VPWR VPWR _26523_/A sky130_fd_sc_hd__mux2_1
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20946_ _33630_/Q _33566_/Q _33502_/Q _33438_/Q _20741_/X _20742_/X VGND VGND VPWR
+ VPWR _20946_/X sky130_fd_sc_hd__mux4_1
X_23734_ _22925_/X _32354_/Q _23748_/S VGND VGND VPWR VPWR _23735_/A sky130_fd_sc_hd__mux2_1
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29241_ _34924_/Q _27103_/X _29255_/S VGND VGND VPWR VPWR _29242_/A sky130_fd_sc_hd__mux2_1
X_26453_ _33669_/Q _23444_/X _26457_/S VGND VGND VPWR VPWR _26454_/A sky130_fd_sc_hd__mux2_1
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20877_ _34140_/Q _34076_/Q _34012_/Q _33948_/Q _20609_/X _20611_/X VGND VGND VPWR
+ VPWR _20877_/X sky130_fd_sc_hd__mux4_1
X_23665_ _23027_/X _32323_/Q _23673_/S VGND VGND VPWR VPWR _23666_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25404_ _25404_/A VGND VGND VPWR VPWR _33173_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29172_ _29172_/A VGND VGND VPWR VPWR _34891_/D sky130_fd_sc_hd__clkbuf_1
X_22616_ _32653_/Q _32589_/Q _32525_/Q _35981_/Q _22582_/X _22366_/X VGND VGND VPWR
+ VPWR _22616_/X sky130_fd_sc_hd__mux4_1
X_23596_ _22925_/X _32290_/Q _23610_/S VGND VGND VPWR VPWR _23597_/A sky130_fd_sc_hd__mux2_1
X_26384_ _33636_/Q _23274_/X _26394_/S VGND VGND VPWR VPWR _26385_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28123_ _28123_/A VGND VGND VPWR VPWR _34395_/D sky130_fd_sc_hd__clkbuf_1
X_22547_ _33931_/Q _33867_/Q _33803_/Q _36107_/Q _22330_/X _22331_/X VGND VGND VPWR
+ VPWR _22547_/X sky130_fd_sc_hd__mux4_1
X_25335_ _33140_/Q _23387_/X _25353_/S VGND VGND VPWR VPWR _25336_/A sky130_fd_sc_hd__mux2_1
XFILLER_220_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28054_ _34363_/Q _27149_/X _28058_/S VGND VGND VPWR VPWR _28055_/A sky130_fd_sc_hd__mux2_1
X_22478_ _33417_/Q _33353_/Q _33289_/Q _33225_/Q _22433_/X _22434_/X VGND VGND VPWR
+ VPWR _22478_/X sky130_fd_sc_hd__mux4_1
X_25266_ _25266_/A VGND VGND VPWR VPWR _33108_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27005_ _33928_/Q _23453_/X _27023_/S VGND VGND VPWR VPWR _27006_/A sky130_fd_sc_hd__mux2_1
X_24217_ _24217_/A VGND VGND VPWR VPWR _32644_/D sky130_fd_sc_hd__clkbuf_1
X_21429_ _21425_/X _21428_/X _21387_/X _21388_/X VGND VGND VPWR VPWR _21444_/B sky130_fd_sc_hd__o211a_1
X_25197_ _25197_/A VGND VGND VPWR VPWR _33075_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24148_ _24148_/A VGND VGND VPWR VPWR _32611_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24079_ _24079_/A VGND VGND VPWR VPWR _32580_/D sky130_fd_sc_hd__clkbuf_1
X_28956_ _34789_/Q _27081_/X _28964_/S VGND VGND VPWR VPWR _28957_/A sky130_fd_sc_hd__mux2_1
X_16970_ _33071_/Q _32047_/Q _35823_/Q _35759_/Q _16725_/X _16726_/X VGND VGND VPWR
+ VPWR _16970_/X sky130_fd_sc_hd__mux4_1
XFILLER_2_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27907_ _27739_/X _34293_/Q _27923_/S VGND VGND VPWR VPWR _27908_/A sky130_fd_sc_hd__mux2_1
XFILLER_237_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28887_ _28887_/A VGND VGND VPWR VPWR _34756_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_237_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18640_ _34397_/Q _36125_/Q _34269_/Q _34205_/Q _18470_/X _18471_/X VGND VGND VPWR
+ VPWR _18640_/X sky130_fd_sc_hd__mux4_1
XTAP_5064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27838_ _27837_/X _34261_/Q _27838_/S VGND VGND VPWR VPWR _27839_/A sky130_fd_sc_hd__mux2_1
XTAP_5075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18571_ _34907_/Q _34843_/Q _34779_/Q _34715_/Q _18396_/X _18398_/X VGND VGND VPWR
+ VPWR _18571_/X sky130_fd_sc_hd__mux4_1
XTAP_4374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27769_ _27769_/A VGND VGND VPWR VPWR _34238_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29508_ _29508_/A VGND VGND VPWR VPWR _35023_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17522_ _33663_/Q _33599_/Q _33535_/Q _33471_/Q _17200_/X _17201_/X VGND VGND VPWR
+ VPWR _17522_/X sky130_fd_sc_hd__mux4_1
XTAP_3673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30780_ _30780_/A VGND VGND VPWR VPWR _35623_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_229_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17453_ _17449_/X _17452_/X _17132_/X VGND VGND VPWR VPWR _17475_/A sky130_fd_sc_hd__o21ba_1
X_29439_ _35001_/Q _29438_/X _29451_/S VGND VGND VPWR VPWR _29440_/A sky130_fd_sc_hd__mux2_1
XTAP_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16404_ _16292_/X _16402_/X _16403_/X _16295_/X VGND VGND VPWR VPWR _16404_/X sky130_fd_sc_hd__a22o_1
X_32450_ _36075_/CLK _32450_/D VGND VGND VPWR VPWR _32450_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17384_ _17059_/X _17382_/X _17383_/X _17065_/X VGND VGND VPWR VPWR _17384_/X sky130_fd_sc_hd__a22o_1
X_31401_ _31401_/A VGND VGND VPWR VPWR _35917_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19123_ _32619_/Q _32555_/Q _32491_/Q _35947_/Q _18870_/X _19007_/X VGND VGND VPWR
+ VPWR _19123_/X sky130_fd_sc_hd__mux4_1
X_16335_ _16297_/X _16333_/X _16334_/X _16300_/X VGND VGND VPWR VPWR _16335_/X sky130_fd_sc_hd__a22o_1
X_32381_ _35964_/CLK _32381_/D VGND VGND VPWR VPWR _32381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34120_ _34185_/CLK _34120_/D VGND VGND VPWR VPWR _34120_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31332_ _31332_/A VGND VGND VPWR VPWR _35884_/D sky130_fd_sc_hd__clkbuf_1
X_19054_ _19050_/X _19053_/X _18734_/X _18735_/X VGND VGND VPWR VPWR _19069_/B sky130_fd_sc_hd__o211a_1
X_16266_ _16262_/X _16265_/X _16075_/X VGND VGND VPWR VPWR _16274_/C sky130_fd_sc_hd__o21ba_1
XFILLER_200_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18005_ _17864_/X _18003_/X _18004_/X _17869_/X VGND VGND VPWR VPWR _18005_/X sky130_fd_sc_hd__a22o_1
X_34051_ _34183_/CLK _34051_/D VGND VGND VPWR VPWR _34051_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31263_ _27810_/X _35852_/Q _31273_/S VGND VGND VPWR VPWR _31264_/A sky130_fd_sc_hd__mux2_1
X_16197_ _35417_/Q _35353_/Q _35289_/Q _35225_/Q _16195_/X _16196_/X VGND VGND VPWR
+ VPWR _16197_/X sky130_fd_sc_hd__mux4_1
X_33002_ _36010_/CLK _33002_/D VGND VGND VPWR VPWR _33002_/Q sky130_fd_sc_hd__dfxtp_1
X_30214_ _35355_/Q _29345_/X _30222_/S VGND VGND VPWR VPWR _30215_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31194_ _27708_/X _35819_/Q _31210_/S VGND VGND VPWR VPWR _31195_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30145_ _30145_/A VGND VGND VPWR VPWR _35322_/D sky130_fd_sc_hd__clkbuf_1
X_19956_ _33667_/Q _33603_/Q _33539_/Q _33475_/Q _19853_/X _19854_/X VGND VGND VPWR
+ VPWR _19956_/X sky130_fd_sc_hd__mux4_1
XFILLER_214_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_218_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18907_ _32101_/Q _32293_/Q _32357_/Q _35877_/Q _18874_/X _18662_/X VGND VGND VPWR
+ VPWR _18907_/X sky130_fd_sc_hd__mux4_1
X_34953_ _34954_/CLK _34953_/D VGND VGND VPWR VPWR _34953_/Q sky130_fd_sc_hd__dfxtp_1
X_30076_ _30076_/A VGND VGND VPWR VPWR _35289_/D sky130_fd_sc_hd__clkbuf_1
X_19887_ _19881_/X _19886_/X _19818_/X VGND VGND VPWR VPWR _19888_/D sky130_fd_sc_hd__o21ba_1
XFILLER_68_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33904_ _33904_/CLK _33904_/D VGND VGND VPWR VPWR _33904_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18838_ _32611_/Q _32547_/Q _32483_/Q _35939_/Q _18517_/X _18654_/X VGND VGND VPWR
+ VPWR _18838_/X sky130_fd_sc_hd__mux4_1
X_34884_ _34949_/CLK _34884_/D VGND VGND VPWR VPWR _34884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33835_ _33895_/CLK _33835_/D VGND VGND VPWR VPWR _33835_/Q sky130_fd_sc_hd__dfxtp_1
X_18769_ _18765_/X _18768_/X _18726_/X VGND VGND VPWR VPWR _18791_/A sky130_fd_sc_hd__o21ba_1
XFILLER_243_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_247_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20800_ _20794_/X _20799_/X _20675_/X VGND VGND VPWR VPWR _20808_/C sky130_fd_sc_hd__o21ba_1
X_33766_ _36066_/CLK _33766_/D VGND VGND VPWR VPWR _33766_/Q sky130_fd_sc_hd__dfxtp_1
X_21780_ _32885_/Q _32821_/Q _32757_/Q _32693_/Q _21593_/X _21594_/X VGND VGND VPWR
+ VPWR _21780_/X sky130_fd_sc_hd__mux4_1
X_30978_ _30978_/A VGND VGND VPWR VPWR _35717_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20731_ _34647_/Q _34583_/Q _34519_/Q _34455_/Q _20679_/X _20680_/X VGND VGND VPWR
+ VPWR _20731_/X sky130_fd_sc_hd__mux4_1
X_35505_ _35697_/CLK _35505_/D VGND VGND VPWR VPWR _35505_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_819 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32717_ _32909_/CLK _32717_/D VGND VGND VPWR VPWR _32717_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33697_ _33697_/CLK _33697_/D VGND VGND VPWR VPWR _33697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23450_ input44/X VGND VGND VPWR VPWR _23450_/X sky130_fd_sc_hd__buf_6
X_20662_ _22450_/A VGND VGND VPWR VPWR _20662_/X sky130_fd_sc_hd__buf_6
XFILLER_211_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32648_ _36040_/CLK _32648_/D VGND VGND VPWR VPWR _32648_/Q sky130_fd_sc_hd__dfxtp_1
X_35436_ _35564_/CLK _35436_/D VGND VGND VPWR VPWR _35436_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22401_ _34183_/Q _34119_/Q _34055_/Q _33991_/Q _22399_/X _22400_/X VGND VGND VPWR
+ VPWR _22401_/X sky130_fd_sc_hd__mux4_1
XFILLER_108_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23381_ input21/X VGND VGND VPWR VPWR _23381_/X sky130_fd_sc_hd__buf_4
X_20593_ _22399_/A VGND VGND VPWR VPWR _20593_/X sky130_fd_sc_hd__buf_4
X_32579_ _35907_/CLK _32579_/D VGND VGND VPWR VPWR _32579_/Q sky130_fd_sc_hd__dfxtp_1
X_35367_ _35367_/CLK _35367_/D VGND VGND VPWR VPWR _35367_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22332_ _33925_/Q _33861_/Q _33797_/Q _36101_/Q _22330_/X _22331_/X VGND VGND VPWR
+ VPWR _22332_/X sky130_fd_sc_hd__mux4_1
X_25120_ _24979_/X _33040_/Q _25122_/S VGND VGND VPWR VPWR _25121_/A sky130_fd_sc_hd__mux2_1
X_34318_ _36176_/CLK _34318_/D VGND VGND VPWR VPWR _34318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35298_ _35553_/CLK _35298_/D VGND VGND VPWR VPWR _35298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_1248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25051_ _24877_/X _33007_/Q _25059_/S VGND VGND VPWR VPWR _25052_/A sky130_fd_sc_hd__mux2_1
X_34249_ _36169_/CLK _34249_/D VGND VGND VPWR VPWR _34249_/Q sky130_fd_sc_hd__dfxtp_1
X_22263_ _32643_/Q _32579_/Q _32515_/Q _35971_/Q _22229_/X _22013_/X VGND VGND VPWR
+ VPWR _22263_/X sky130_fd_sc_hd__mux4_1
X_24002_ _24113_/S VGND VGND VPWR VPWR _24021_/S sky130_fd_sc_hd__buf_4
XFILLER_3_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21214_ _35621_/Q _34981_/Q _34341_/Q _33701_/Q _21038_/X _21039_/X VGND VGND VPWR
+ VPWR _21214_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22194_ _33921_/Q _33857_/Q _33793_/Q _36097_/Q _21977_/X _21978_/X VGND VGND VPWR
+ VPWR _22194_/X sky130_fd_sc_hd__mux4_1
XFILLER_219_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28810_ _28921_/S VGND VGND VPWR VPWR _28829_/S sky130_fd_sc_hd__buf_4
X_21145_ _35683_/Q _32190_/Q _35555_/Q _35491_/Q _20858_/X _20859_/X VGND VGND VPWR
+ VPWR _21145_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29790_ _29790_/A VGND VGND VPWR VPWR _35154_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_6_14__f_CLK clkbuf_5_7_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_14__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_28741_ _34688_/Q _27165_/X _28755_/S VGND VGND VPWR VPWR _28742_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25953_ _24806_/X _33432_/Q _25967_/S VGND VGND VPWR VPWR _25954_/A sky130_fd_sc_hd__mux2_1
X_21076_ _21072_/X _21075_/X _21034_/X _21035_/X VGND VGND VPWR VPWR _21091_/B sky130_fd_sc_hd__o211a_1
XFILLER_63_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20027_ _34181_/Q _34117_/Q _34053_/Q _33989_/Q _19746_/X _19747_/X VGND VGND VPWR
+ VPWR _20027_/X sky130_fd_sc_hd__mux4_1
X_24904_ _24904_/A VGND VGND VPWR VPWR _32951_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_219_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28672_ _28672_/A VGND VGND VPWR VPWR _34655_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25884_ _25884_/A VGND VGND VPWR VPWR _33399_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27623_ _34190_/Q _27208_/X _27629_/S VGND VGND VPWR VPWR _27624_/A sky130_fd_sc_hd__mux2_1
X_24835_ _24834_/X _32929_/Q _24859_/S VGND VGND VPWR VPWR _24836_/A sky130_fd_sc_hd__mux2_1
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27554_ _34157_/Q _27106_/X _27566_/S VGND VGND VPWR VPWR _27555_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24766_ _24766_/A VGND VGND VPWR VPWR _32903_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21978_ _22451_/A VGND VGND VPWR VPWR _21978_/X sky130_fd_sc_hd__buf_6
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_1090 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26505_ _24821_/X _33693_/Q _26509_/S VGND VGND VPWR VPWR _26506_/A sky130_fd_sc_hd__mux2_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23717_ _22900_/X _32346_/Q _23727_/S VGND VGND VPWR VPWR _23718_/A sky130_fd_sc_hd__mux2_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27485_ _27485_/A VGND VGND VPWR VPWR _34124_/D sky130_fd_sc_hd__clkbuf_1
X_20929_ _20925_/X _20928_/X _20644_/X _20646_/X VGND VGND VPWR VPWR _20944_/B sky130_fd_sc_hd__o211a_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24697_ _24697_/A VGND VGND VPWR VPWR _32870_/D sky130_fd_sc_hd__clkbuf_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29224_ _34916_/Q _27078_/X _29234_/S VGND VGND VPWR VPWR _29225_/A sky130_fd_sc_hd__mux2_1
X_26436_ _33661_/Q _23417_/X _26436_/S VGND VGND VPWR VPWR _26437_/A sky130_fd_sc_hd__mux2_1
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23648_ _23002_/X _32315_/Q _23652_/S VGND VGND VPWR VPWR _23649_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29155_ _29155_/A VGND VGND VPWR VPWR _34883_/D sky130_fd_sc_hd__clkbuf_1
X_26367_ _33628_/Q _23249_/X _26373_/S VGND VGND VPWR VPWR _26368_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_195_CLK clkbuf_6_49__f_CLK/X VGND VGND VPWR VPWR _35853_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_211_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23579_ _22900_/X _32282_/Q _23589_/S VGND VGND VPWR VPWR _23580_/A sky130_fd_sc_hd__mux2_1
X_16120_ _32087_/Q _32279_/Q _32343_/Q _35863_/Q _16032_/X _17867_/A VGND VGND VPWR
+ VPWR _16120_/X sky130_fd_sc_hd__mux4_1
XFILLER_195_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28106_ _34388_/Q _27226_/X _28108_/S VGND VGND VPWR VPWR _28107_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25318_ _33132_/Q _23299_/X _25332_/S VGND VGND VPWR VPWR _25319_/A sky130_fd_sc_hd__mux2_1
X_29086_ _29086_/A VGND VGND VPWR VPWR _34850_/D sky130_fd_sc_hd__clkbuf_1
X_26298_ _24917_/X _33596_/Q _26300_/S VGND VGND VPWR VPWR _26299_/A sky130_fd_sc_hd__mux2_1
X_16051_ _35670_/Q _32175_/Q _35542_/Q _35478_/Q _16049_/X _16050_/X VGND VGND VPWR
+ VPWR _16051_/X sky130_fd_sc_hd__mux4_1
X_28037_ _34355_/Q _27124_/X _28037_/S VGND VGND VPWR VPWR _28038_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25249_ _33100_/Q _23469_/X _25259_/S VGND VGND VPWR VPWR _25250_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1050 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19810_ _19806_/X _19807_/X _19808_/X _19809_/X VGND VGND VPWR VPWR _19810_/X sky130_fd_sc_hd__a22o_1
XFILLER_237_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29988_ _35248_/Q _29410_/X _29994_/S VGND VGND VPWR VPWR _29989_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16953_ _33391_/Q _33327_/Q _33263_/Q _33199_/Q _16774_/X _16775_/X VGND VGND VPWR
+ VPWR _16953_/X sky130_fd_sc_hd__mux4_1
X_19741_ _19458_/X _19739_/X _19740_/X _19463_/X VGND VGND VPWR VPWR _19741_/X sky130_fd_sc_hd__a22o_1
X_28939_ _34781_/Q _27056_/X _28943_/S VGND VGND VPWR VPWR _28940_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31950_ _23487_/X _36178_/Q _31956_/S VGND VGND VPWR VPWR _31951_/A sky130_fd_sc_hd__mux2_1
X_19672_ _19672_/A VGND VGND VPWR VPWR _32442_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_237_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16884_ _33645_/Q _33581_/Q _33517_/Q _33453_/Q _16847_/X _16848_/X VGND VGND VPWR
+ VPWR _16884_/X sky130_fd_sc_hd__mux4_1
XFILLER_42_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18623_ _32605_/Q _32541_/Q _32477_/Q _35933_/Q _18517_/X _20017_/A VGND VGND VPWR
+ VPWR _18623_/X sky130_fd_sc_hd__mux4_1
XFILLER_37_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30901_ _30901_/A VGND VGND VPWR VPWR _35680_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_237_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31881_ _23364_/X _36145_/Q _31885_/S VGND VGND VPWR VPWR _31882_/A sky130_fd_sc_hd__mux2_1
XFILLER_237_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33620_ _33685_/CLK _33620_/D VGND VGND VPWR VPWR _33620_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18554_ _32091_/Q _32283_/Q _32347_/Q _35867_/Q _18521_/X _20167_/A VGND VGND VPWR
+ VPWR _18554_/X sky130_fd_sc_hd__mux4_1
X_30832_ _35648_/Q input37/X _30846_/S VGND VGND VPWR VPWR _30833_/A sky130_fd_sc_hd__mux2_1
XTAP_3470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17505_ _17500_/X _17503_/X _17504_/X VGND VGND VPWR VPWR _17520_/C sky130_fd_sc_hd__o21ba_1
XTAP_3492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33551_ _34441_/CLK _33551_/D VGND VGND VPWR VPWR _33551_/Q sky130_fd_sc_hd__dfxtp_1
X_18485_ _32601_/Q _32537_/Q _32473_/Q _35929_/Q _20166_/A _20017_/A VGND VGND VPWR
+ VPWR _18485_/X sky130_fd_sc_hd__mux4_1
X_30763_ _30763_/A VGND VGND VPWR VPWR _35615_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_206_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32502_ _36021_/CLK _32502_/D VGND VGND VPWR VPWR _32502_/Q sky130_fd_sc_hd__dfxtp_1
X_17436_ _34684_/Q _34620_/Q _34556_/Q _34492_/Q _17292_/X _17293_/X VGND VGND VPWR
+ VPWR _17436_/X sky130_fd_sc_hd__mux4_1
X_33482_ _33869_/CLK _33482_/D VGND VGND VPWR VPWR _33482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30694_ _30694_/A VGND VGND VPWR VPWR _35582_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_242_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35221_ _35221_/CLK _35221_/D VGND VGND VPWR VPWR _35221_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_1464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32433_ _33895_/CLK _32433_/D VGND VGND VPWR VPWR _32433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_186_CLK clkbuf_leaf_65_CLK/A VGND VGND VPWR VPWR _36049_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_144_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17367_ _34426_/Q _36154_/Q _34298_/Q _34234_/Q _17229_/X _17230_/X VGND VGND VPWR
+ VPWR _17367_/X sky130_fd_sc_hd__mux4_1
XFILLER_14_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19106_ _34410_/Q _36138_/Q _34282_/Q _34218_/Q _18823_/X _18824_/X VGND VGND VPWR
+ VPWR _19106_/X sky130_fd_sc_hd__mux4_1
X_35152_ _36115_/CLK _35152_/D VGND VGND VPWR VPWR _35152_/Q sky130_fd_sc_hd__dfxtp_1
X_16318_ _17850_/A VGND VGND VPWR VPWR _16318_/X sky130_fd_sc_hd__buf_6
XFILLER_140_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32364_ _35949_/CLK _32364_/D VGND VGND VPWR VPWR _32364_/Q sky130_fd_sc_hd__dfxtp_1
X_17298_ _34936_/Q _34872_/Q _34808_/Q _34744_/Q _17160_/X _17161_/X VGND VGND VPWR
+ VPWR _17298_/X sky130_fd_sc_hd__mux4_1
X_34103_ _35704_/CLK _34103_/D VGND VGND VPWR VPWR _34103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19037_ _19037_/A _19037_/B _19037_/C _19037_/D VGND VGND VPWR VPWR _19038_/A sky130_fd_sc_hd__or4_2
X_31315_ _31315_/A VGND VGND VPWR VPWR _35876_/D sky130_fd_sc_hd__clkbuf_1
X_35083_ _35212_/CLK _35083_/D VGND VGND VPWR VPWR _35083_/Q sky130_fd_sc_hd__dfxtp_1
X_16249_ _16147_/X _16247_/X _16248_/X _16150_/X VGND VGND VPWR VPWR _16249_/X sky130_fd_sc_hd__a22o_1
X_32295_ _35947_/CLK _32295_/D VGND VGND VPWR VPWR _32295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput102 _31978_/Q VGND VGND VPWR VPWR D1[20] sky130_fd_sc_hd__buf_2
XFILLER_86_1131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34034_ _35635_/CLK _34034_/D VGND VGND VPWR VPWR _34034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput113 _31988_/Q VGND VGND VPWR VPWR D1[30] sky130_fd_sc_hd__buf_2
X_31246_ _27785_/X _35844_/Q _31252_/S VGND VGND VPWR VPWR _31247_/A sky130_fd_sc_hd__mux2_1
Xoutput124 _31998_/Q VGND VGND VPWR VPWR D1[40] sky130_fd_sc_hd__buf_2
XFILLER_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput135 _32008_/Q VGND VGND VPWR VPWR D1[50] sky130_fd_sc_hd__buf_2
XFILLER_99_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput146 _32018_/Q VGND VGND VPWR VPWR D1[60] sky130_fd_sc_hd__buf_2
Xoutput157 _36194_/Q VGND VGND VPWR VPWR D2[12] sky130_fd_sc_hd__buf_2
XFILLER_142_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput168 _36204_/Q VGND VGND VPWR VPWR D2[22] sky130_fd_sc_hd__buf_2
Xoutput179 _36214_/Q VGND VGND VPWR VPWR D2[32] sky130_fd_sc_hd__buf_2
XFILLER_130_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31177_ _27683_/X _35811_/Q _31189_/S VGND VGND VPWR VPWR _31178_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30128_ _30128_/A VGND VGND VPWR VPWR _35314_/D sky130_fd_sc_hd__clkbuf_1
X_19939_ _35650_/Q _35010_/Q _34370_/Q _33730_/Q _19797_/X _19798_/X VGND VGND VPWR
+ VPWR _19939_/X sky130_fd_sc_hd__mux4_1
X_35985_ _35985_/CLK _35985_/D VGND VGND VPWR VPWR _35985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_110_CLK clkbuf_6_22__f_CLK/X VGND VGND VPWR VPWR _35801_/CLK sky130_fd_sc_hd__clkbuf_16
X_30059_ _35282_/Q _29515_/X _30065_/S VGND VGND VPWR VPWR _30060_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34936_ _36152_/CLK _34936_/D VGND VGND VPWR VPWR _34936_/Q sky130_fd_sc_hd__dfxtp_1
X_22950_ _23083_/S VGND VGND VPWR VPWR _22978_/S sky130_fd_sc_hd__buf_4
XFILLER_229_878 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21901_ _21901_/A _21901_/B _21901_/C _21901_/D VGND VGND VPWR VPWR _21902_/A sky130_fd_sc_hd__or4_1
XFILLER_228_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_5_8_0_CLK clkbuf_5_9_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_8_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_95_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22881_ _22881_/A VGND VGND VPWR VPWR _31147_/A sky130_fd_sc_hd__buf_8
X_34867_ _35056_/CLK _34867_/D VGND VGND VPWR VPWR _34867_/Q sky130_fd_sc_hd__dfxtp_1
X_24620_ _23024_/X _32834_/Q _24630_/S VGND VGND VPWR VPWR _24621_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33818_ _33818_/CLK _33818_/D VGND VGND VPWR VPWR _33818_/Q sky130_fd_sc_hd__dfxtp_1
X_21832_ _34934_/Q _34870_/Q _34806_/Q _34742_/Q _21760_/X _21761_/X VGND VGND VPWR
+ VPWR _21832_/X sky130_fd_sc_hd__mux4_1
XFILLER_83_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34798_ _35183_/CLK _34798_/D VGND VGND VPWR VPWR _34798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24551_ _22922_/X _32801_/Q _24567_/S VGND VGND VPWR VPWR _24552_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21763_ _21763_/A VGND VGND VPWR VPWR _21763_/X sky130_fd_sc_hd__buf_4
XFILLER_224_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33749_ _35669_/CLK _33749_/D VGND VGND VPWR VPWR _33749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_1277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20714_ _33879_/Q _33815_/Q _33751_/Q _36055_/Q _20712_/X _20713_/X VGND VGND VPWR
+ VPWR _20714_/X sky130_fd_sc_hd__mux4_1
XFILLER_169_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23502_ _23502_/A VGND VGND VPWR VPWR _32246_/D sky130_fd_sc_hd__clkbuf_1
X_27270_ _27270_/A VGND VGND VPWR VPWR _34022_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24482_ _24482_/A VGND VGND VPWR VPWR _32768_/D sky130_fd_sc_hd__clkbuf_1
X_21694_ _22561_/A VGND VGND VPWR VPWR _21694_/X sky130_fd_sc_hd__buf_4
XFILLER_52_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26221_ _24803_/X _33559_/Q _26237_/S VGND VGND VPWR VPWR _26222_/A sky130_fd_sc_hd__mux2_1
XFILLER_221_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35419_ _36059_/CLK _35419_/D VGND VGND VPWR VPWR _35419_/Q sky130_fd_sc_hd__dfxtp_1
X_20645_ input76/X VGND VGND VPWR VPWR _22447_/A sky130_fd_sc_hd__buf_6
X_23433_ _32223_/Q _23432_/X _23451_/S VGND VGND VPWR VPWR _23434_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_177_CLK clkbuf_6_27__f_CLK/X VGND VGND VPWR VPWR _35858_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_137_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26152_ _26152_/A VGND VGND VPWR VPWR _33526_/D sky130_fd_sc_hd__clkbuf_1
X_23364_ input20/X VGND VGND VPWR VPWR _23364_/X sky130_fd_sc_hd__buf_4
X_20576_ _20572_/X _20575_/X _20171_/A VGND VGND VPWR VPWR _20577_/D sky130_fd_sc_hd__o21ba_1
XFILLER_137_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25103_ _25130_/S VGND VGND VPWR VPWR _25122_/S sky130_fd_sc_hd__buf_4
XFILLER_30_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22315_ _34692_/Q _34628_/Q _34564_/Q _34500_/Q _22245_/X _22246_/X VGND VGND VPWR
+ VPWR _22315_/X sky130_fd_sc_hd__mux4_1
XFILLER_194_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26083_ _26215_/S VGND VGND VPWR VPWR _26102_/S sky130_fd_sc_hd__buf_6
X_23295_ _23295_/A VGND VGND VPWR VPWR _32170_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29911_ _29911_/A VGND VGND VPWR VPWR _35211_/D sky130_fd_sc_hd__clkbuf_1
X_22246_ _22599_/A VGND VGND VPWR VPWR _22246_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_180_847 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25034_ _24852_/X _32999_/Q _25038_/S VGND VGND VPWR VPWR _25035_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_1354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29842_ _29842_/A VGND VGND VPWR VPWR _35178_/D sky130_fd_sc_hd__clkbuf_1
X_22177_ _21956_/X _22175_/X _22176_/X _21959_/X VGND VGND VPWR VPWR _22177_/X sky130_fd_sc_hd__a22o_1
XFILLER_191_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_1086 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21128_ _21122_/X _21127_/X _21059_/X VGND VGND VPWR VPWR _21129_/D sky130_fd_sc_hd__o21ba_1
X_29773_ _35146_/Q _29491_/X _29787_/S VGND VGND VPWR VPWR _29774_/A sky130_fd_sc_hd__mux2_1
X_26985_ _26985_/A VGND VGND VPWR VPWR _33918_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28724_ _34680_/Q _27140_/X _28734_/S VGND VGND VPWR VPWR _28725_/A sky130_fd_sc_hd__mux2_1
X_25936_ _25936_/A VGND VGND VPWR VPWR _33424_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_101_CLK clkbuf_leaf_99_CLK/A VGND VGND VPWR VPWR _36212_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_4_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21059_ _22471_/A VGND VGND VPWR VPWR _21059_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_19_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28655_ _34647_/Q _27038_/X _28671_/S VGND VGND VPWR VPWR _28656_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25867_ _25867_/A VGND VGND VPWR VPWR _33391_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27606_ _34182_/Q _27183_/X _27608_/S VGND VGND VPWR VPWR _27607_/A sky130_fd_sc_hd__mux2_1
XFILLER_189_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24818_ input61/X VGND VGND VPWR VPWR _24818_/X sky130_fd_sc_hd__buf_2
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28586_ _27745_/X _34615_/Q _28598_/S VGND VGND VPWR VPWR _28587_/A sky130_fd_sc_hd__mux2_1
X_25798_ _24976_/X _33359_/Q _25802_/S VGND VGND VPWR VPWR _25799_/A sky130_fd_sc_hd__mux2_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_931 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27537_ _34149_/Q _27081_/X _27545_/S VGND VGND VPWR VPWR _27538_/A sky130_fd_sc_hd__mux2_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24749_ _23015_/X _32895_/Q _24765_/S VGND VGND VPWR VPWR _24750_/A sky130_fd_sc_hd__mux2_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18270_ _34709_/Q _34645_/Q _34581_/Q _34517_/Q _17998_/X _17999_/X VGND VGND VPWR
+ VPWR _18270_/X sky130_fd_sc_hd__mux4_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27468_ _27468_/A VGND VGND VPWR VPWR _34116_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_226_1057 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29207_ _34908_/Q _27053_/X _29213_/S VGND VGND VPWR VPWR _29208_/A sky130_fd_sc_hd__mux2_1
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17221_ _16998_/X _17219_/X _17220_/X _17001_/X VGND VGND VPWR VPWR _17221_/X sky130_fd_sc_hd__a22o_1
X_26419_ _26419_/A VGND VGND VPWR VPWR _33652_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1041 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_168_CLK clkbuf_6_30__f_CLK/X VGND VGND VPWR VPWR _36114_/CLK sky130_fd_sc_hd__clkbuf_16
X_27399_ _27399_/A VGND VGND VPWR VPWR _34083_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17152_ _17147_/X _17150_/X _17151_/X VGND VGND VPWR VPWR _17167_/C sky130_fd_sc_hd__o21ba_1
X_29138_ _29138_/A VGND VGND VPWR VPWR _34875_/D sky130_fd_sc_hd__clkbuf_1
Xinput15 DW[22] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__buf_4
XFILLER_11_883 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput26 DW[32] VGND VGND VPWR VPWR input26/X sky130_fd_sc_hd__clkbuf_4
XFILLER_122_1055 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput37 DW[42] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__buf_6
X_16103_ input70/X input69/X VGND VGND VPWR VPWR _17871_/A sky130_fd_sc_hd__or2b_4
Xinput48 DW[52] VGND VGND VPWR VPWR input48/X sky130_fd_sc_hd__buf_8
Xinput59 DW[62] VGND VGND VPWR VPWR input59/X sky130_fd_sc_hd__clkbuf_16
X_29069_ _29069_/A VGND VGND VPWR VPWR _34842_/D sky130_fd_sc_hd__clkbuf_1
X_17083_ _34674_/Q _34610_/Q _34546_/Q _34482_/Q _16939_/X _16940_/X VGND VGND VPWR
+ VPWR _17083_/X sky130_fd_sc_hd__mux4_1
XFILLER_157_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31100_ _35775_/Q input36/X _31116_/S VGND VGND VPWR VPWR _31101_/A sky130_fd_sc_hd__mux2_1
X_16034_ _17774_/A VGND VGND VPWR VPWR _17867_/A sky130_fd_sc_hd__buf_8
XFILLER_109_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32080_ _35855_/CLK _32080_/D VGND VGND VPWR VPWR _32080_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31031_ _31031_/A VGND VGND VPWR VPWR _35742_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_233_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_340_CLK clkbuf_6_45__f_CLK/X VGND VGND VPWR VPWR _32891_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_112_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17985_ _17765_/X _17983_/X _17984_/X _17771_/X VGND VGND VPWR VPWR _17985_/X sky130_fd_sc_hd__a22o_1
XFILLER_123_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19724_ _20215_/A VGND VGND VPWR VPWR _19724_/X sky130_fd_sc_hd__clkbuf_4
X_16936_ _33070_/Q _32046_/Q _35822_/Q _35758_/Q _16725_/X _16726_/X VGND VGND VPWR
+ VPWR _16936_/X sky130_fd_sc_hd__mux4_1
XFILLER_96_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32982_ _35992_/CLK _32982_/D VGND VGND VPWR VPWR _32982_/Q sky130_fd_sc_hd__dfxtp_1
X_35770_ _35835_/CLK _35770_/D VGND VGND VPWR VPWR _35770_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_6_60__f_CLK clkbuf_5_30_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_60__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_37_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34721_ _34915_/CLK _34721_/D VGND VGND VPWR VPWR _34721_/Q sky130_fd_sc_hd__dfxtp_1
X_31933_ _31933_/A VGND VGND VPWR VPWR _36169_/D sky130_fd_sc_hd__clkbuf_1
X_16867_ _35628_/Q _34988_/Q _34348_/Q _33708_/Q _16791_/X _16792_/X VGND VGND VPWR
+ VPWR _16867_/X sky130_fd_sc_hd__mux4_1
X_19655_ _19651_/X _19652_/X _19653_/X _19654_/X VGND VGND VPWR VPWR _19655_/X sky130_fd_sc_hd__a22o_1
XFILLER_93_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_226_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18606_ _35164_/Q _35100_/Q _35036_/Q _32156_/Q _18604_/X _18605_/X VGND VGND VPWR
+ VPWR _18606_/X sky130_fd_sc_hd__mux4_1
X_34652_ _36229_/CLK _34652_/D VGND VGND VPWR VPWR _34652_/Q sky130_fd_sc_hd__dfxtp_1
X_19586_ _35640_/Q _35000_/Q _34360_/Q _33720_/Q _19444_/X _19445_/X VGND VGND VPWR
+ VPWR _19586_/X sky130_fd_sc_hd__mux4_1
X_31864_ _23289_/X _36137_/Q _31864_/S VGND VGND VPWR VPWR _31865_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16798_ _17857_/A VGND VGND VPWR VPWR _16798_/X sky130_fd_sc_hd__buf_2
XFILLER_20_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33603_ _34180_/CLK _33603_/D VGND VGND VPWR VPWR _33603_/Q sky130_fd_sc_hd__dfxtp_1
X_18537_ _18378_/X _18535_/X _18536_/X _18388_/X VGND VGND VPWR VPWR _18537_/X sky130_fd_sc_hd__a22o_1
X_30815_ _35640_/Q input28/X _30825_/S VGND VGND VPWR VPWR _30816_/A sky130_fd_sc_hd__mux2_1
XFILLER_244_1113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34583_ _34647_/CLK _34583_/D VGND VGND VPWR VPWR _34583_/Q sky130_fd_sc_hd__dfxtp_1
X_31795_ _36104_/Q input46/X _31813_/S VGND VGND VPWR VPWR _31796_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18468_ _35160_/Q _35096_/Q _35032_/Q _32152_/Q _18383_/X _18385_/X VGND VGND VPWR
+ VPWR _18468_/X sky130_fd_sc_hd__mux4_1
X_30746_ _35607_/Q input12/X _30762_/S VGND VGND VPWR VPWR _30747_/A sky130_fd_sc_hd__mux2_1
X_33534_ _35453_/CLK _33534_/D VGND VGND VPWR VPWR _33534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17419_ _17412_/X _17414_/X _17417_/X _17418_/X VGND VGND VPWR VPWR _17419_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_159_CLK clkbuf_6_31__f_CLK/X VGND VGND VPWR VPWR _36175_/CLK sky130_fd_sc_hd__clkbuf_16
X_33465_ _33913_/CLK _33465_/D VGND VGND VPWR VPWR _33465_/Q sky130_fd_sc_hd__dfxtp_1
X_18399_ _34902_/Q _34838_/Q _34774_/Q _34710_/Q _18396_/X _18398_/X VGND VGND VPWR
+ VPWR _18399_/X sky130_fd_sc_hd__mux4_1
X_30677_ _30677_/A VGND VGND VPWR VPWR _35574_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_991 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20430_ _34193_/Q _34129_/Q _34065_/Q _34001_/Q _18349_/X _18350_/X VGND VGND VPWR
+ VPWR _20430_/X sky130_fd_sc_hd__mux4_1
X_35204_ _35717_/CLK _35204_/D VGND VGND VPWR VPWR _35204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32416_ _33573_/CLK _32416_/D VGND VGND VPWR VPWR _32416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36184_ _36191_/CLK _36184_/D VGND VGND VPWR VPWR _36184_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33396_ _34100_/CLK _33396_/D VGND VGND VPWR VPWR _33396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20361_ _35214_/Q _35150_/Q _35086_/Q _32270_/Q _18392_/X _18394_/X VGND VGND VPWR
+ VPWR _20361_/X sky130_fd_sc_hd__mux4_1
X_35135_ _36100_/CLK _35135_/D VGND VGND VPWR VPWR _35135_/Q sky130_fd_sc_hd__dfxtp_1
X_32347_ _35995_/CLK _32347_/D VGND VGND VPWR VPWR _32347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22100_ _21951_/X _22096_/X _22099_/X _21954_/X VGND VGND VPWR VPWR _22100_/X sky130_fd_sc_hd__a22o_1
XFILLER_134_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23080_ _23079_/X _32084_/Q _23083_/S VGND VGND VPWR VPWR _23081_/A sky130_fd_sc_hd__mux2_1
X_35066_ _35194_/CLK _35066_/D VGND VGND VPWR VPWR _35066_/Q sky130_fd_sc_hd__dfxtp_1
X_32278_ _35221_/CLK _32278_/D VGND VGND VPWR VPWR _32278_/Q sky130_fd_sc_hd__dfxtp_1
X_20292_ _35660_/Q _35020_/Q _34380_/Q _33740_/Q _20150_/X _20151_/X VGND VGND VPWR
+ VPWR _20292_/X sky130_fd_sc_hd__mux4_1
XFILLER_164_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22031_ _22535_/A VGND VGND VPWR VPWR _22031_/X sky130_fd_sc_hd__buf_6
X_34017_ _34594_/CLK _34017_/D VGND VGND VPWR VPWR _34017_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31229_ _27760_/X _35836_/Q _31231_/S VGND VGND VPWR VPWR _31230_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_331_CLK clkbuf_6_38__f_CLK/X VGND VGND VPWR VPWR _36023_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_88_614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26770_ _26770_/A VGND VGND VPWR VPWR _33816_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23982_ _22879_/X _32534_/Q _24000_/S VGND VGND VPWR VPWR _23983_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35968_ _36030_/CLK _35968_/D VGND VGND VPWR VPWR _35968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25721_ _24861_/X _33322_/Q _25739_/S VGND VGND VPWR VPWR _25722_/A sky130_fd_sc_hd__mux2_1
XFILLER_228_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34919_ _34921_/CLK _34919_/D VGND VGND VPWR VPWR _34919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22933_ _22933_/A VGND VGND VPWR VPWR _32036_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_216_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35899_ _36027_/CLK _35899_/D VGND VGND VPWR VPWR _35899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28440_ _27729_/X _34546_/Q _28442_/S VGND VGND VPWR VPWR _28441_/A sky130_fd_sc_hd__mux2_1
X_25652_ _25652_/A VGND VGND VPWR VPWR _33289_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22864_ _35669_/Q _35029_/Q _34389_/Q _33749_/Q _20712_/X _20713_/X VGND VGND VPWR
+ VPWR _22864_/X sky130_fd_sc_hd__mux4_1
XFILLER_37_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24603_ _22999_/X _32826_/Q _24609_/S VGND VGND VPWR VPWR _24604_/A sky130_fd_sc_hd__mux2_1
XFILLER_227_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28371_ _28371_/A VGND VGND VPWR VPWR _34513_/D sky130_fd_sc_hd__clkbuf_1
X_21815_ _32118_/Q _32310_/Q _32374_/Q _35894_/Q _21527_/X _21668_/X VGND VGND VPWR
+ VPWR _21815_/X sky130_fd_sc_hd__mux4_1
XFILLER_25_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25583_ _24858_/X _33257_/Q _25583_/S VGND VGND VPWR VPWR _25584_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_398_CLK clkbuf_6_35__f_CLK/X VGND VGND VPWR VPWR _35126_/CLK sky130_fd_sc_hd__clkbuf_16
X_22795_ _22791_/X _22794_/X _22438_/A VGND VGND VPWR VPWR _22817_/A sky130_fd_sc_hd__o21ba_1
XPHY_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27322_ _34047_/Q _27162_/X _27338_/S VGND VGND VPWR VPWR _27323_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24534_ _22897_/X _32793_/Q _24546_/S VGND VGND VPWR VPWR _24535_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21746_ _35636_/Q _34996_/Q _34356_/Q _33716_/Q _21744_/X _21745_/X VGND VGND VPWR
+ VPWR _21746_/X sky130_fd_sc_hd__mux4_1
XFILLER_40_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27253_ _27253_/A VGND VGND VPWR VPWR _34014_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_185_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24465_ _24465_/A VGND VGND VPWR VPWR _32760_/D sky130_fd_sc_hd__clkbuf_1
X_21677_ _35442_/Q _35378_/Q _35314_/Q _35250_/Q _21501_/X _21502_/X VGND VGND VPWR
+ VPWR _21677_/X sky130_fd_sc_hd__mux4_1
XFILLER_225_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26204_ _26204_/A VGND VGND VPWR VPWR _33551_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23416_ _23416_/A VGND VGND VPWR VPWR _32217_/D sky130_fd_sc_hd__clkbuf_1
X_27184_ _33990_/Q _27183_/X _27187_/S VGND VGND VPWR VPWR _27185_/A sky130_fd_sc_hd__mux2_1
X_20628_ _20618_/X _20623_/X _20626_/X _20627_/X VGND VGND VPWR VPWR _20628_/X sky130_fd_sc_hd__a22o_1
X_24396_ _24396_/A VGND VGND VPWR VPWR _32727_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26135_ _26135_/A VGND VGND VPWR VPWR _33518_/D sky130_fd_sc_hd__clkbuf_1
X_20559_ _32149_/Q _32341_/Q _32405_/Q _35925_/Q _20286_/X _19311_/A VGND VGND VPWR
+ VPWR _20559_/X sky130_fd_sc_hd__mux4_1
XFILLER_125_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23347_ _32190_/Q _23271_/X _23359_/S VGND VGND VPWR VPWR _23348_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26066_ _24973_/X _33486_/Q _26072_/S VGND VGND VPWR VPWR _26067_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23278_ _32165_/Q _23277_/X _23290_/S VGND VGND VPWR VPWR _23279_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25017_ _24827_/X _32991_/Q _25017_/S VGND VGND VPWR VPWR _25018_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22229_ _22582_/A VGND VGND VPWR VPWR _22229_/X sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_322_CLK clkbuf_6_39__f_CLK/X VGND VGND VPWR VPWR _32904_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_6810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_880 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29825_ _29825_/A VGND VGND VPWR VPWR _35170_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17770_ _33158_/Q _36038_/Q _33030_/Q _32966_/Q _17768_/X _17769_/X VGND VGND VPWR
+ VPWR _17770_/X sky130_fd_sc_hd__mux4_1
XFILLER_43_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29756_ _35138_/Q _29466_/X _29766_/S VGND VGND VPWR VPWR _29757_/A sky130_fd_sc_hd__mux2_1
X_26968_ _26968_/A VGND VGND VPWR VPWR _33910_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16721_ _35688_/Q _32195_/Q _35560_/Q _35496_/Q _16611_/X _16612_/X VGND VGND VPWR
+ VPWR _16721_/X sky130_fd_sc_hd__mux4_1
X_25919_ _24954_/X _33416_/Q _25937_/S VGND VGND VPWR VPWR _25920_/A sky130_fd_sc_hd__mux2_1
X_28707_ _34672_/Q _27115_/X _28713_/S VGND VGND VPWR VPWR _28708_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29687_ _35105_/Q _29364_/X _29703_/S VGND VGND VPWR VPWR _29688_/A sky130_fd_sc_hd__mux2_1
X_26899_ _27031_/S VGND VGND VPWR VPWR _26918_/S sky130_fd_sc_hd__buf_6
XFILLER_86_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19440_ _20146_/A VGND VGND VPWR VPWR _19440_/X sky130_fd_sc_hd__clkbuf_4
X_28638_ _27822_/X _34640_/Q _28640_/S VGND VGND VPWR VPWR _28639_/A sky130_fd_sc_hd__mux2_1
X_16652_ _33062_/Q _32038_/Q _35814_/Q _35750_/Q _16372_/X _16373_/X VGND VGND VPWR
+ VPWR _16652_/X sky130_fd_sc_hd__mux4_1
XFILLER_235_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19371_ _20215_/A VGND VGND VPWR VPWR _19371_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_389_CLK clkbuf_6_40__f_CLK/X VGND VGND VPWR VPWR _33911_/CLK sky130_fd_sc_hd__clkbuf_16
X_28569_ _27720_/X _34607_/Q _28577_/S VGND VGND VPWR VPWR _28570_/A sky130_fd_sc_hd__mux2_1
X_16583_ _33060_/Q _32036_/Q _35812_/Q _35748_/Q _16372_/X _16373_/X VGND VGND VPWR
+ VPWR _16583_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30600_ _30600_/A VGND VGND VPWR VPWR _35538_/D sky130_fd_sc_hd__clkbuf_1
X_18322_ _20066_/A VGND VGND VPWR VPWR _20017_/A sky130_fd_sc_hd__buf_8
XFILLER_15_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31580_ _27680_/X _36002_/Q _31594_/S VGND VGND VPWR VPWR _31581_/A sky130_fd_sc_hd__mux2_1
XFILLER_187_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18253_ _33941_/Q _33877_/Q _33813_/Q _36117_/Q _16062_/X _16064_/X VGND VGND VPWR
+ VPWR _18253_/X sky130_fd_sc_hd__mux4_1
XFILLER_124_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30531_ _30531_/A VGND VGND VPWR VPWR _35505_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17204_ _17910_/A VGND VGND VPWR VPWR _17204_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_187_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33250_ _33827_/CLK _33250_/D VGND VGND VPWR VPWR _33250_/Q sky130_fd_sc_hd__dfxtp_1
X_18184_ _34962_/Q _34898_/Q _34834_/Q _34770_/Q _16083_/X _16085_/X VGND VGND VPWR
+ VPWR _18184_/X sky130_fd_sc_hd__mux4_1
XFILLER_175_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30462_ _35473_/Q _29512_/X _30462_/S VGND VGND VPWR VPWR _30463_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32201_ _35693_/CLK _32201_/D VGND VGND VPWR VPWR _32201_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17135_ _33140_/Q _36020_/Q _33012_/Q _32948_/Q _17062_/X _17063_/X VGND VGND VPWR
+ VPWR _17135_/X sky130_fd_sc_hd__mux4_1
X_33181_ _36205_/CLK _33181_/D VGND VGND VPWR VPWR _33181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30393_ _35440_/Q _29410_/X _30399_/S VGND VGND VPWR VPWR _30394_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32132_ _35973_/CLK _32132_/D VGND VGND VPWR VPWR _32132_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17066_ _17059_/X _17061_/X _17064_/X _17065_/X VGND VGND VPWR VPWR _17066_/X sky130_fd_sc_hd__a22o_1
XFILLER_170_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16017_ _17765_/A VGND VGND VPWR VPWR _17905_/A sky130_fd_sc_hd__buf_12
XFILLER_100_1172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32063_ _35454_/CLK _32063_/D VGND VGND VPWR VPWR _32063_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_313_CLK clkbuf_6_48__f_CLK/X VGND VGND VPWR VPWR _36040_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_98_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31014_ _35734_/Q input1/X _31032_/S VGND VGND VPWR VPWR _31015_/A sky130_fd_sc_hd__mux2_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_1115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35822_ _35822_/CLK _35822_/D VGND VGND VPWR VPWR _35822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17968_ _17859_/X _17966_/X _17967_/X _17862_/X VGND VGND VPWR VPWR _17968_/X sky130_fd_sc_hd__a22o_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19707_ _19499_/X _19705_/X _19706_/X _19504_/X VGND VGND VPWR VPWR _19707_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16919_ _33390_/Q _33326_/Q _33262_/Q _33198_/Q _16774_/X _16775_/X VGND VGND VPWR
+ VPWR _16919_/X sky130_fd_sc_hd__mux4_1
X_35753_ _35753_/CLK _35753_/D VGND VGND VPWR VPWR _35753_/Q sky130_fd_sc_hd__dfxtp_1
X_32965_ _36037_/CLK _32965_/D VGND VGND VPWR VPWR _32965_/Q sky130_fd_sc_hd__dfxtp_1
X_17899_ _34441_/Q _36169_/Q _34313_/Q _34249_/Q _17582_/X _17583_/X VGND VGND VPWR
+ VPWR _17899_/X sky130_fd_sc_hd__mux4_1
X_34704_ _34705_/CLK _34704_/D VGND VGND VPWR VPWR _34704_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31916_ _31916_/A VGND VGND VPWR VPWR _36161_/D sky130_fd_sc_hd__clkbuf_1
X_19638_ _33402_/Q _33338_/Q _33274_/Q _33210_/Q _19427_/X _19428_/X VGND VGND VPWR
+ VPWR _19638_/X sky130_fd_sc_hd__mux4_1
X_35684_ _35684_/CLK _35684_/D VGND VGND VPWR VPWR _35684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32896_ _32896_/CLK _32896_/D VGND VGND VPWR VPWR _32896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_829 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34635_ _35208_/CLK _34635_/D VGND VGND VPWR VPWR _34635_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31847_ _31847_/A VGND VGND VPWR VPWR _36128_/D sky130_fd_sc_hd__clkbuf_1
X_19569_ _33656_/Q _33592_/Q _33528_/Q _33464_/Q _19500_/X _19501_/X VGND VGND VPWR
+ VPWR _19569_/X sky130_fd_sc_hd__mux4_1
XFILLER_18_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21600_ _35632_/Q _34992_/Q _34352_/Q _33712_/Q _21391_/X _21392_/X VGND VGND VPWR
+ VPWR _21600_/X sky130_fd_sc_hd__mux4_1
XFILLER_55_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22580_ _22512_/X _22578_/X _22579_/X _22515_/X VGND VGND VPWR VPWR _22580_/X sky130_fd_sc_hd__a22o_1
XFILLER_209_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34566_ _34694_/CLK _34566_/D VGND VGND VPWR VPWR _34566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31778_ _36096_/Q input37/X _31792_/S VGND VGND VPWR VPWR _31779_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33517_ _34093_/CLK _33517_/D VGND VGND VPWR VPWR _33517_/Q sky130_fd_sc_hd__dfxtp_1
X_21531_ _21526_/X _21530_/X _21387_/X _21388_/X VGND VGND VPWR VPWR _21548_/B sky130_fd_sc_hd__o211a_1
XFILLER_107_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30729_ _30729_/A VGND VGND VPWR VPWR _35599_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34497_ _34626_/CLK _34497_/D VGND VGND VPWR VPWR _34497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36236_ _36242_/CLK _36236_/D VGND VGND VPWR VPWR _36236_/Q sky130_fd_sc_hd__dfxtp_1
X_24250_ _24250_/A VGND VGND VPWR VPWR _32660_/D sky130_fd_sc_hd__clkbuf_1
X_21462_ _32108_/Q _32300_/Q _32364_/Q _35884_/Q _21174_/X _21315_/X VGND VGND VPWR
+ VPWR _21462_/X sky130_fd_sc_hd__mux4_1
X_33448_ _35622_/CLK _33448_/D VGND VGND VPWR VPWR _33448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20413_ _35728_/Q _32239_/Q _35600_/Q _35536_/Q _18293_/X _18295_/X VGND VGND VPWR
+ VPWR _20413_/X sky130_fd_sc_hd__mux4_1
X_23201_ _23049_/X _32138_/Q _23215_/S VGND VGND VPWR VPWR _23202_/A sky130_fd_sc_hd__mux2_1
X_36167_ _36167_/CLK _36167_/D VGND VGND VPWR VPWR _36167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33379_ _33828_/CLK _33379_/D VGND VGND VPWR VPWR _33379_/Q sky130_fd_sc_hd__dfxtp_1
X_21393_ _35626_/Q _34986_/Q _34346_/Q _33706_/Q _21391_/X _21392_/X VGND VGND VPWR
+ VPWR _21393_/X sky130_fd_sc_hd__mux4_1
X_24181_ _24181_/A VGND VGND VPWR VPWR _32627_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20344_ _20212_/X _20342_/X _20343_/X _20215_/X VGND VGND VPWR VPWR _20344_/X sky130_fd_sc_hd__a22o_1
X_35118_ _36142_/CLK _35118_/D VGND VGND VPWR VPWR _35118_/Q sky130_fd_sc_hd__dfxtp_1
X_23132_ _23132_/A VGND VGND VPWR VPWR _32105_/D sky130_fd_sc_hd__clkbuf_1
X_36098_ _36099_/CLK _36098_/D VGND VGND VPWR VPWR _36098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1078 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27940_ _27788_/X _34309_/Q _27944_/S VGND VGND VPWR VPWR _27941_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23063_ _23063_/A VGND VGND VPWR VPWR _32078_/D sky130_fd_sc_hd__clkbuf_1
X_20275_ _33676_/Q _33612_/Q _33548_/Q _33484_/Q _20206_/X _20207_/X VGND VGND VPWR
+ VPWR _20275_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_304_CLK clkbuf_6_51__f_CLK/X VGND VGND VPWR VPWR _35845_/CLK sky130_fd_sc_hd__clkbuf_16
X_35049_ _36137_/CLK _35049_/D VGND VGND VPWR VPWR _35049_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22014_ _32636_/Q _32572_/Q _32508_/Q _35964_/Q _21876_/X _22013_/X VGND VGND VPWR
+ VPWR _22014_/X sky130_fd_sc_hd__mux4_1
XTAP_6139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27871_ _27686_/X _34276_/Q _27881_/S VGND VGND VPWR VPWR _27872_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26822_ _26822_/A VGND VGND VPWR VPWR _33841_/D sky130_fd_sc_hd__clkbuf_1
X_29610_ _35069_/Q _29450_/X _29610_/S VGND VGND VPWR VPWR _29611_/A sky130_fd_sc_hd__mux2_1
XTAP_5449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29541_ _35036_/Q _29348_/X _29547_/S VGND VGND VPWR VPWR _29542_/A sky130_fd_sc_hd__mux2_1
XTAP_4737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26753_ _33809_/Q _23484_/X _26753_/S VGND VGND VPWR VPWR _26754_/A sky130_fd_sc_hd__mux2_1
XTAP_4748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23965_ _23064_/X _32527_/Q _23969_/S VGND VGND VPWR VPWR _23966_/A sky130_fd_sc_hd__mux2_1
X_25704_ _24837_/X _33314_/Q _25718_/S VGND VGND VPWR VPWR _25705_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29472_ input41/X VGND VGND VPWR VPWR _29472_/X sky130_fd_sc_hd__buf_2
X_22916_ _22915_/X _32031_/Q _22916_/S VGND VGND VPWR VPWR _22917_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26684_ _33776_/Q _23340_/X _26690_/S VGND VGND VPWR VPWR _26685_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23896_ _22962_/X _32494_/Q _23906_/S VGND VGND VPWR VPWR _23897_/A sky130_fd_sc_hd__mux2_1
X_28423_ _28513_/S VGND VGND VPWR VPWR _28442_/S sky130_fd_sc_hd__buf_4
X_25635_ _25635_/A VGND VGND VPWR VPWR _33281_/D sky130_fd_sc_hd__clkbuf_1
X_22847_ _22847_/A _22847_/B _22847_/C _22847_/D VGND VGND VPWR VPWR _22848_/A sky130_fd_sc_hd__or4_4
XFILLER_204_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_1188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28354_ _27801_/X _34505_/Q _28370_/S VGND VGND VPWR VPWR _28355_/A sky130_fd_sc_hd__mux2_1
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25566_ _25566_/A VGND VGND VPWR VPWR _33248_/D sky130_fd_sc_hd__clkbuf_1
X_22778_ _20601_/X _22776_/X _22777_/X _20607_/X VGND VGND VPWR VPWR _22778_/X sky130_fd_sc_hd__a22o_1
XFILLER_231_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27305_ _34039_/Q _27137_/X _27317_/S VGND VGND VPWR VPWR _27306_/A sky130_fd_sc_hd__mux2_1
XFILLER_212_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24517_ _24517_/A VGND VGND VPWR VPWR _32785_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21729_ _33396_/Q _33332_/Q _33268_/Q _33204_/Q _21727_/X _21728_/X VGND VGND VPWR
+ VPWR _21729_/X sky130_fd_sc_hd__mux4_1
X_28285_ _28285_/A VGND VGND VPWR VPWR _34472_/D sky130_fd_sc_hd__clkbuf_1
X_25497_ _24930_/X _33216_/Q _25511_/S VGND VGND VPWR VPWR _25498_/A sky130_fd_sc_hd__mux2_1
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27236_ _34006_/Q _27033_/X _27254_/S VGND VGND VPWR VPWR _27237_/A sky130_fd_sc_hd__mux2_1
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24448_ _24448_/A VGND VGND VPWR VPWR _32752_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27167_ _27167_/A VGND VGND VPWR VPWR _33984_/D sky130_fd_sc_hd__clkbuf_1
X_24379_ _23067_/X _32720_/Q _24381_/S VGND VGND VPWR VPWR _24380_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26118_ _26118_/A VGND VGND VPWR VPWR _33510_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27098_ _33962_/Q _27096_/X _27125_/S VGND VGND VPWR VPWR _27099_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26049_ _24948_/X _33478_/Q _26051_/S VGND VGND VPWR VPWR _26050_/A sky130_fd_sc_hd__mux2_1
X_18940_ _20133_/A VGND VGND VPWR VPWR _18940_/X sky130_fd_sc_hd__buf_4
XFILLER_165_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18871_ _32612_/Q _32548_/Q _32484_/Q _35940_/Q _18870_/X _18654_/X VGND VGND VPWR
+ VPWR _18871_/X sky130_fd_sc_hd__mux4_1
XTAP_6640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29808_ _29808_/A VGND VGND VPWR VPWR _35162_/D sky130_fd_sc_hd__clkbuf_1
X_17822_ _35207_/Q _35143_/Q _35079_/Q _32263_/Q _17716_/X _17717_/X VGND VGND VPWR
+ VPWR _17822_/X sky130_fd_sc_hd__mux4_1
XTAP_6684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17753_ _34949_/Q _34885_/Q _34821_/Q _34757_/Q _17513_/X _17514_/X VGND VGND VPWR
+ VPWR _17753_/X sky130_fd_sc_hd__mux4_1
XTAP_5983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29739_ _35130_/Q _29441_/X _29745_/S VGND VGND VPWR VPWR _29740_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16704_ _16500_/X _16702_/X _16703_/X _16503_/X VGND VGND VPWR VPWR _16704_/X sky130_fd_sc_hd__a22o_1
X_17684_ _17511_/X _17682_/X _17683_/X _17516_/X VGND VGND VPWR VPWR _17684_/X sky130_fd_sc_hd__a22o_1
X_32750_ _32877_/CLK _32750_/D VGND VGND VPWR VPWR _32750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31701_ _31701_/A VGND VGND VPWR VPWR _36059_/D sky130_fd_sc_hd__clkbuf_1
X_16635_ _16631_/X _16634_/X _16426_/X VGND VGND VPWR VPWR _16665_/A sky130_fd_sc_hd__o21ba_1
X_19423_ _19423_/A VGND VGND VPWR VPWR _32435_/D sky130_fd_sc_hd__clkbuf_1
X_32681_ _32808_/CLK _32681_/D VGND VGND VPWR VPWR _32681_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_245_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34420_ _36149_/CLK _34420_/D VGND VGND VPWR VPWR _34420_/Q sky130_fd_sc_hd__dfxtp_1
X_31632_ _27757_/X _36027_/Q _31636_/S VGND VGND VPWR VPWR _31633_/A sky130_fd_sc_hd__mux2_1
XFILLER_206_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19354_ _19146_/X _19352_/X _19353_/X _19151_/X VGND VGND VPWR VPWR _19354_/X sky130_fd_sc_hd__a22o_1
X_16566_ _33380_/Q _33316_/Q _33252_/Q _33188_/Q _16421_/X _16422_/X VGND VGND VPWR
+ VPWR _16566_/X sky130_fd_sc_hd__mux4_1
XFILLER_245_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18305_ input80/X input79/X VGND VGND VPWR VPWR _20077_/A sky130_fd_sc_hd__nor2b_4
XFILLER_15_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31563_ _27655_/X _35994_/Q _31573_/S VGND VGND VPWR VPWR _31564_/A sky130_fd_sc_hd__mux2_1
X_19285_ _33392_/Q _33328_/Q _33264_/Q _33200_/Q _19074_/X _19075_/X VGND VGND VPWR
+ VPWR _19285_/X sky130_fd_sc_hd__mux4_1
X_34351_ _35630_/CLK _34351_/D VGND VGND VPWR VPWR _34351_/Q sky130_fd_sc_hd__dfxtp_1
X_16497_ _34146_/Q _34082_/Q _34018_/Q _33954_/Q _16387_/X _16388_/X VGND VGND VPWR
+ VPWR _16497_/X sky130_fd_sc_hd__mux4_1
XFILLER_200_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18236_ _35476_/Q _35412_/Q _35348_/Q _35284_/Q _17960_/X _17961_/X VGND VGND VPWR
+ VPWR _18236_/X sky130_fd_sc_hd__mux4_1
X_33302_ _35804_/CLK _33302_/D VGND VGND VPWR VPWR _33302_/Q sky130_fd_sc_hd__dfxtp_1
X_30514_ _30514_/A VGND VGND VPWR VPWR _35497_/D sky130_fd_sc_hd__clkbuf_1
X_34282_ _36140_/CLK _34282_/D VGND VGND VPWR VPWR _34282_/Q sky130_fd_sc_hd__dfxtp_1
X_31494_ _31494_/A VGND VGND VPWR VPWR _35961_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33233_ _36106_/CLK _33233_/D VGND VGND VPWR VPWR _33233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36021_ _36021_/CLK _36021_/D VGND VGND VPWR VPWR _36021_/Q sky130_fd_sc_hd__dfxtp_1
X_30445_ _30445_/A VGND VGND VPWR VPWR _35464_/D sky130_fd_sc_hd__clkbuf_1
X_18167_ _33170_/Q _36050_/Q _33042_/Q _32978_/Q _16032_/X _17161_/A VGND VGND VPWR
+ VPWR _18167_/X sky130_fd_sc_hd__mux4_1
XFILLER_15_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_90_CLK clkbuf_leaf_96_CLK/A VGND VGND VPWR VPWR _35615_/CLK sky130_fd_sc_hd__clkbuf_16
X_17118_ _34419_/Q _36147_/Q _34291_/Q _34227_/Q _16876_/X _16877_/X VGND VGND VPWR
+ VPWR _17118_/X sky130_fd_sc_hd__mux4_1
XFILLER_209_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33164_ _36044_/CLK _33164_/D VGND VGND VPWR VPWR _33164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18098_ _18098_/A VGND VGND VPWR VPWR _32015_/D sky130_fd_sc_hd__buf_2
X_30376_ _35432_/Q _29385_/X _30378_/S VGND VGND VPWR VPWR _30377_/A sky130_fd_sc_hd__mux2_1
XFILLER_209_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32115_ _32882_/CLK _32115_/D VGND VGND VPWR VPWR _32115_/Q sky130_fd_sc_hd__dfxtp_1
X_17049_ _17045_/X _17048_/X _16812_/X VGND VGND VPWR VPWR _17050_/D sky130_fd_sc_hd__o21ba_1
X_33095_ _35845_/CLK _33095_/D VGND VGND VPWR VPWR _33095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20060_ _19852_/X _20058_/X _20059_/X _19857_/X VGND VGND VPWR VPWR _20060_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32046_ _36015_/CLK _32046_/D VGND VGND VPWR VPWR _32046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_1070 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35805_ _35805_/CLK _35805_/D VGND VGND VPWR VPWR _35805_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33997_ _34193_/CLK _33997_/D VGND VGND VPWR VPWR _33997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35736_ _35800_/CLK _35736_/D VGND VGND VPWR VPWR _35736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23750_ _23840_/S VGND VGND VPWR VPWR _23769_/S sky130_fd_sc_hd__buf_4
XFILLER_226_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20962_ _22374_/A VGND VGND VPWR VPWR _20962_/X sky130_fd_sc_hd__buf_4
X_32948_ _36020_/CLK _32948_/D VGND VGND VPWR VPWR _32948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22701_ _22505_/X _22699_/X _22700_/X _22510_/X VGND VGND VPWR VPWR _22701_/X sky130_fd_sc_hd__a22o_1
XFILLER_241_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35667_ _35729_/CLK _35667_/D VGND VGND VPWR VPWR _35667_/Q sky130_fd_sc_hd__dfxtp_1
X_23681_ _23681_/A VGND VGND VPWR VPWR _32330_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20893_ _35676_/Q _32182_/Q _35548_/Q _35484_/Q _20858_/X _20859_/X VGND VGND VPWR
+ VPWR _20893_/X sky130_fd_sc_hd__mux4_1
X_32879_ _32879_/CLK _32879_/D VGND VGND VPWR VPWR _32879_/Q sky130_fd_sc_hd__dfxtp_1
X_25420_ _25420_/A VGND VGND VPWR VPWR _33179_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_242_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22632_ _22459_/X _22630_/X _22631_/X _22462_/X VGND VGND VPWR VPWR _22632_/X sky130_fd_sc_hd__a22o_1
X_34618_ _35835_/CLK _34618_/D VGND VGND VPWR VPWR _34618_/Q sky130_fd_sc_hd__dfxtp_1
X_35598_ _35599_/CLK _35598_/D VGND VGND VPWR VPWR _35598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1044 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25351_ _33148_/Q _23414_/X _25353_/S VGND VGND VPWR VPWR _25352_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22563_ _33099_/Q _32075_/Q _35851_/Q _35787_/Q _22384_/X _22385_/X VGND VGND VPWR
+ VPWR _22563_/X sky130_fd_sc_hd__mux4_1
X_34549_ _36149_/CLK _34549_/D VGND VGND VPWR VPWR _34549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24302_ _22953_/X _32683_/Q _24318_/S VGND VGND VPWR VPWR _24303_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28070_ _28070_/A VGND VGND VPWR VPWR _34370_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21514_ _21514_/A _21514_/B _21514_/C _21514_/D VGND VGND VPWR VPWR _21515_/A sky130_fd_sc_hd__or4_4
XFILLER_210_876 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25282_ _33115_/Q _23246_/X _25290_/S VGND VGND VPWR VPWR _25283_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22494_ _22309_/X _22492_/X _22493_/X _22312_/X VGND VGND VPWR VPWR _22494_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_908 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27021_ _33936_/Q _23481_/X _27023_/S VGND VGND VPWR VPWR _27022_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_898 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36219_ _36219_/CLK _36219_/D VGND VGND VPWR VPWR _36219_/Q sky130_fd_sc_hd__dfxtp_1
X_24233_ _32652_/Q _23469_/X _24243_/S VGND VGND VPWR VPWR _24234_/A sky130_fd_sc_hd__mux2_1
X_21445_ _21445_/A VGND VGND VPWR VPWR _36203_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_81_CLK clkbuf_leaf_81_CLK/A VGND VGND VPWR VPWR _35804_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_68_1416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21376_ _33386_/Q _33322_/Q _33258_/Q _33194_/Q _21374_/X _21375_/X VGND VGND VPWR
+ VPWR _21376_/X sky130_fd_sc_hd__mux4_1
X_24164_ _32619_/Q _23296_/X _24180_/S VGND VGND VPWR VPWR _24165_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20327_ _33101_/Q _32077_/Q _35853_/Q _35789_/Q _20084_/X _20085_/X VGND VGND VPWR
+ VPWR _20327_/X sky130_fd_sc_hd__mux4_1
X_23115_ _22922_/X _32097_/Q _23131_/S VGND VGND VPWR VPWR _23116_/A sky130_fd_sc_hd__mux2_1
XFILLER_235_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24095_ _23055_/X _32588_/Q _24105_/S VGND VGND VPWR VPWR _24096_/A sky130_fd_sc_hd__mux2_1
X_28972_ _28972_/A VGND VGND VPWR VPWR _34796_/D sky130_fd_sc_hd__clkbuf_1
X_20258_ _35659_/Q _35019_/Q _34379_/Q _33739_/Q _20150_/X _20151_/X VGND VGND VPWR
+ VPWR _20258_/X sky130_fd_sc_hd__mux4_1
XFILLER_122_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23046_ input47/X VGND VGND VPWR VPWR _23046_/X sky130_fd_sc_hd__buf_2
X_27923_ _27763_/X _34301_/Q _27923_/S VGND VGND VPWR VPWR _27924_/A sky130_fd_sc_hd__mux2_1
XTAP_5202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27854_ _27661_/X _34268_/Q _27860_/S VGND VGND VPWR VPWR _27855_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20189_ _35721_/Q _32232_/Q _35593_/Q _35529_/Q _19970_/X _19971_/X VGND VGND VPWR
+ VPWR _20189_/X sky130_fd_sc_hd__mux4_1
XTAP_5235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26805_ _26805_/A VGND VGND VPWR VPWR _33833_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27785_ input41/X VGND VGND VPWR VPWR _27785_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24997_ _28380_/A _31553_/B VGND VGND VPWR VPWR _25130_/S sky130_fd_sc_hd__nand2_8
XTAP_4556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26736_ _26736_/A VGND VGND VPWR VPWR _33800_/D sky130_fd_sc_hd__clkbuf_1
X_29524_ input60/X VGND VGND VPWR VPWR _29524_/X sky130_fd_sc_hd__clkbuf_4
XTAP_4578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23948_ _23039_/X _32519_/Q _23948_/S VGND VGND VPWR VPWR _23949_/A sky130_fd_sc_hd__mux2_1
XTAP_3844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29455_ _35006_/Q _29453_/X _29482_/S VGND VGND VPWR VPWR _29456_/A sky130_fd_sc_hd__mux2_1
XTAP_3877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26667_ _33768_/Q _23286_/X _26669_/S VGND VGND VPWR VPWR _26668_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_867 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23879_ _22937_/X _32486_/Q _23885_/S VGND VGND VPWR VPWR _23880_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16420_ _16140_/X _16418_/X _16419_/X _16145_/X VGND VGND VPWR VPWR _16420_/X sky130_fd_sc_hd__a22o_1
X_25618_ _25618_/A VGND VGND VPWR VPWR _33273_/D sky130_fd_sc_hd__clkbuf_1
X_28406_ _28406_/A VGND VGND VPWR VPWR _34529_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29386_ _34984_/Q _29385_/X _29389_/S VGND VGND VPWR VPWR _29387_/A sky130_fd_sc_hd__mux2_1
X_26598_ _24958_/X _33737_/Q _26614_/S VGND VGND VPWR VPWR _26599_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28337_ _27776_/X _34497_/Q _28349_/S VGND VGND VPWR VPWR _28338_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16351_ _16147_/X _16349_/X _16350_/X _16150_/X VGND VGND VPWR VPWR _16351_/X sky130_fd_sc_hd__a22o_1
X_25549_ _25549_/A VGND VGND VPWR VPWR _33240_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19070_ _19070_/A VGND VGND VPWR VPWR _32425_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_185_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16282_ _16278_/X _16281_/X _16015_/X VGND VGND VPWR VPWR _16312_/A sky130_fd_sc_hd__o21ba_1
X_28268_ _27673_/X _34464_/Q _28286_/S VGND VGND VPWR VPWR _28269_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18021_ _17773_/X _18019_/X _18020_/X _17777_/X VGND VGND VPWR VPWR _18021_/X sky130_fd_sc_hd__a22o_1
X_27219_ _27219_/A VGND VGND VPWR VPWR _34001_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28199_ _28199_/A VGND VGND VPWR VPWR _34431_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_72_CLK clkbuf_leaf_73_CLK/A VGND VGND VPWR VPWR _32797_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30230_ _30230_/A VGND VGND VPWR VPWR _35362_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_1_0_CLK clkbuf_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_9_0_CLK/A sky130_fd_sc_hd__clkbuf_8
XFILLER_5_974 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30161_ _35330_/Q _29466_/X _30171_/S VGND VGND VPWR VPWR _30162_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19972_ _35715_/Q _32225_/Q _35587_/Q _35523_/Q _19970_/X _19971_/X VGND VGND VPWR
+ VPWR _19972_/X sky130_fd_sc_hd__mux4_1
XFILLER_141_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18923_ _34405_/Q _36133_/Q _34277_/Q _34213_/Q _18823_/X _18824_/X VGND VGND VPWR
+ VPWR _18923_/X sky130_fd_sc_hd__mux4_1
X_30092_ _35297_/Q _29364_/X _30108_/S VGND VGND VPWR VPWR _30093_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33920_ _33921_/CLK _33920_/D VGND VGND VPWR VPWR _33920_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18854_ _34659_/Q _34595_/Q _34531_/Q _34467_/Q _18533_/X _18534_/X VGND VGND VPWR
+ VPWR _18854_/X sky130_fd_sc_hd__mux4_1
XTAP_6470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17805_ _17559_/X _17803_/X _17804_/X _17562_/X VGND VGND VPWR VPWR _17805_/X sky130_fd_sc_hd__a22o_1
XFILLER_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33851_ _36092_/CLK _33851_/D VGND VGND VPWR VPWR _33851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15997_ _15981_/X _15988_/X _15991_/X _15996_/X VGND VGND VPWR VPWR _15997_/X sky130_fd_sc_hd__a22o_1
X_18785_ _35169_/Q _35105_/Q _35041_/Q _32161_/Q _18604_/X _18605_/X VGND VGND VPWR
+ VPWR _18785_/X sky130_fd_sc_hd__mux4_1
XFILLER_95_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32802_ _32802_/CLK _32802_/D VGND VGND VPWR VPWR _32802_/Q sky130_fd_sc_hd__dfxtp_1
X_17736_ _33157_/Q _36037_/Q _33029_/Q _32965_/Q _17415_/X _17416_/X VGND VGND VPWR
+ VPWR _17736_/X sky130_fd_sc_hd__mux4_1
X_30994_ _35725_/Q input51/X _31002_/S VGND VGND VPWR VPWR _30995_/A sky130_fd_sc_hd__mux2_1
X_33782_ _33910_/CLK _33782_/D VGND VGND VPWR VPWR _33782_/Q sky130_fd_sc_hd__dfxtp_1
X_35521_ _35646_/CLK _35521_/D VGND VGND VPWR VPWR _35521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32733_ _32797_/CLK _32733_/D VGND VGND VPWR VPWR _32733_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17667_ _32899_/Q _32835_/Q _32771_/Q _32707_/Q _17346_/X _17347_/X VGND VGND VPWR
+ VPWR _17667_/X sky130_fd_sc_hd__mux4_1
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19406_ _19367_/X _19404_/X _19405_/X _19371_/X VGND VGND VPWR VPWR _19406_/X sky130_fd_sc_hd__a22o_1
X_16618_ _16297_/X _16616_/X _16617_/X _16300_/X VGND VGND VPWR VPWR _16618_/X sky130_fd_sc_hd__a22o_1
X_35452_ _35708_/CLK _35452_/D VGND VGND VPWR VPWR _35452_/Q sky130_fd_sc_hd__dfxtp_1
X_32664_ _36119_/CLK _32664_/D VGND VGND VPWR VPWR _32664_/Q sky130_fd_sc_hd__dfxtp_1
X_17598_ _33153_/Q _36033_/Q _33025_/Q _32961_/Q _17415_/X _17416_/X VGND VGND VPWR
+ VPWR _17598_/X sky130_fd_sc_hd__mux4_1
XFILLER_50_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34403_ _34405_/CLK _34403_/D VGND VGND VPWR VPWR _34403_/Q sky130_fd_sc_hd__dfxtp_1
X_19337_ _35633_/Q _34993_/Q _34353_/Q _33713_/Q _19091_/X _19092_/X VGND VGND VPWR
+ VPWR _19337_/X sky130_fd_sc_hd__mux4_1
X_16549_ _17961_/A VGND VGND VPWR VPWR _16549_/X sky130_fd_sc_hd__clkbuf_4
X_31615_ _27732_/X _36019_/Q _31615_/S VGND VGND VPWR VPWR _31616_/A sky130_fd_sc_hd__mux2_1
X_35383_ _35769_/CLK _35383_/D VGND VGND VPWR VPWR _35383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32595_ _36049_/CLK _32595_/D VGND VGND VPWR VPWR _32595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34334_ _35615_/CLK _34334_/D VGND VGND VPWR VPWR _34334_/Q sky130_fd_sc_hd__dfxtp_1
X_31546_ _31546_/A VGND VGND VPWR VPWR _35986_/D sky130_fd_sc_hd__clkbuf_1
X_19268_ _18945_/X _19266_/X _19267_/X _18948_/X VGND VGND VPWR VPWR _19268_/X sky130_fd_sc_hd__a22o_1
X_18219_ _33684_/Q _33620_/Q _33556_/Q _33492_/Q _16024_/X _16025_/X VGND VGND VPWR
+ VPWR _18219_/X sky130_fd_sc_hd__mux4_1
X_34265_ _36121_/CLK _34265_/D VGND VGND VPWR VPWR _34265_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_507_CLK clkbuf_leaf_2_CLK/A VGND VGND VPWR VPWR _34151_/CLK sky130_fd_sc_hd__clkbuf_16
X_19199_ _35629_/Q _34989_/Q _34349_/Q _33709_/Q _19091_/X _19092_/X VGND VGND VPWR
+ VPWR _19199_/X sky130_fd_sc_hd__mux4_1
X_31477_ _31477_/A VGND VGND VPWR VPWR _35953_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_63_CLK clkbuf_leaf_65_CLK/A VGND VGND VPWR VPWR _35985_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_102_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21230_ _34150_/Q _34086_/Q _34022_/Q _33958_/Q _20987_/X _20988_/X VGND VGND VPWR
+ VPWR _21230_/X sky130_fd_sc_hd__mux4_1
X_36004_ _36005_/CLK _36004_/D VGND VGND VPWR VPWR _36004_/Q sky130_fd_sc_hd__dfxtp_1
X_33216_ _33921_/CLK _33216_/D VGND VGND VPWR VPWR _33216_/Q sky130_fd_sc_hd__dfxtp_1
X_30428_ _30428_/A VGND VGND VPWR VPWR _35456_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34196_ _34773_/CLK _34196_/D VGND VGND VPWR VPWR _34196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21161_ _21161_/A _21161_/B _21161_/C _21161_/D VGND VGND VPWR VPWR _21162_/A sky130_fd_sc_hd__or4_1
XFILLER_137_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30359_ _30470_/S VGND VGND VPWR VPWR _30378_/S sky130_fd_sc_hd__buf_4
X_33147_ _35835_/CLK _33147_/D VGND VGND VPWR VPWR _33147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20112_ _20073_/X _20110_/X _20111_/X _20077_/X VGND VGND VPWR VPWR _20112_/X sky130_fd_sc_hd__a22o_1
X_21092_ _21092_/A VGND VGND VPWR VPWR _36193_/D sky130_fd_sc_hd__clkbuf_1
X_33078_ _35830_/CLK _33078_/D VGND VGND VPWR VPWR _33078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20043_ _35653_/Q _35013_/Q _34373_/Q _33733_/Q _19797_/X _19798_/X VGND VGND VPWR
+ VPWR _20043_/X sky130_fd_sc_hd__mux4_1
X_32029_ _35998_/CLK _32029_/D VGND VGND VPWR VPWR _32029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24920_ input33/X VGND VGND VPWR VPWR _24920_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_112_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24851_ _24851_/A VGND VGND VPWR VPWR _32934_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23802_ _23802_/A VGND VGND VPWR VPWR _32386_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27570_ _27570_/A VGND VGND VPWR VPWR _34164_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_227_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24782_ _23064_/X _32911_/Q _24786_/S VGND VGND VPWR VPWR _24783_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21994_ _21956_/X _21992_/X _21993_/X _21959_/X VGND VGND VPWR VPWR _21994_/X sky130_fd_sc_hd__a22o_1
XFILLER_38_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26521_ _26521_/A VGND VGND VPWR VPWR _33700_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35719_ _35721_/CLK _35719_/D VGND VGND VPWR VPWR _35719_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23733_ _23733_/A VGND VGND VPWR VPWR _32353_/D sky130_fd_sc_hd__clkbuf_1
X_20945_ _20945_/A VGND VGND VPWR VPWR _36189_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29240_ _29240_/A VGND VGND VPWR VPWR _34923_/D sky130_fd_sc_hd__clkbuf_1
X_26452_ _26452_/A VGND VGND VPWR VPWR _33668_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23664_ _23664_/A VGND VGND VPWR VPWR _32322_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20876_ _33628_/Q _33564_/Q _33500_/Q _33436_/Q _20741_/X _20742_/X VGND VGND VPWR
+ VPWR _20876_/X sky130_fd_sc_hd__mux4_1
XFILLER_144_1109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25403_ _33173_/Q _23498_/X _25403_/S VGND VGND VPWR VPWR _25404_/A sky130_fd_sc_hd__mux2_1
X_29171_ _34891_/Q _27199_/X _29183_/S VGND VGND VPWR VPWR _29172_/A sky130_fd_sc_hd__mux2_1
X_22615_ _22611_/X _22614_/X _22438_/X VGND VGND VPWR VPWR _22637_/A sky130_fd_sc_hd__o21ba_1
XFILLER_201_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26383_ _26383_/A VGND VGND VPWR VPWR _33635_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23595_ _23595_/A VGND VGND VPWR VPWR _32289_/D sky130_fd_sc_hd__clkbuf_1
X_28122_ _27658_/X _34395_/Q _28130_/S VGND VGND VPWR VPWR _28123_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_6_37__f_CLK clkbuf_5_18_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_37__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_210_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25334_ _25403_/S VGND VGND VPWR VPWR _25353_/S sky130_fd_sc_hd__buf_4
X_22546_ _33419_/Q _33355_/Q _33291_/Q _33227_/Q _22433_/X _22434_/X VGND VGND VPWR
+ VPWR _22546_/X sky130_fd_sc_hd__mux4_1
XFILLER_220_1008 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28053_ _28053_/A VGND VGND VPWR VPWR _34362_/D sky130_fd_sc_hd__clkbuf_1
X_25265_ _33108_/Q _23495_/X _25267_/S VGND VGND VPWR VPWR _25266_/A sky130_fd_sc_hd__mux2_1
X_22477_ _22152_/X _22475_/X _22476_/X _22157_/X VGND VGND VPWR VPWR _22477_/X sky130_fd_sc_hd__a22o_1
XFILLER_120_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_54_CLK clkbuf_leaf_57_CLK/A VGND VGND VPWR VPWR _32804_/CLK sky130_fd_sc_hd__clkbuf_16
X_27004_ _27031_/S VGND VGND VPWR VPWR _27023_/S sky130_fd_sc_hd__buf_4
X_24216_ _32644_/Q _23441_/X _24222_/S VGND VGND VPWR VPWR _24217_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21428_ _21314_/X _21426_/X _21427_/X _21318_/X VGND VGND VPWR VPWR _21428_/X sky130_fd_sc_hd__a22o_1
XFILLER_107_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25196_ _33075_/Q _23384_/X _25196_/S VGND VGND VPWR VPWR _25197_/A sky130_fd_sc_hd__mux2_1
XFILLER_205_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24147_ _32611_/Q _23271_/X _24159_/S VGND VGND VPWR VPWR _24148_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21359_ _33065_/Q _32041_/Q _35817_/Q _35753_/Q _21325_/X _21326_/X VGND VGND VPWR
+ VPWR _21359_/X sky130_fd_sc_hd__mux4_1
XFILLER_190_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24078_ _23030_/X _32580_/Q _24084_/S VGND VGND VPWR VPWR _24079_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28955_ _28955_/A VGND VGND VPWR VPWR _34788_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23029_ _23029_/A VGND VGND VPWR VPWR _32067_/D sky130_fd_sc_hd__clkbuf_1
X_27906_ _27906_/A VGND VGND VPWR VPWR _34292_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28886_ _34756_/Q _27177_/X _28892_/S VGND VGND VPWR VPWR _28887_/A sky130_fd_sc_hd__mux2_1
XTAP_5032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27837_ input60/X VGND VGND VPWR VPWR _27837_/X sky130_fd_sc_hd__clkbuf_4
XTAP_5065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18570_ _34395_/Q _36123_/Q _34267_/Q _34203_/Q _18470_/X _18471_/X VGND VGND VPWR
+ VPWR _18570_/X sky130_fd_sc_hd__mux4_1
X_27768_ _27766_/X _34238_/Q _27795_/S VGND VGND VPWR VPWR _27769_/A sky130_fd_sc_hd__mux2_1
XTAP_4375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29507_ _35023_/Q _29506_/X _29513_/S VGND VGND VPWR VPWR _29508_/A sky130_fd_sc_hd__mux2_1
X_17521_ _17521_/A VGND VGND VPWR VPWR _31998_/D sky130_fd_sc_hd__buf_4
XTAP_3663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26719_ _26719_/A VGND VGND VPWR VPWR _33792_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27699_ _27698_/X _34216_/Q _27702_/S VGND VGND VPWR VPWR _27700_/A sky130_fd_sc_hd__mux2_1
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17452_ _17206_/X _17450_/X _17451_/X _17209_/X VGND VGND VPWR VPWR _17452_/X sky130_fd_sc_hd__a22o_1
XTAP_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29438_ input29/X VGND VGND VPWR VPWR _29438_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16403_ _35615_/Q _34975_/Q _34335_/Q _33695_/Q _16053_/X _16055_/X VGND VGND VPWR
+ VPWR _16403_/X sky130_fd_sc_hd__mux4_1
XFILLER_177_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17383_ _33147_/Q _36027_/Q _33019_/Q _32955_/Q _17062_/X _17063_/X VGND VGND VPWR
+ VPWR _17383_/X sky130_fd_sc_hd__mux4_1
X_29369_ _29369_/A VGND VGND VPWR VPWR _34978_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16334_ _33053_/Q _32029_/Q _35805_/Q _35741_/Q _16067_/X _16069_/X VGND VGND VPWR
+ VPWR _16334_/X sky130_fd_sc_hd__mux4_1
X_31400_ _27813_/X _35917_/Q _31408_/S VGND VGND VPWR VPWR _31401_/A sky130_fd_sc_hd__mux2_1
X_19122_ _19118_/X _19121_/X _19079_/X VGND VGND VPWR VPWR _19144_/A sky130_fd_sc_hd__o21ba_1
X_32380_ _35964_/CLK _32380_/D VGND VGND VPWR VPWR _32380_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31331_ _27711_/X _35884_/Q _31345_/S VGND VGND VPWR VPWR _31332_/A sky130_fd_sc_hd__mux2_1
X_19053_ _19014_/X _19051_/X _19052_/X _19018_/X VGND VGND VPWR VPWR _19053_/X sky130_fd_sc_hd__a22o_1
X_16265_ _16060_/X _16263_/X _16264_/X _16072_/X VGND VGND VPWR VPWR _16265_/X sky130_fd_sc_hd__a22o_1
XFILLER_16_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_1250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_45_CLK clkbuf_6_6__f_CLK/X VGND VGND VPWR VPWR _35814_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_195_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18004_ _34956_/Q _34892_/Q _34828_/Q _34764_/Q _17866_/X _17867_/X VGND VGND VPWR
+ VPWR _18004_/X sky130_fd_sc_hd__mux4_1
X_34050_ _34945_/CLK _34050_/D VGND VGND VPWR VPWR _34050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31262_ _31262_/A VGND VGND VPWR VPWR _35851_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16196_ _17851_/A VGND VGND VPWR VPWR _16196_/X sky130_fd_sc_hd__buf_4
X_30213_ _30213_/A VGND VGND VPWR VPWR _35354_/D sky130_fd_sc_hd__clkbuf_1
X_33001_ _35755_/CLK _33001_/D VGND VGND VPWR VPWR _33001_/Q sky130_fd_sc_hd__dfxtp_1
X_31193_ _31193_/A VGND VGND VPWR VPWR _35818_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30144_ _35322_/Q _29441_/X _30150_/S VGND VGND VPWR VPWR _30145_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19955_ _19955_/A VGND VGND VPWR VPWR _32450_/D sky130_fd_sc_hd__buf_2
XFILLER_68_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18906_ _18653_/X _18904_/X _18905_/X _18659_/X VGND VGND VPWR VPWR _18906_/X sky130_fd_sc_hd__a22o_1
X_34952_ _34954_/CLK _34952_/D VGND VGND VPWR VPWR _34952_/Q sky130_fd_sc_hd__dfxtp_1
X_30075_ _35289_/Q _29339_/X _30087_/S VGND VGND VPWR VPWR _30076_/A sky130_fd_sc_hd__mux2_1
X_19886_ _19811_/X _19884_/X _19885_/X _19816_/X VGND VGND VPWR VPWR _19886_/X sky130_fd_sc_hd__a22o_1
XFILLER_45_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33903_ _36080_/CLK _33903_/D VGND VGND VPWR VPWR _33903_/Q sky130_fd_sc_hd__dfxtp_1
X_18837_ _18833_/X _18836_/X _18726_/X VGND VGND VPWR VPWR _18861_/A sky130_fd_sc_hd__o21ba_1
X_34883_ _36105_/CLK _34883_/D VGND VGND VPWR VPWR _34883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33834_ _34091_/CLK _33834_/D VGND VGND VPWR VPWR _33834_/Q sky130_fd_sc_hd__dfxtp_1
X_18768_ _18447_/X _18766_/X _18767_/X _18450_/X VGND VGND VPWR VPWR _18768_/X sky130_fd_sc_hd__a22o_1
XFILLER_215_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17719_ _17506_/X _17715_/X _17718_/X _17509_/X VGND VGND VPWR VPWR _17719_/X sky130_fd_sc_hd__a22o_1
X_33765_ _36070_/CLK _33765_/D VGND VGND VPWR VPWR _33765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30977_ _35717_/Q input42/X _30981_/S VGND VGND VPWR VPWR _30978_/A sky130_fd_sc_hd__mux2_1
X_18699_ _32863_/Q _32799_/Q _32735_/Q _32671_/Q _18587_/X _18588_/X VGND VGND VPWR
+ VPWR _18699_/X sky130_fd_sc_hd__mux4_1
XFILLER_224_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35504_ _35567_/CLK _35504_/D VGND VGND VPWR VPWR _35504_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20730_ _20726_/X _20729_/X _20675_/X VGND VGND VPWR VPWR _20738_/C sky130_fd_sc_hd__o21ba_1
X_32716_ _32879_/CLK _32716_/D VGND VGND VPWR VPWR _32716_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33696_ _35618_/CLK _33696_/D VGND VGND VPWR VPWR _33696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35435_ _35753_/CLK _35435_/D VGND VGND VPWR VPWR _35435_/Q sky130_fd_sc_hd__dfxtp_1
X_20661_ _20661_/A VGND VGND VPWR VPWR _22450_/A sky130_fd_sc_hd__buf_12
X_32647_ _36038_/CLK _32647_/D VGND VGND VPWR VPWR _32647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22400_ _22400_/A VGND VGND VPWR VPWR _22400_/X sky130_fd_sc_hd__buf_4
XFILLER_51_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20592_ _20661_/A VGND VGND VPWR VPWR _22399_/A sky130_fd_sc_hd__buf_12
X_23380_ _23380_/A VGND VGND VPWR VPWR _32205_/D sky130_fd_sc_hd__clkbuf_1
X_35366_ _35367_/CLK _35366_/D VGND VGND VPWR VPWR _35366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32578_ _35970_/CLK _32578_/D VGND VGND VPWR VPWR _32578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34317_ _36176_/CLK _34317_/D VGND VGND VPWR VPWR _34317_/Q sky130_fd_sc_hd__dfxtp_1
X_22331_ _22451_/A VGND VGND VPWR VPWR _22331_/X sky130_fd_sc_hd__buf_4
X_31529_ _27804_/X _35978_/Q _31543_/S VGND VGND VPWR VPWR _31530_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_36_CLK clkbuf_6_7__f_CLK/X VGND VGND VPWR VPWR _36002_/CLK sky130_fd_sc_hd__clkbuf_16
X_35297_ _35297_/CLK _35297_/D VGND VGND VPWR VPWR _35297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25050_ _25050_/A VGND VGND VPWR VPWR _33006_/D sky130_fd_sc_hd__clkbuf_1
X_34248_ _35212_/CLK _34248_/D VGND VGND VPWR VPWR _34248_/Q sky130_fd_sc_hd__dfxtp_1
X_22262_ _22258_/X _22261_/X _22085_/X VGND VGND VPWR VPWR _22286_/A sky130_fd_sc_hd__o21ba_1
XFILLER_191_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24001_ _24001_/A VGND VGND VPWR VPWR _32543_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21213_ _35685_/Q _32192_/Q _35557_/Q _35493_/Q _21211_/X _21212_/X VGND VGND VPWR
+ VPWR _21213_/X sky130_fd_sc_hd__mux4_2
X_22193_ _33409_/Q _33345_/Q _33281_/Q _33217_/Q _22080_/X _22081_/X VGND VGND VPWR
+ VPWR _22193_/X sky130_fd_sc_hd__mux4_1
X_34179_ _34179_/CLK _34179_/D VGND VGND VPWR VPWR _34179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21144_ _21140_/X _21143_/X _21034_/X _21035_/X VGND VGND VPWR VPWR _21161_/B sky130_fd_sc_hd__o211a_1
XFILLER_232_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28740_ _28740_/A VGND VGND VPWR VPWR _34687_/D sky130_fd_sc_hd__clkbuf_1
X_25952_ _25952_/A VGND VGND VPWR VPWR _33431_/D sky130_fd_sc_hd__clkbuf_1
X_21075_ _20961_/X _21073_/X _21074_/X _20965_/X VGND VGND VPWR VPWR _21075_/X sky130_fd_sc_hd__a22o_1
XFILLER_247_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20026_ _33669_/Q _33605_/Q _33541_/Q _33477_/Q _19853_/X _19854_/X VGND VGND VPWR
+ VPWR _20026_/X sky130_fd_sc_hd__mux4_1
X_24903_ _24902_/X _32951_/Q _24921_/S VGND VGND VPWR VPWR _24904_/A sky130_fd_sc_hd__mux2_1
X_28671_ _34655_/Q _27062_/X _28671_/S VGND VGND VPWR VPWR _28672_/A sky130_fd_sc_hd__mux2_1
X_25883_ _24902_/X _33399_/Q _25895_/S VGND VGND VPWR VPWR _25884_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27622_ _27622_/A VGND VGND VPWR VPWR _34189_/D sky130_fd_sc_hd__clkbuf_1
X_24834_ input3/X VGND VGND VPWR VPWR _24834_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_206_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27553_ _27553_/A VGND VGND VPWR VPWR _34156_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_215_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24765_ _23039_/X _32903_/Q _24765_/S VGND VGND VPWR VPWR _24766_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21977_ _22450_/A VGND VGND VPWR VPWR _21977_/X sky130_fd_sc_hd__buf_8
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26504_ _26504_/A VGND VGND VPWR VPWR _33692_/D sky130_fd_sc_hd__clkbuf_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23716_ _23716_/A VGND VGND VPWR VPWR _32345_/D sky130_fd_sc_hd__clkbuf_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27484_ _34124_/Q _27202_/X _27494_/S VGND VGND VPWR VPWR _27485_/A sky130_fd_sc_hd__mux2_1
XFILLER_214_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20928_ _20630_/X _20926_/X _20927_/X _20641_/X VGND VGND VPWR VPWR _20928_/X sky130_fd_sc_hd__a22o_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24696_ _22937_/X _32870_/Q _24702_/S VGND VGND VPWR VPWR _24697_/A sky130_fd_sc_hd__mux2_1
XFILLER_226_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26435_ _26435_/A VGND VGND VPWR VPWR _33660_/D sky130_fd_sc_hd__clkbuf_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29223_ _29223_/A VGND VGND VPWR VPWR _34915_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23647_ _23647_/A VGND VGND VPWR VPWR _32314_/D sky130_fd_sc_hd__clkbuf_1
X_20859_ _22400_/A VGND VGND VPWR VPWR _20859_/X sky130_fd_sc_hd__buf_4
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_870 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29154_ _34883_/Q _27174_/X _29162_/S VGND VGND VPWR VPWR _29155_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26366_ _26366_/A VGND VGND VPWR VPWR _33627_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23578_ _23578_/A VGND VGND VPWR VPWR _32281_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28105_ _28105_/A VGND VGND VPWR VPWR _34387_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25317_ _25317_/A VGND VGND VPWR VPWR _33131_/D sky130_fd_sc_hd__clkbuf_1
X_22529_ _33098_/Q _32074_/Q _35850_/Q _35786_/Q _22384_/X _22385_/X VGND VGND VPWR
+ VPWR _22529_/X sky130_fd_sc_hd__mux4_1
X_29085_ _34850_/Q _27072_/X _29099_/S VGND VGND VPWR VPWR _29086_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26297_ _26297_/A VGND VGND VPWR VPWR _33595_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_27_CLK clkbuf_6_5__f_CLK/X VGND VGND VPWR VPWR _34594_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_183_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16050_ _17800_/A VGND VGND VPWR VPWR _16050_/X sky130_fd_sc_hd__buf_6
X_28036_ _28036_/A VGND VGND VPWR VPWR _34354_/D sky130_fd_sc_hd__clkbuf_1
X_25248_ _25248_/A VGND VGND VPWR VPWR _33099_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25179_ _25179_/A VGND VGND VPWR VPWR _33066_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1062 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29987_ _29987_/A VGND VGND VPWR VPWR _35247_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19740_ _34940_/Q _34876_/Q _34812_/Q _34748_/Q _19460_/X _19461_/X VGND VGND VPWR
+ VPWR _19740_/X sky130_fd_sc_hd__mux4_1
X_28938_ _28938_/A VGND VGND VPWR VPWR _34780_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16952_ _16846_/X _16950_/X _16951_/X _16851_/X VGND VGND VPWR VPWR _16952_/X sky130_fd_sc_hd__a22o_1
XFILLER_238_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19671_ _19671_/A _19671_/B _19671_/C _19671_/D VGND VGND VPWR VPWR _19672_/A sky130_fd_sc_hd__or4_2
X_16883_ _16883_/A VGND VGND VPWR VPWR _31980_/D sky130_fd_sc_hd__clkbuf_1
X_28869_ _34748_/Q _27152_/X _28871_/S VGND VGND VPWR VPWR _28870_/A sky130_fd_sc_hd__mux2_1
X_18622_ _18616_/X _18621_/X _18315_/X VGND VGND VPWR VPWR _18644_/A sky130_fd_sc_hd__o21ba_1
X_30900_ _35680_/Q input2/X _30918_/S VGND VGND VPWR VPWR _30901_/A sky130_fd_sc_hd__mux2_1
XTAP_4150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31880_ _31880_/A VGND VGND VPWR VPWR _36144_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18553_ _18318_/X _18551_/X _18552_/X _18327_/X VGND VGND VPWR VPWR _18553_/X sky130_fd_sc_hd__a22o_1
X_30831_ _30831_/A VGND VGND VPWR VPWR _35647_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17504_ _17857_/A VGND VGND VPWR VPWR _17504_/X sky130_fd_sc_hd__buf_4
XTAP_3493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33550_ _34064_/CLK _33550_/D VGND VGND VPWR VPWR _33550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18484_ _18480_/X _18483_/X _18315_/X VGND VGND VPWR VPWR _18508_/A sky130_fd_sc_hd__o21ba_1
X_30762_ _35615_/Q input64/X _30762_/S VGND VGND VPWR VPWR _30763_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1036 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32501_ _35956_/CLK _32501_/D VGND VGND VPWR VPWR _32501_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17435_ _17429_/X _17434_/X _17151_/X VGND VGND VPWR VPWR _17443_/C sky130_fd_sc_hd__o21ba_1
X_33481_ _34121_/CLK _33481_/D VGND VGND VPWR VPWR _33481_/Q sky130_fd_sc_hd__dfxtp_1
X_30693_ _35582_/Q _29453_/X _30711_/S VGND VGND VPWR VPWR _30694_/A sky130_fd_sc_hd__mux2_1
X_35220_ _35221_/CLK _35220_/D VGND VGND VPWR VPWR _35220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32432_ _36075_/CLK _32432_/D VGND VGND VPWR VPWR _32432_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17366_ _17153_/X _17362_/X _17365_/X _17156_/X VGND VGND VPWR VPWR _17366_/X sky130_fd_sc_hd__a22o_1
XFILLER_18_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_20__f_CLK clkbuf_5_10_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_20__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_158_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19105_ _19458_/A VGND VGND VPWR VPWR _19105_/X sky130_fd_sc_hd__buf_2
X_35151_ _35217_/CLK _35151_/D VGND VGND VPWR VPWR _35151_/Q sky130_fd_sc_hd__dfxtp_1
X_16317_ _33373_/Q _33309_/Q _33245_/Q _33181_/Q _16002_/X _16003_/X VGND VGND VPWR
+ VPWR _16317_/X sky130_fd_sc_hd__mux4_1
XFILLER_105_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17297_ _34424_/Q _36152_/Q _34296_/Q _34232_/Q _17229_/X _17230_/X VGND VGND VPWR
+ VPWR _17297_/X sky130_fd_sc_hd__mux4_1
X_32363_ _35946_/CLK _32363_/D VGND VGND VPWR VPWR _32363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_18_CLK clkbuf_6_4__f_CLK/X VGND VGND VPWR VPWR _35553_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_185_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34102_ _34166_/CLK _34102_/D VGND VGND VPWR VPWR _34102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16248_ _33883_/Q _33819_/Q _33755_/Q _36059_/Q _16112_/X _16113_/X VGND VGND VPWR
+ VPWR _16248_/X sky130_fd_sc_hd__mux4_1
X_19036_ _19032_/X _19035_/X _18759_/X VGND VGND VPWR VPWR _19037_/D sky130_fd_sc_hd__o21ba_1
X_31314_ _27686_/X _35876_/Q _31324_/S VGND VGND VPWR VPWR _31315_/A sky130_fd_sc_hd__mux2_1
X_35082_ _35212_/CLK _35082_/D VGND VGND VPWR VPWR _35082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32294_ _32552_/CLK _32294_/D VGND VGND VPWR VPWR _32294_/Q sky130_fd_sc_hd__dfxtp_1
X_31245_ _31245_/A VGND VGND VPWR VPWR _35843_/D sky130_fd_sc_hd__clkbuf_1
X_34033_ _35632_/CLK _34033_/D VGND VGND VPWR VPWR _34033_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput103 _31979_/Q VGND VGND VPWR VPWR D1[21] sky130_fd_sc_hd__buf_2
X_16179_ _34137_/Q _34073_/Q _34009_/Q _33945_/Q _16009_/X _16011_/X VGND VGND VPWR
+ VPWR _16179_/X sky130_fd_sc_hd__mux4_1
Xoutput114 _31989_/Q VGND VGND VPWR VPWR D1[31] sky130_fd_sc_hd__buf_2
XFILLER_86_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput125 _31999_/Q VGND VGND VPWR VPWR D1[41] sky130_fd_sc_hd__buf_2
Xoutput136 _32009_/Q VGND VGND VPWR VPWR D1[51] sky130_fd_sc_hd__buf_2
Xoutput147 _32019_/Q VGND VGND VPWR VPWR D1[61] sky130_fd_sc_hd__buf_2
Xoutput158 _36195_/Q VGND VGND VPWR VPWR D2[13] sky130_fd_sc_hd__buf_2
X_31176_ _31176_/A VGND VGND VPWR VPWR _35810_/D sky130_fd_sc_hd__clkbuf_1
Xoutput169 _36205_/Q VGND VGND VPWR VPWR D2[23] sky130_fd_sc_hd__buf_2
XFILLER_47_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30127_ _35314_/Q _29416_/X _30129_/S VGND VGND VPWR VPWR _30128_/A sky130_fd_sc_hd__mux2_1
X_19938_ _35714_/Q _32224_/Q _35586_/Q _35522_/Q _19617_/X _19618_/X VGND VGND VPWR
+ VPWR _19938_/X sky130_fd_sc_hd__mux4_1
XFILLER_138_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35984_ _35985_/CLK _35984_/D VGND VGND VPWR VPWR _35984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30058_ _30058_/A VGND VGND VPWR VPWR _35281_/D sky130_fd_sc_hd__clkbuf_1
X_34935_ _36151_/CLK _34935_/D VGND VGND VPWR VPWR _34935_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_233_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19869_ _32896_/Q _32832_/Q _32768_/Q _32704_/Q _19646_/X _19647_/X VGND VGND VPWR
+ VPWR _19869_/X sky130_fd_sc_hd__mux4_1
X_21900_ _21896_/X _21899_/X _21765_/X VGND VGND VPWR VPWR _21901_/D sky130_fd_sc_hd__o21ba_1
X_22880_ input88/X input87/X input86/X VGND VGND VPWR VPWR _22881_/A sky130_fd_sc_hd__or3_1
X_34866_ _35633_/CLK _34866_/D VGND VGND VPWR VPWR _34866_/Q sky130_fd_sc_hd__dfxtp_1
X_33817_ _34009_/CLK _33817_/D VGND VGND VPWR VPWR _33817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21831_ _34422_/Q _36150_/Q _34294_/Q _34230_/Q _21829_/X _21830_/X VGND VGND VPWR
+ VPWR _21831_/X sky130_fd_sc_hd__mux4_1
X_34797_ _34924_/CLK _34797_/D VGND VGND VPWR VPWR _34797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24550_ _24550_/A VGND VGND VPWR VPWR _32800_/D sky130_fd_sc_hd__clkbuf_1
X_33748_ _35669_/CLK _33748_/D VGND VGND VPWR VPWR _33748_/Q sky130_fd_sc_hd__dfxtp_1
X_21762_ _34932_/Q _34868_/Q _34804_/Q _34740_/Q _21760_/X _21761_/X VGND VGND VPWR
+ VPWR _21762_/X sky130_fd_sc_hd__mux4_1
XFILLER_149_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_954 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23501_ _32246_/Q _23396_/X _23515_/S VGND VGND VPWR VPWR _23502_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20713_ _22451_/A VGND VGND VPWR VPWR _20713_/X sky130_fd_sc_hd__buf_4
XFILLER_12_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24481_ _23018_/X _32768_/Q _24495_/S VGND VGND VPWR VPWR _24482_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33679_ _34440_/CLK _33679_/D VGND VGND VPWR VPWR _33679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_212_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21693_ _22560_/A VGND VGND VPWR VPWR _21693_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_211_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26220_ _26220_/A VGND VGND VPWR VPWR _33558_/D sky130_fd_sc_hd__clkbuf_1
X_35418_ _35802_/CLK _35418_/D VGND VGND VPWR VPWR _35418_/Q sky130_fd_sc_hd__dfxtp_1
X_23432_ input38/X VGND VGND VPWR VPWR _23432_/X sky130_fd_sc_hd__clkbuf_8
X_20644_ _22446_/A VGND VGND VPWR VPWR _20644_/X sky130_fd_sc_hd__buf_4
XFILLER_149_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26151_ _24899_/X _33526_/Q _26165_/S VGND VGND VPWR VPWR _26152_/A sky130_fd_sc_hd__mux2_1
X_35349_ _36055_/CLK _35349_/D VGND VGND VPWR VPWR _35349_/Q sky130_fd_sc_hd__dfxtp_1
X_23363_ _23363_/A VGND VGND VPWR VPWR _32197_/D sky130_fd_sc_hd__clkbuf_1
X_20575_ _18360_/X _20573_/X _20574_/X _18372_/X VGND VGND VPWR VPWR _20575_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25102_ _25102_/A VGND VGND VPWR VPWR _33031_/D sky130_fd_sc_hd__clkbuf_1
X_22314_ _22308_/X _22313_/X _22104_/X VGND VGND VPWR VPWR _22324_/C sky130_fd_sc_hd__o21ba_1
XFILLER_137_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26082_ _28380_/A _26352_/B VGND VGND VPWR VPWR _26215_/S sky130_fd_sc_hd__nand2_8
X_23294_ _32170_/Q _23292_/X _23424_/S VGND VGND VPWR VPWR _23295_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29910_ _35211_/Q _29494_/X _29922_/S VGND VGND VPWR VPWR _29911_/A sky130_fd_sc_hd__mux2_1
XFILLER_191_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25033_ _25033_/A VGND VGND VPWR VPWR _32998_/D sky130_fd_sc_hd__clkbuf_1
X_22245_ _22598_/A VGND VGND VPWR VPWR _22245_/X sky130_fd_sc_hd__buf_6
XFILLER_117_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29841_ _35178_/Q _29391_/X _29859_/S VGND VGND VPWR VPWR _29842_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22176_ _33088_/Q _32064_/Q _35840_/Q _35776_/Q _22031_/X _22032_/X VGND VGND VPWR
+ VPWR _22176_/X sky130_fd_sc_hd__mux4_1
XFILLER_156_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21127_ _21052_/X _21125_/X _21126_/X _21057_/X VGND VGND VPWR VPWR _21127_/X sky130_fd_sc_hd__a22o_1
X_29772_ _29772_/A VGND VGND VPWR VPWR _35145_/D sky130_fd_sc_hd__clkbuf_1
X_26984_ _33918_/Q _23420_/X _27002_/S VGND VGND VPWR VPWR _26985_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28723_ _28723_/A VGND VGND VPWR VPWR _34679_/D sky130_fd_sc_hd__clkbuf_1
X_25935_ _24979_/X _33424_/Q _25937_/S VGND VGND VPWR VPWR _25936_/A sky130_fd_sc_hd__mux2_1
X_21058_ _21052_/X _21053_/X _21056_/X _21057_/X VGND VGND VPWR VPWR _21058_/X sky130_fd_sc_hd__a22o_1
XFILLER_93_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_1131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20009_ _20164_/A VGND VGND VPWR VPWR _20009_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_246_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28654_ _28654_/A VGND VGND VPWR VPWR _34646_/D sky130_fd_sc_hd__clkbuf_1
X_25866_ _24877_/X _33391_/Q _25874_/S VGND VGND VPWR VPWR _25867_/A sky130_fd_sc_hd__mux2_1
XFILLER_219_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27605_ _27605_/A VGND VGND VPWR VPWR _34181_/D sky130_fd_sc_hd__clkbuf_1
X_24817_ _24817_/A VGND VGND VPWR VPWR _32923_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25797_ _25797_/A VGND VGND VPWR VPWR _33358_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28585_ _28585_/A VGND VGND VPWR VPWR _34614_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24748_ _24748_/A VGND VGND VPWR VPWR _32894_/D sky130_fd_sc_hd__clkbuf_1
X_27536_ _27536_/A VGND VGND VPWR VPWR _34148_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27467_ _34116_/Q _27177_/X _27473_/S VGND VGND VPWR VPWR _27468_/A sky130_fd_sc_hd__mux2_1
XFILLER_203_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24679_ _22912_/X _32862_/Q _24681_/S VGND VGND VPWR VPWR _24680_/A sky130_fd_sc_hd__mux2_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29206_ _29206_/A VGND VGND VPWR VPWR _34907_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_208_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17220_ _35638_/Q _34998_/Q _34358_/Q _33718_/Q _17144_/X _17145_/X VGND VGND VPWR
+ VPWR _17220_/X sky130_fd_sc_hd__mux4_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26418_ _33652_/Q _23387_/X _26436_/S VGND VGND VPWR VPWR _26419_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27398_ _34083_/Q _27075_/X _27410_/S VGND VGND VPWR VPWR _27399_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17151_ _17857_/A VGND VGND VPWR VPWR _17151_/X sky130_fd_sc_hd__buf_4
X_26349_ _26349_/A VGND VGND VPWR VPWR _33620_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_862 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29137_ _34875_/Q _27149_/X _29141_/S VGND VGND VPWR VPWR _29138_/A sky130_fd_sc_hd__mux2_1
Xinput16 DW[23] VGND VGND VPWR VPWR input16/X sky130_fd_sc_hd__buf_4
XFILLER_122_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput27 DW[33] VGND VGND VPWR VPWR input27/X sky130_fd_sc_hd__clkbuf_4
X_16102_ _16091_/X _16095_/X _16099_/X _16101_/X VGND VGND VPWR VPWR _16102_/X sky130_fd_sc_hd__a22o_1
XFILLER_11_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput38 DW[43] VGND VGND VPWR VPWR input38/X sky130_fd_sc_hd__buf_6
X_29068_ _34842_/Q _27047_/X _29078_/S VGND VGND VPWR VPWR _29069_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput49 DW[53] VGND VGND VPWR VPWR input49/X sky130_fd_sc_hd__clkbuf_16
X_17082_ _17076_/X _17081_/X _16798_/X VGND VGND VPWR VPWR _17090_/C sky130_fd_sc_hd__o21ba_1
XFILLER_196_1135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16033_ _16063_/A VGND VGND VPWR VPWR _17774_/A sky130_fd_sc_hd__buf_8
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28019_ _34346_/Q _27096_/X _28037_/S VGND VGND VPWR VPWR _28020_/A sky130_fd_sc_hd__mux2_1
XFILLER_237_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31030_ _35742_/Q input63/X _31032_/S VGND VGND VPWR VPWR _31031_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17984_ _33164_/Q _36044_/Q _33036_/Q _32972_/Q _17768_/X _17769_/X VGND VGND VPWR
+ VPWR _17984_/X sky130_fd_sc_hd__mux4_1
XFILLER_46_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19723_ _32892_/Q _32828_/Q _32764_/Q _32700_/Q _19646_/X _19647_/X VGND VGND VPWR
+ VPWR _19723_/X sky130_fd_sc_hd__mux4_1
XFILLER_111_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16935_ _35438_/Q _35374_/Q _35310_/Q _35246_/Q _16901_/X _16902_/X VGND VGND VPWR
+ VPWR _16935_/X sky130_fd_sc_hd__mux4_1
XFILLER_238_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32981_ _36052_/CLK _32981_/D VGND VGND VPWR VPWR _32981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_1163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34720_ _34914_/CLK _34720_/D VGND VGND VPWR VPWR _34720_/Q sky130_fd_sc_hd__dfxtp_1
X_31932_ _23460_/X _36169_/Q _31948_/S VGND VGND VPWR VPWR _31933_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19654_ _20162_/A VGND VGND VPWR VPWR _19654_/X sky130_fd_sc_hd__buf_6
X_16866_ _35692_/Q _32200_/Q _35564_/Q _35500_/Q _16611_/X _16612_/X VGND VGND VPWR
+ VPWR _16866_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_7_CLK clkbuf_leaf_9_CLK/A VGND VGND VPWR VPWR _34915_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_225_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18605_ _19311_/A VGND VGND VPWR VPWR _18605_/X sky130_fd_sc_hd__buf_6
X_34651_ _35544_/CLK _34651_/D VGND VGND VPWR VPWR _34651_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19585_ _35704_/Q _32213_/Q _35576_/Q _35512_/Q _19264_/X _19265_/X VGND VGND VPWR
+ VPWR _19585_/X sky130_fd_sc_hd__mux4_1
X_31863_ _31863_/A VGND VGND VPWR VPWR _36136_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16797_ _16650_/X _16795_/X _16796_/X _16653_/X VGND VGND VPWR VPWR _16797_/X sky130_fd_sc_hd__a22o_1
XFILLER_53_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33602_ _36161_/CLK _33602_/D VGND VGND VPWR VPWR _33602_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_248_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18536_ _35162_/Q _35098_/Q _35034_/Q _32154_/Q _18383_/X _18385_/X VGND VGND VPWR
+ VPWR _18536_/X sky130_fd_sc_hd__mux4_1
X_30814_ _30814_/A VGND VGND VPWR VPWR _35639_/D sky130_fd_sc_hd__clkbuf_1
X_34582_ _34647_/CLK _34582_/D VGND VGND VPWR VPWR _34582_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31794_ _31821_/S VGND VGND VPWR VPWR _31813_/S sky130_fd_sc_hd__buf_4
XFILLER_244_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33533_ _33661_/CLK _33533_/D VGND VGND VPWR VPWR _33533_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18467_ _34648_/Q _34584_/Q _34520_/Q _34456_/Q _18379_/X _18380_/X VGND VGND VPWR
+ VPWR _18467_/X sky130_fd_sc_hd__mux4_1
X_30745_ _30745_/A VGND VGND VPWR VPWR _35606_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17418_ _17910_/A VGND VGND VPWR VPWR _17418_/X sky130_fd_sc_hd__clkbuf_4
X_33464_ _33850_/CLK _33464_/D VGND VGND VPWR VPWR _33464_/Q sky130_fd_sc_hd__dfxtp_1
X_18398_ _19461_/A VGND VGND VPWR VPWR _18398_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_194_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30676_ _35574_/Q _29429_/X _30690_/S VGND VGND VPWR VPWR _30677_/A sky130_fd_sc_hd__mux2_1
X_35203_ _35655_/CLK _35203_/D VGND VGND VPWR VPWR _35203_/Q sky130_fd_sc_hd__dfxtp_1
X_32415_ _33573_/CLK _32415_/D VGND VGND VPWR VPWR _32415_/Q sky130_fd_sc_hd__dfxtp_1
X_36183_ _36191_/CLK _36183_/D VGND VGND VPWR VPWR _36183_/Q sky130_fd_sc_hd__dfxtp_1
X_17349_ _17067_/X _17345_/X _17348_/X _17071_/X VGND VGND VPWR VPWR _17349_/X sky130_fd_sc_hd__a22o_1
X_33395_ _36082_/CLK _33395_/D VGND VGND VPWR VPWR _33395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35134_ _36099_/CLK _35134_/D VGND VGND VPWR VPWR _35134_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20360_ _34702_/Q _34638_/Q _34574_/Q _34510_/Q _20298_/X _20299_/X VGND VGND VPWR
+ VPWR _20360_/X sky130_fd_sc_hd__mux4_1
X_32346_ _35995_/CLK _32346_/D VGND VGND VPWR VPWR _32346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19019_ _19014_/X _19016_/X _19017_/X _19018_/X VGND VGND VPWR VPWR _19019_/X sky130_fd_sc_hd__a22o_1
X_20291_ _35724_/Q _32235_/Q _35596_/Q _35532_/Q _19970_/X _19971_/X VGND VGND VPWR
+ VPWR _20291_/X sky130_fd_sc_hd__mux4_1
X_35065_ _35191_/CLK _35065_/D VGND VGND VPWR VPWR _35065_/Q sky130_fd_sc_hd__dfxtp_1
X_32277_ _35221_/CLK _32277_/D VGND VGND VPWR VPWR _32277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22030_ _35452_/Q _35388_/Q _35324_/Q _35260_/Q _21854_/X _21855_/X VGND VGND VPWR
+ VPWR _22030_/X sky130_fd_sc_hd__mux4_1
X_34016_ _36209_/CLK _34016_/D VGND VGND VPWR VPWR _34016_/Q sky130_fd_sc_hd__dfxtp_1
X_31228_ _31228_/A VGND VGND VPWR VPWR _35835_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31159_ _31159_/A VGND VGND VPWR VPWR _35802_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_248_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23981_ _24113_/S VGND VGND VPWR VPWR _24000_/S sky130_fd_sc_hd__buf_6
X_35967_ _36031_/CLK _35967_/D VGND VGND VPWR VPWR _35967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25720_ _25810_/S VGND VGND VPWR VPWR _25739_/S sky130_fd_sc_hd__buf_4
XFILLER_69_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34918_ _34918_/CLK _34918_/D VGND VGND VPWR VPWR _34918_/Q sky130_fd_sc_hd__dfxtp_1
X_22932_ _22931_/X _32036_/Q _22947_/S VGND VGND VPWR VPWR _22933_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35898_ _35962_/CLK _35898_/D VGND VGND VPWR VPWR _35898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_244_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25651_ _24958_/X _33289_/Q _25667_/S VGND VGND VPWR VPWR _25652_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22863_ _35733_/Q _32245_/Q _35605_/Q _35541_/Q _20593_/X _20595_/X VGND VGND VPWR
+ VPWR _22863_/X sky130_fd_sc_hd__mux4_1
X_34849_ _34913_/CLK _34849_/D VGND VGND VPWR VPWR _34849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24602_ _24602_/A VGND VGND VPWR VPWR _32825_/D sky130_fd_sc_hd__clkbuf_1
X_28370_ _27825_/X _34513_/Q _28370_/S VGND VGND VPWR VPWR _28371_/A sky130_fd_sc_hd__mux2_1
X_21814_ _21659_/X _21812_/X _21813_/X _21665_/X VGND VGND VPWR VPWR _21814_/X sky130_fd_sc_hd__a22o_1
X_25582_ _25582_/A VGND VGND VPWR VPWR _33256_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22794_ _22512_/X _22792_/X _22793_/X _22515_/X VGND VGND VPWR VPWR _22794_/X sky130_fd_sc_hd__a22o_1
XFILLER_19_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27321_ _27321_/A VGND VGND VPWR VPWR _34046_/D sky130_fd_sc_hd__clkbuf_1
X_24533_ _24533_/A VGND VGND VPWR VPWR _32792_/D sky130_fd_sc_hd__clkbuf_1
XPHY_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21745_ _22599_/A VGND VGND VPWR VPWR _21745_/X sky130_fd_sc_hd__buf_4
XFILLER_197_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27252_ _34014_/Q _27059_/X _27254_/S VGND VGND VPWR VPWR _27253_/A sky130_fd_sc_hd__mux2_1
X_24464_ _22993_/X _32760_/Q _24474_/S VGND VGND VPWR VPWR _24465_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21676_ _21598_/X _21674_/X _21675_/X _21601_/X VGND VGND VPWR VPWR _21676_/X sky130_fd_sc_hd__a22o_1
XFILLER_145_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26203_ _24976_/X _33551_/Q _26207_/S VGND VGND VPWR VPWR _26204_/A sky130_fd_sc_hd__mux2_1
XFILLER_200_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23415_ _32217_/Q _23414_/X _23418_/S VGND VGND VPWR VPWR _23416_/A sky130_fd_sc_hd__mux2_1
X_20627_ _22510_/A VGND VGND VPWR VPWR _20627_/X sky130_fd_sc_hd__clkbuf_4
X_27183_ input43/X VGND VGND VPWR VPWR _27183_/X sky130_fd_sc_hd__buf_4
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24395_ _22891_/X _32727_/Q _24411_/S VGND VGND VPWR VPWR _24396_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26134_ _24874_/X _33518_/Q _26144_/S VGND VGND VPWR VPWR _26135_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23346_ _23346_/A VGND VGND VPWR VPWR _32189_/D sky130_fd_sc_hd__clkbuf_1
X_20558_ _19453_/A _20556_/X _20557_/X _19456_/A VGND VGND VPWR VPWR _20558_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26065_ _26065_/A VGND VGND VPWR VPWR _33485_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23277_ input7/X VGND VGND VPWR VPWR _23277_/X sky130_fd_sc_hd__buf_6
X_20489_ _33683_/Q _33619_/Q _33555_/Q _33491_/Q _20206_/X _20207_/X VGND VGND VPWR
+ VPWR _20489_/X sky130_fd_sc_hd__mux4_1
XFILLER_180_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25016_ _25016_/A VGND VGND VPWR VPWR _32990_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22228_ _22224_/X _22227_/X _22085_/X VGND VGND VPWR VPWR _22254_/A sky130_fd_sc_hd__o21ba_1
XFILLER_65_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29824_ _35170_/Q _29367_/X _29838_/S VGND VGND VPWR VPWR _29825_/A sky130_fd_sc_hd__mux2_1
X_22159_ _22512_/A VGND VGND VPWR VPWR _22159_/X sky130_fd_sc_hd__buf_4
XFILLER_117_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29755_ _29755_/A VGND VGND VPWR VPWR _35137_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26967_ _33910_/Q _23396_/X _26981_/S VGND VGND VPWR VPWR _26968_/A sky130_fd_sc_hd__mux2_1
XTAP_6899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28706_ _28706_/A VGND VGND VPWR VPWR _34671_/D sky130_fd_sc_hd__clkbuf_1
X_16720_ _16713_/X _16719_/X _16434_/X _16435_/X VGND VGND VPWR VPWR _16737_/B sky130_fd_sc_hd__o211a_1
X_25918_ _25945_/S VGND VGND VPWR VPWR _25937_/S sky130_fd_sc_hd__buf_4
XFILLER_219_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29686_ _29686_/A VGND VGND VPWR VPWR _35104_/D sky130_fd_sc_hd__clkbuf_1
X_26898_ _30337_/A _31688_/B VGND VGND VPWR VPWR _27031_/S sky130_fd_sc_hd__nor2_8
XFILLER_247_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28637_ _28637_/A VGND VGND VPWR VPWR _34639_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16651_ _35430_/Q _35366_/Q _35302_/Q _35238_/Q _16548_/X _16549_/X VGND VGND VPWR
+ VPWR _16651_/X sky130_fd_sc_hd__mux4_1
XFILLER_74_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25849_ _24852_/X _33383_/Q _25853_/S VGND VGND VPWR VPWR _25850_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19370_ _32882_/Q _32818_/Q _32754_/Q _32690_/Q _19293_/X _19294_/X VGND VGND VPWR
+ VPWR _19370_/X sky130_fd_sc_hd__mux4_1
X_28568_ _28568_/A VGND VGND VPWR VPWR _34606_/D sky130_fd_sc_hd__clkbuf_1
X_16582_ _35428_/Q _35364_/Q _35300_/Q _35236_/Q _16548_/X _16549_/X VGND VGND VPWR
+ VPWR _16582_/X sky130_fd_sc_hd__mux4_1
XFILLER_188_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18321_ _18363_/A VGND VGND VPWR VPWR _20066_/A sky130_fd_sc_hd__buf_12
XFILLER_231_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27519_ _27519_/A VGND VGND VPWR VPWR _34140_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28499_ _27816_/X _34574_/Q _28505_/S VGND VGND VPWR VPWR _28500_/A sky130_fd_sc_hd__mux2_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18252_ _33429_/Q _33365_/Q _33301_/Q _33237_/Q _16037_/X _16039_/X VGND VGND VPWR
+ VPWR _18252_/X sky130_fd_sc_hd__mux4_1
XFILLER_179_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30530_ _35505_/Q _29413_/X _30534_/S VGND VGND VPWR VPWR _30531_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17203_ _34166_/Q _34102_/Q _34038_/Q _33974_/Q _17093_/X _17094_/X VGND VGND VPWR
+ VPWR _17203_/X sky130_fd_sc_hd__mux4_1
X_30461_ _30461_/A VGND VGND VPWR VPWR _35472_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18183_ _34450_/Q _36178_/Q _34322_/Q _34258_/Q _17935_/X _17936_/X VGND VGND VPWR
+ VPWR _18183_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32200_ _35564_/CLK _32200_/D VGND VGND VPWR VPWR _32200_/Q sky130_fd_sc_hd__dfxtp_1
X_17134_ _32628_/Q _32564_/Q _32500_/Q _35956_/Q _16923_/X _17060_/X VGND VGND VPWR
+ VPWR _17134_/X sky130_fd_sc_hd__mux4_1
X_33180_ _33818_/CLK _33180_/D VGND VGND VPWR VPWR _33180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30392_ _30392_/A VGND VGND VPWR VPWR _35439_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_5_7_0_CLK clkbuf_5_7_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_7_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_144_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32131_ _35907_/CLK _32131_/D VGND VGND VPWR VPWR _32131_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17065_ _17910_/A VGND VGND VPWR VPWR _17065_/X sky130_fd_sc_hd__clkbuf_4
X_16016_ _15997_/X _16013_/X _16015_/X VGND VGND VPWR VPWR _16106_/A sky130_fd_sc_hd__o21ba_1
XFILLER_170_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32062_ _32575_/CLK _32062_/D VGND VGND VPWR VPWR _32062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31013_ _31145_/S VGND VGND VPWR VPWR _31032_/S sky130_fd_sc_hd__buf_6
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35821_ _36141_/CLK _35821_/D VGND VGND VPWR VPWR _35821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17967_ _35211_/Q _35147_/Q _35083_/Q _32267_/Q _17716_/X _17717_/X VGND VGND VPWR
+ VPWR _17967_/X sky130_fd_sc_hd__mux4_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19706_ _34172_/Q _34108_/Q _34044_/Q _33980_/Q _19393_/X _19394_/X VGND VGND VPWR
+ VPWR _19706_/X sky130_fd_sc_hd__mux4_1
X_16918_ _16846_/X _16916_/X _16917_/X _16851_/X VGND VGND VPWR VPWR _16918_/X sky130_fd_sc_hd__a22o_1
X_35752_ _35817_/CLK _35752_/D VGND VGND VPWR VPWR _35752_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32964_ _36038_/CLK _32964_/D VGND VGND VPWR VPWR _32964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17898_ _17859_/X _17896_/X _17897_/X _17862_/X VGND VGND VPWR VPWR _17898_/X sky130_fd_sc_hd__a22o_1
XFILLER_226_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34703_ _35147_/CLK _34703_/D VGND VGND VPWR VPWR _34703_/Q sky130_fd_sc_hd__dfxtp_1
X_31915_ _23432_/X _36161_/Q _31927_/S VGND VGND VPWR VPWR _31916_/A sky130_fd_sc_hd__mux2_1
X_19637_ _19499_/X _19635_/X _19636_/X _19504_/X VGND VGND VPWR VPWR _19637_/X sky130_fd_sc_hd__a22o_1
X_16849_ _33644_/Q _33580_/Q _33516_/Q _33452_/Q _16847_/X _16848_/X VGND VGND VPWR
+ VPWR _16849_/X sky130_fd_sc_hd__mux4_1
X_35683_ _35684_/CLK _35683_/D VGND VGND VPWR VPWR _35683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32895_ _32895_/CLK _32895_/D VGND VGND VPWR VPWR _32895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34634_ _35210_/CLK _34634_/D VGND VGND VPWR VPWR _34634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19568_ _19568_/A VGND VGND VPWR VPWR _32439_/D sky130_fd_sc_hd__buf_2
X_31846_ _23261_/X _36128_/Q _31864_/S VGND VGND VPWR VPWR _31847_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_248_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18519_ _33114_/Q _35994_/Q _32986_/Q _32922_/Q _18324_/X _18325_/X VGND VGND VPWR
+ VPWR _18519_/X sky130_fd_sc_hd__mux4_1
X_34565_ _34694_/CLK _34565_/D VGND VGND VPWR VPWR _34565_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31777_ _31777_/A VGND VGND VPWR VPWR _36095_/D sky130_fd_sc_hd__clkbuf_1
X_19499_ _20205_/A VGND VGND VPWR VPWR _19499_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_90_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33516_ _34093_/CLK _33516_/D VGND VGND VPWR VPWR _33516_/Q sky130_fd_sc_hd__dfxtp_1
X_21530_ _21314_/X _21528_/X _21529_/X _21318_/X VGND VGND VPWR VPWR _21530_/X sky130_fd_sc_hd__a22o_1
X_30728_ _35599_/Q _29506_/X _30732_/S VGND VGND VPWR VPWR _30729_/A sky130_fd_sc_hd__mux2_1
X_34496_ _34690_/CLK _34496_/D VGND VGND VPWR VPWR _34496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36235_ _36235_/CLK _36235_/D VGND VGND VPWR VPWR _36235_/Q sky130_fd_sc_hd__dfxtp_1
X_33447_ _36068_/CLK _33447_/D VGND VGND VPWR VPWR _33447_/Q sky130_fd_sc_hd__dfxtp_1
X_21461_ _21306_/X _21459_/X _21460_/X _21312_/X VGND VGND VPWR VPWR _21461_/X sky130_fd_sc_hd__a22o_1
X_30659_ _35566_/Q _29404_/X _30669_/S VGND VGND VPWR VPWR _30660_/A sky130_fd_sc_hd__mux2_1
X_23200_ _23200_/A VGND VGND VPWR VPWR _32137_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20412_ _20408_/X _20411_/X _20146_/X _20147_/X VGND VGND VPWR VPWR _20427_/B sky130_fd_sc_hd__o211a_1
XFILLER_105_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36166_ _36167_/CLK _36166_/D VGND VGND VPWR VPWR _36166_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24180_ _32627_/Q _23384_/X _24180_/S VGND VGND VPWR VPWR _24181_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33378_ _33828_/CLK _33378_/D VGND VGND VPWR VPWR _33378_/Q sky130_fd_sc_hd__dfxtp_1
X_21392_ _22599_/A VGND VGND VPWR VPWR _21392_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_105_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35117_ _35181_/CLK _35117_/D VGND VGND VPWR VPWR _35117_/Q sky130_fd_sc_hd__dfxtp_1
X_23131_ _22946_/X _32105_/Q _23131_/S VGND VGND VPWR VPWR _23132_/A sky130_fd_sc_hd__mux2_1
X_20343_ _33934_/Q _33870_/Q _33806_/Q _36110_/Q _20030_/X _20031_/X VGND VGND VPWR
+ VPWR _20343_/X sky130_fd_sc_hd__mux4_1
XFILLER_134_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32329_ _35978_/CLK _32329_/D VGND VGND VPWR VPWR _32329_/Q sky130_fd_sc_hd__dfxtp_1
X_36097_ _36097_/CLK _36097_/D VGND VGND VPWR VPWR _36097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23062_ _23061_/X _32078_/Q _23071_/S VGND VGND VPWR VPWR _23063_/A sky130_fd_sc_hd__mux2_1
X_35048_ _35176_/CLK _35048_/D VGND VGND VPWR VPWR _35048_/Q sky130_fd_sc_hd__dfxtp_1
X_20274_ _20274_/A VGND VGND VPWR VPWR _32459_/D sky130_fd_sc_hd__clkbuf_4
XTAP_6107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22013_ _22366_/A VGND VGND VPWR VPWR _22013_/X sky130_fd_sc_hd__buf_4
XTAP_6129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27870_ _27870_/A VGND VGND VPWR VPWR _34275_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1057 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26821_ _33841_/Q _23364_/X _26825_/S VGND VGND VPWR VPWR _26822_/A sky130_fd_sc_hd__mux2_1
XTAP_5439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29540_ _29540_/A VGND VGND VPWR VPWR _35035_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26752_ _26752_/A VGND VGND VPWR VPWR _33808_/D sky130_fd_sc_hd__clkbuf_1
X_23964_ _23964_/A VGND VGND VPWR VPWR _32526_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22915_ input64/X VGND VGND VPWR VPWR _22915_/X sky130_fd_sc_hd__buf_2
X_25703_ _25703_/A VGND VGND VPWR VPWR _33313_/D sky130_fd_sc_hd__clkbuf_1
X_29471_ _29471_/A VGND VGND VPWR VPWR _35011_/D sky130_fd_sc_hd__clkbuf_1
X_26683_ _26683_/A VGND VGND VPWR VPWR _33775_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23895_ _23895_/A VGND VGND VPWR VPWR _32493_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28422_ _28422_/A VGND VGND VPWR VPWR _34537_/D sky130_fd_sc_hd__clkbuf_1
X_22846_ _22842_/X _22845_/X _22471_/A VGND VGND VPWR VPWR _22847_/D sky130_fd_sc_hd__o21ba_1
X_25634_ _24933_/X _33281_/Q _25646_/S VGND VGND VPWR VPWR _25635_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_244_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28353_ _28353_/A VGND VGND VPWR VPWR _34504_/D sky130_fd_sc_hd__clkbuf_1
X_25565_ _24830_/X _33248_/Q _25583_/S VGND VGND VPWR VPWR _25566_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22777_ _33106_/Q _32082_/Q _35858_/Q _35794_/Q _20679_/X _20680_/X VGND VGND VPWR
+ VPWR _22777_/X sky130_fd_sc_hd__mux4_1
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_240_CLK clkbuf_6_61__f_CLK/X VGND VGND VPWR VPWR _34949_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_890 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24516_ _23070_/X _32785_/Q _24516_/S VGND VGND VPWR VPWR _24517_/A sky130_fd_sc_hd__mux2_1
X_27304_ _27304_/A VGND VGND VPWR VPWR _34038_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21728_ _22434_/A VGND VGND VPWR VPWR _21728_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_38_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25496_ _25496_/A VGND VGND VPWR VPWR _33215_/D sky130_fd_sc_hd__clkbuf_1
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28284_ _27698_/X _34472_/Q _28286_/S VGND VGND VPWR VPWR _28285_/A sky130_fd_sc_hd__mux2_1
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27235_ _27367_/S VGND VGND VPWR VPWR _27254_/S sky130_fd_sc_hd__buf_6
X_24447_ _22968_/X _32752_/Q _24453_/S VGND VGND VPWR VPWR _24448_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21659_ _22505_/A VGND VGND VPWR VPWR _21659_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_12_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27166_ _33984_/Q _27165_/X _27187_/S VGND VGND VPWR VPWR _27167_/A sky130_fd_sc_hd__mux2_1
X_24378_ _24378_/A VGND VGND VPWR VPWR _32719_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26117_ _24849_/X _33510_/Q _26123_/S VGND VGND VPWR VPWR _26118_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23329_ _32182_/Q _23249_/X _23335_/S VGND VGND VPWR VPWR _23330_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27097_ _27230_/S VGND VGND VPWR VPWR _27125_/S sky130_fd_sc_hd__buf_4
XFILLER_67_1108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26048_ _26048_/A VGND VGND VPWR VPWR _33477_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18870_ _20282_/A VGND VGND VPWR VPWR _18870_/X sky130_fd_sc_hd__buf_6
XTAP_6630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29807_ _35162_/Q _29342_/X _29817_/S VGND VGND VPWR VPWR _29808_/A sky130_fd_sc_hd__mux2_1
X_17821_ _34695_/Q _34631_/Q _34567_/Q _34503_/Q _17645_/X _17646_/X VGND VGND VPWR
+ VPWR _17821_/X sky130_fd_sc_hd__mux4_1
XTAP_6663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27999_ _27999_/A VGND VGND VPWR VPWR _34336_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17752_ _34437_/Q _36165_/Q _34309_/Q _34245_/Q _17582_/X _17583_/X VGND VGND VPWR
+ VPWR _17752_/X sky130_fd_sc_hd__mux4_1
XFILLER_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29738_ _29738_/A VGND VGND VPWR VPWR _35129_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16703_ _33896_/Q _33832_/Q _33768_/Q _36072_/Q _16671_/X _16672_/X VGND VGND VPWR
+ VPWR _16703_/X sky130_fd_sc_hd__mux4_1
X_29669_ _29669_/A VGND VGND VPWR VPWR _35096_/D sky130_fd_sc_hd__clkbuf_1
X_17683_ _34947_/Q _34883_/Q _34819_/Q _34755_/Q _17513_/X _17514_/X VGND VGND VPWR
+ VPWR _17683_/X sky130_fd_sc_hd__mux4_1
XFILLER_75_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31700_ _36059_/Q input56/X _31708_/S VGND VGND VPWR VPWR _31701_/A sky130_fd_sc_hd__mux2_1
X_19422_ _19422_/A _19422_/B _19422_/C _19422_/D VGND VGND VPWR VPWR _19423_/A sky130_fd_sc_hd__or4_4
X_16634_ _16500_/X _16632_/X _16633_/X _16503_/X VGND VGND VPWR VPWR _16634_/X sky130_fd_sc_hd__a22o_1
XFILLER_207_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32680_ _32871_/CLK _32680_/D VGND VGND VPWR VPWR _32680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19353_ _34162_/Q _34098_/Q _34034_/Q _33970_/Q _19040_/X _19041_/X VGND VGND VPWR
+ VPWR _19353_/X sky130_fd_sc_hd__mux4_1
X_31631_ _31631_/A VGND VGND VPWR VPWR _36026_/D sky130_fd_sc_hd__clkbuf_1
X_16565_ _16493_/X _16563_/X _16564_/X _16498_/X VGND VGND VPWR VPWR _16565_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_231_CLK clkbuf_6_55__f_CLK/X VGND VGND VPWR VPWR _33869_/CLK sky130_fd_sc_hd__clkbuf_16
X_18304_ _33366_/Q _33302_/Q _33238_/Q _33174_/Q _18302_/X _18303_/X VGND VGND VPWR
+ VPWR _18304_/X sky130_fd_sc_hd__mux4_1
X_34350_ _35694_/CLK _34350_/D VGND VGND VPWR VPWR _34350_/Q sky130_fd_sc_hd__dfxtp_1
X_31562_ _31562_/A VGND VGND VPWR VPWR _35993_/D sky130_fd_sc_hd__clkbuf_1
X_19284_ _19146_/X _19282_/X _19283_/X _19151_/X VGND VGND VPWR VPWR _19284_/X sky130_fd_sc_hd__a22o_1
XFILLER_31_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16496_ _33634_/Q _33570_/Q _33506_/Q _33442_/Q _16494_/X _16495_/X VGND VGND VPWR
+ VPWR _16496_/X sky130_fd_sc_hd__mux4_1
XFILLER_206_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33301_ _33685_/CLK _33301_/D VGND VGND VPWR VPWR _33301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18235_ _15981_/X _18233_/X _18234_/X _15991_/X VGND VGND VPWR VPWR _18235_/X sky130_fd_sc_hd__a22o_1
XFILLER_175_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30513_ _35497_/Q _29388_/X _30513_/S VGND VGND VPWR VPWR _30514_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34281_ _34915_/CLK _34281_/D VGND VGND VPWR VPWR _34281_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31493_ _27751_/X _35961_/Q _31501_/S VGND VGND VPWR VPWR _31494_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36020_ _36020_/CLK _36020_/D VGND VGND VPWR VPWR _36020_/Q sky130_fd_sc_hd__dfxtp_1
X_33232_ _34186_/CLK _33232_/D VGND VGND VPWR VPWR _33232_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30444_ _35464_/Q _29484_/X _30462_/S VGND VGND VPWR VPWR _30445_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18166_ _32658_/Q _32594_/Q _32530_/Q _35986_/Q _17982_/X _16877_/A VGND VGND VPWR
+ VPWR _18166_/X sky130_fd_sc_hd__mux4_1
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17117_ _16800_/X _17115_/X _17116_/X _16803_/X VGND VGND VPWR VPWR _17117_/X sky130_fd_sc_hd__a22o_1
XFILLER_171_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33163_ _36044_/CLK _33163_/D VGND VGND VPWR VPWR _33163_/Q sky130_fd_sc_hd__dfxtp_1
X_18097_ _18097_/A _18097_/B _18097_/C _18097_/D VGND VGND VPWR VPWR _18098_/A sky130_fd_sc_hd__or4_2
XFILLER_144_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30375_ _30375_/A VGND VGND VPWR VPWR _35431_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_239_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32114_ _32882_/CLK _32114_/D VGND VGND VPWR VPWR _32114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1079 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17048_ _16805_/X _17046_/X _17047_/X _16810_/X VGND VGND VPWR VPWR _17048_/X sky130_fd_sc_hd__a22o_1
X_33094_ _35845_/CLK _33094_/D VGND VGND VPWR VPWR _33094_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_298_CLK clkbuf_6_57__f_CLK/X VGND VGND VPWR VPWR _35841_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_48_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32045_ _35822_/CLK _32045_/D VGND VGND VPWR VPWR _32045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1074 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_1366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18999_ _33640_/Q _33576_/Q _33512_/Q _33448_/Q _18794_/X _18795_/X VGND VGND VPWR
+ VPWR _18999_/X sky130_fd_sc_hd__mux4_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35804_ _35804_/CLK _35804_/D VGND VGND VPWR VPWR _35804_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33996_ _34188_/CLK _33996_/D VGND VGND VPWR VPWR _33996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35735_ _35735_/CLK _35735_/D VGND VGND VPWR VPWR _35735_/Q sky130_fd_sc_hd__dfxtp_1
X_20961_ _22512_/A VGND VGND VPWR VPWR _20961_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_54_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32947_ _36019_/CLK _32947_/D VGND VGND VPWR VPWR _32947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22700_ _34192_/Q _34128_/Q _34064_/Q _34000_/Q _22399_/X _22400_/X VGND VGND VPWR
+ VPWR _22700_/X sky130_fd_sc_hd__mux4_1
XFILLER_187_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_470_CLK clkbuf_6_11__f_CLK/X VGND VGND VPWR VPWR _35694_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_54_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35666_ _35666_/CLK _35666_/D VGND VGND VPWR VPWR _35666_/Q sky130_fd_sc_hd__dfxtp_1
X_23680_ _23049_/X _32330_/Q _23694_/S VGND VGND VPWR VPWR _23681_/A sky130_fd_sc_hd__mux2_1
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20892_ _22459_/A VGND VGND VPWR VPWR _20892_/X sky130_fd_sc_hd__buf_4
X_32878_ _32911_/CLK _32878_/D VGND VGND VPWR VPWR _32878_/Q sky130_fd_sc_hd__dfxtp_1
X_22631_ _35213_/Q _35149_/Q _35085_/Q _32269_/Q _22316_/X _22317_/X VGND VGND VPWR
+ VPWR _22631_/X sky130_fd_sc_hd__mux4_1
X_34617_ _35193_/CLK _34617_/D VGND VGND VPWR VPWR _34617_/Q sky130_fd_sc_hd__dfxtp_1
X_31829_ _23237_/X _36120_/Q _31843_/S VGND VGND VPWR VPWR _31830_/A sky130_fd_sc_hd__mux2_1
X_35597_ _35727_/CLK _35597_/D VGND VGND VPWR VPWR _35597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_1072 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_222_CLK clkbuf_6_53__f_CLK/X VGND VGND VPWR VPWR _34957_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_34_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25350_ _25350_/A VGND VGND VPWR VPWR _33147_/D sky130_fd_sc_hd__clkbuf_1
X_22562_ _35467_/Q _35403_/Q _35339_/Q _35275_/Q _22560_/X _22561_/X VGND VGND VPWR
+ VPWR _22562_/X sky130_fd_sc_hd__mux4_1
X_34548_ _34612_/CLK _34548_/D VGND VGND VPWR VPWR _34548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24301_ _24301_/A VGND VGND VPWR VPWR _32682_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_221_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21513_ _21509_/X _21512_/X _21412_/X VGND VGND VPWR VPWR _21514_/D sky130_fd_sc_hd__o21ba_1
X_25281_ _25281_/A VGND VGND VPWR VPWR _33114_/D sky130_fd_sc_hd__clkbuf_1
X_22493_ _33097_/Q _32073_/Q _35849_/Q _35785_/Q _22384_/X _22385_/X VGND VGND VPWR
+ VPWR _22493_/X sky130_fd_sc_hd__mux4_1
XFILLER_37_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34479_ _36142_/CLK _34479_/D VGND VGND VPWR VPWR _34479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27020_ _27020_/A VGND VGND VPWR VPWR _33935_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36218_ _36223_/CLK _36218_/D VGND VGND VPWR VPWR _36218_/Q sky130_fd_sc_hd__dfxtp_1
X_24232_ _24232_/A VGND VGND VPWR VPWR _32651_/D sky130_fd_sc_hd__clkbuf_1
X_21444_ _21444_/A _21444_/B _21444_/C _21444_/D VGND VGND VPWR VPWR _21445_/A sky130_fd_sc_hd__or4_4
XFILLER_194_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36149_ _36149_/CLK _36149_/D VGND VGND VPWR VPWR _36149_/Q sky130_fd_sc_hd__dfxtp_1
X_24163_ _24163_/A VGND VGND VPWR VPWR _32618_/D sky130_fd_sc_hd__clkbuf_1
X_21375_ _22434_/A VGND VGND VPWR VPWR _21375_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_135_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23114_ _23114_/A VGND VGND VPWR VPWR _32096_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20326_ _35469_/Q _35405_/Q _35341_/Q _35277_/Q _20260_/X _20261_/X VGND VGND VPWR
+ VPWR _20326_/X sky130_fd_sc_hd__mux4_1
X_24094_ _24094_/A VGND VGND VPWR VPWR _32587_/D sky130_fd_sc_hd__clkbuf_1
X_28971_ _34796_/Q _27103_/X _28985_/S VGND VGND VPWR VPWR _28972_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_289_CLK clkbuf_6_58__f_CLK/X VGND VGND VPWR VPWR _36030_/CLK sky130_fd_sc_hd__clkbuf_16
X_23045_ _23045_/A VGND VGND VPWR VPWR _32072_/D sky130_fd_sc_hd__clkbuf_1
X_27922_ _27922_/A VGND VGND VPWR VPWR _34300_/D sky130_fd_sc_hd__clkbuf_1
X_20257_ _35723_/Q _32234_/Q _35595_/Q _35531_/Q _19970_/X _19971_/X VGND VGND VPWR
+ VPWR _20257_/X sky130_fd_sc_hd__mux4_1
XFILLER_118_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27853_ _27853_/A VGND VGND VPWR VPWR _34267_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20188_ _20184_/X _20187_/X _20146_/X _20147_/X VGND VGND VPWR VPWR _20203_/B sky130_fd_sc_hd__o211a_1
XTAP_5247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26804_ _33833_/Q _23289_/X _26804_/S VGND VGND VPWR VPWR _26805_/A sky130_fd_sc_hd__mux2_1
XTAP_5269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27784_ _27784_/A VGND VGND VPWR VPWR _34243_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24996_ _24996_/A VGND VGND VPWR VPWR _32981_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29523_ _29523_/A VGND VGND VPWR VPWR _35028_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26735_ _33800_/Q _23453_/X _26753_/S VGND VGND VPWR VPWR _26736_/A sky130_fd_sc_hd__mux2_1
XTAP_4568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_966 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23947_ _23947_/A VGND VGND VPWR VPWR _32518_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_461_CLK clkbuf_6_9__f_CLK/X VGND VGND VPWR VPWR _35434_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_72_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29454_ _29525_/S VGND VGND VPWR VPWR _29482_/S sky130_fd_sc_hd__buf_4
XTAP_3878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26666_ _26666_/A VGND VGND VPWR VPWR _33767_/D sky130_fd_sc_hd__clkbuf_1
X_23878_ _23878_/A VGND VGND VPWR VPWR _32485_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_233_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28405_ _27677_/X _34529_/Q _28421_/S VGND VGND VPWR VPWR _28406_/A sky130_fd_sc_hd__mux2_1
X_22829_ _32148_/Q _32340_/Q _32404_/Q _35924_/Q _22586_/X _21611_/A VGND VGND VPWR
+ VPWR _22829_/X sky130_fd_sc_hd__mux4_1
X_25617_ _24908_/X _33273_/Q _25625_/S VGND VGND VPWR VPWR _25618_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29385_ input10/X VGND VGND VPWR VPWR _29385_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_204_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26597_ _26597_/A VGND VGND VPWR VPWR _33736_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_213_CLK clkbuf_6_52__f_CLK/X VGND VGND VPWR VPWR _35661_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_164_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28336_ _28336_/A VGND VGND VPWR VPWR _34496_/D sky130_fd_sc_hd__clkbuf_1
X_16350_ _33886_/Q _33822_/Q _33758_/Q _36062_/Q _16318_/X _16319_/X VGND VGND VPWR
+ VPWR _16350_/X sky130_fd_sc_hd__mux4_1
XFILLER_44_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25548_ _24806_/X _33240_/Q _25562_/S VGND VGND VPWR VPWR _25549_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16281_ _16147_/X _16279_/X _16280_/X _16150_/X VGND VGND VPWR VPWR _16281_/X sky130_fd_sc_hd__a22o_1
XFILLER_12_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25479_ _25479_/A VGND VGND VPWR VPWR _33207_/D sky130_fd_sc_hd__clkbuf_1
X_28267_ _28378_/S VGND VGND VPWR VPWR _28286_/S sky130_fd_sc_hd__buf_6
XFILLER_139_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18020_ _32909_/Q _32845_/Q _32781_/Q _32717_/Q _17699_/X _17700_/X VGND VGND VPWR
+ VPWR _18020_/X sky130_fd_sc_hd__mux4_1
X_27218_ _34001_/Q _27217_/X _27218_/S VGND VGND VPWR VPWR _27219_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28198_ _27770_/X _34431_/Q _28214_/S VGND VGND VPWR VPWR _28199_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27149_ input31/X VGND VGND VPWR VPWR _27149_/X sky130_fd_sc_hd__buf_2
XFILLER_126_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30160_ _30160_/A VGND VGND VPWR VPWR _35329_/D sky130_fd_sc_hd__clkbuf_1
X_19971_ _20100_/A VGND VGND VPWR VPWR _19971_/X sky130_fd_sc_hd__buf_4
XFILLER_180_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18922_ _18747_/X _18920_/X _18921_/X _18750_/X VGND VGND VPWR VPWR _18922_/X sky130_fd_sc_hd__a22o_1
XFILLER_45_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30091_ _30091_/A VGND VGND VPWR VPWR _35296_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18853_ _18847_/X _18852_/X _18745_/X VGND VGND VPWR VPWR _18861_/C sky130_fd_sc_hd__o21ba_1
XTAP_6460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17804_ _33927_/Q _33863_/Q _33799_/Q _36103_/Q _17730_/X _17731_/X VGND VGND VPWR
+ VPWR _17804_/X sky130_fd_sc_hd__mux4_1
XFILLER_95_746 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33850_ _33850_/CLK _33850_/D VGND VGND VPWR VPWR _33850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18784_ _34657_/Q _34593_/Q _34529_/Q _34465_/Q _18533_/X _18534_/X VGND VGND VPWR
+ VPWR _18784_/X sky130_fd_sc_hd__mux4_1
XTAP_5770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15996_ _34134_/Q _34070_/Q _34006_/Q _33942_/Q _15993_/X _15995_/X VGND VGND VPWR
+ VPWR _15996_/X sky130_fd_sc_hd__mux4_1
XTAP_5781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32801_ _32804_/CLK _32801_/D VGND VGND VPWR VPWR _32801_/Q sky130_fd_sc_hd__dfxtp_1
X_17735_ _32645_/Q _32581_/Q _32517_/Q _35973_/Q _17629_/X _17413_/X VGND VGND VPWR
+ VPWR _17735_/X sky130_fd_sc_hd__mux4_1
X_33781_ _36085_/CLK _33781_/D VGND VGND VPWR VPWR _33781_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30993_ _30993_/A VGND VGND VPWR VPWR _35724_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35520_ _35648_/CLK _35520_/D VGND VGND VPWR VPWR _35520_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_452_CLK clkbuf_6_14__f_CLK/X VGND VGND VPWR VPWR _36142_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_224_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32732_ _36053_/CLK _32732_/D VGND VGND VPWR VPWR _32732_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_1162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17666_ _32131_/Q _32323_/Q _32387_/Q _35907_/Q _17633_/X _17421_/X VGND VGND VPWR
+ VPWR _17666_/X sky130_fd_sc_hd__mux4_1
XFILLER_165_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19405_ _32883_/Q _32819_/Q _32755_/Q _32691_/Q _19293_/X _19294_/X VGND VGND VPWR
+ VPWR _19405_/X sky130_fd_sc_hd__mux4_1
XFILLER_211_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16617_ _33061_/Q _32037_/Q _35813_/Q _35749_/Q _16372_/X _16373_/X VGND VGND VPWR
+ VPWR _16617_/X sky130_fd_sc_hd__mux4_1
X_35451_ _35451_/CLK _35451_/D VGND VGND VPWR VPWR _35451_/Q sky130_fd_sc_hd__dfxtp_1
X_32663_ _35863_/CLK _32663_/D VGND VGND VPWR VPWR _32663_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17597_ _32641_/Q _32577_/Q _32513_/Q _35969_/Q _17276_/X _17413_/X VGND VGND VPWR
+ VPWR _17597_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_204_CLK clkbuf_6_51__f_CLK/X VGND VGND VPWR VPWR _35721_/CLK sky130_fd_sc_hd__clkbuf_16
X_34402_ _36210_/CLK _34402_/D VGND VGND VPWR VPWR _34402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_245_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19336_ _35697_/Q _32205_/Q _35569_/Q _35505_/Q _19264_/X _19265_/X VGND VGND VPWR
+ VPWR _19336_/X sky130_fd_sc_hd__mux4_1
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31614_ _31614_/A VGND VGND VPWR VPWR _36018_/D sky130_fd_sc_hd__clkbuf_1
X_35382_ _35446_/CLK _35382_/D VGND VGND VPWR VPWR _35382_/Q sky130_fd_sc_hd__dfxtp_1
X_16548_ _17960_/A VGND VGND VPWR VPWR _16548_/X sky130_fd_sc_hd__buf_4
XFILLER_182_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32594_ _35986_/CLK _32594_/D VGND VGND VPWR VPWR _32594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34333_ _36060_/CLK _34333_/D VGND VGND VPWR VPWR _34333_/Q sky130_fd_sc_hd__dfxtp_1
X_31545_ _27828_/X _35986_/Q _31551_/S VGND VGND VPWR VPWR _31546_/A sky130_fd_sc_hd__mux2_1
X_19267_ _35631_/Q _34991_/Q _34351_/Q _33711_/Q _19091_/X _19092_/X VGND VGND VPWR
+ VPWR _19267_/X sky130_fd_sc_hd__mux4_1
XFILLER_91_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16479_ _16292_/X _16477_/X _16478_/X _16295_/X VGND VGND VPWR VPWR _16479_/X sky130_fd_sc_hd__a22o_1
X_18218_ _18218_/A VGND VGND VPWR VPWR _32019_/D sky130_fd_sc_hd__clkbuf_2
X_34264_ _34907_/CLK _34264_/D VGND VGND VPWR VPWR _34264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19198_ _35693_/Q _32201_/Q _35565_/Q _35501_/Q _18911_/X _18912_/X VGND VGND VPWR
+ VPWR _19198_/X sky130_fd_sc_hd__mux4_1
X_31476_ _27726_/X _35953_/Q _31480_/S VGND VGND VPWR VPWR _31477_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36003_ _36003_/CLK _36003_/D VGND VGND VPWR VPWR _36003_/Q sky130_fd_sc_hd__dfxtp_1
X_33215_ _36096_/CLK _33215_/D VGND VGND VPWR VPWR _33215_/Q sky130_fd_sc_hd__dfxtp_1
X_18149_ _18145_/X _18148_/X _17857_/X VGND VGND VPWR VPWR _18157_/C sky130_fd_sc_hd__o21ba_1
X_30427_ _35456_/Q _29460_/X _30441_/S VGND VGND VPWR VPWR _30428_/A sky130_fd_sc_hd__mux2_1
X_34195_ _34897_/CLK _34195_/D VGND VGND VPWR VPWR _34195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21160_ _21156_/X _21159_/X _21059_/X VGND VGND VPWR VPWR _21161_/D sky130_fd_sc_hd__o21ba_1
X_33146_ _36026_/CLK _33146_/D VGND VGND VPWR VPWR _33146_/Q sky130_fd_sc_hd__dfxtp_1
X_30358_ _30358_/A VGND VGND VPWR VPWR _35423_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20111_ _32903_/Q _32839_/Q _32775_/Q _32711_/Q _19999_/X _20000_/X VGND VGND VPWR
+ VPWR _20111_/X sky130_fd_sc_hd__mux4_1
XFILLER_176_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33077_ _35765_/CLK _33077_/D VGND VGND VPWR VPWR _33077_/Q sky130_fd_sc_hd__dfxtp_1
X_21091_ _21091_/A _21091_/B _21091_/C _21091_/D VGND VGND VPWR VPWR _21092_/A sky130_fd_sc_hd__or4_1
X_30289_ _30289_/A VGND VGND VPWR VPWR _35390_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_217_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20042_ _35717_/Q _32227_/Q _35589_/Q _35525_/Q _19970_/X _19971_/X VGND VGND VPWR
+ VPWR _20042_/X sky130_fd_sc_hd__mux4_1
X_32028_ _35998_/CLK _32028_/D VGND VGND VPWR VPWR _32028_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24850_ _24849_/X _32934_/Q _24859_/S VGND VGND VPWR VPWR _24851_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23801_ _23024_/X _32386_/Q _23811_/S VGND VGND VPWR VPWR _23802_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24781_ _24781_/A VGND VGND VPWR VPWR _32910_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33979_ _35449_/CLK _33979_/D VGND VGND VPWR VPWR _33979_/Q sky130_fd_sc_hd__dfxtp_1
X_21993_ _33083_/Q _32059_/Q _35835_/Q _35771_/Q _21678_/X _21679_/X VGND VGND VPWR
+ VPWR _21993_/X sky130_fd_sc_hd__mux4_1
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_443_CLK clkbuf_6_37__f_CLK/X VGND VGND VPWR VPWR _32879_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_54_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26520_ _24843_/X _33700_/Q _26530_/S VGND VGND VPWR VPWR _26521_/A sky130_fd_sc_hd__mux2_1
X_23732_ _22922_/X _32353_/Q _23748_/S VGND VGND VPWR VPWR _23733_/A sky130_fd_sc_hd__mux2_1
X_35718_ _35718_/CLK _35718_/D VGND VGND VPWR VPWR _35718_/Q sky130_fd_sc_hd__dfxtp_1
X_20944_ _20944_/A _20944_/B _20944_/C _20944_/D VGND VGND VPWR VPWR _20945_/A sky130_fd_sc_hd__or4_1
XFILLER_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26451_ _33668_/Q _23441_/X _26457_/S VGND VGND VPWR VPWR _26452_/A sky130_fd_sc_hd__mux2_1
X_23663_ _23024_/X _32322_/Q _23673_/S VGND VGND VPWR VPWR _23664_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35649_ _36099_/CLK _35649_/D VGND VGND VPWR VPWR _35649_/Q sky130_fd_sc_hd__dfxtp_1
X_20875_ _20875_/A VGND VGND VPWR VPWR _36187_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22614_ _22512_/X _22612_/X _22613_/X _22515_/X VGND VGND VPWR VPWR _22614_/X sky130_fd_sc_hd__a22o_1
XFILLER_198_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25402_ _25402_/A VGND VGND VPWR VPWR _33172_/D sky130_fd_sc_hd__clkbuf_1
X_29170_ _29170_/A VGND VGND VPWR VPWR _34890_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26382_ _33635_/Q _23271_/X _26394_/S VGND VGND VPWR VPWR _26383_/A sky130_fd_sc_hd__mux2_1
XFILLER_224_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23594_ _22922_/X _32289_/Q _23610_/S VGND VGND VPWR VPWR _23595_/A sky130_fd_sc_hd__mux2_1
X_28121_ _28121_/A VGND VGND VPWR VPWR _34394_/D sky130_fd_sc_hd__clkbuf_1
X_25333_ _25333_/A VGND VGND VPWR VPWR _33139_/D sky130_fd_sc_hd__clkbuf_1
X_22545_ _22505_/X _22543_/X _22544_/X _22510_/X VGND VGND VPWR VPWR _22545_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25264_ _25264_/A VGND VGND VPWR VPWR _33107_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28052_ _34362_/Q _27146_/X _28058_/S VGND VGND VPWR VPWR _28053_/A sky130_fd_sc_hd__mux2_1
X_22476_ _34185_/Q _34121_/Q _34057_/Q _33993_/Q _22399_/X _22400_/X VGND VGND VPWR
+ VPWR _22476_/X sky130_fd_sc_hd__mux4_1
XFILLER_155_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27003_ _27003_/A VGND VGND VPWR VPWR _33927_/D sky130_fd_sc_hd__clkbuf_1
X_24215_ _24215_/A VGND VGND VPWR VPWR _32643_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21427_ _32875_/Q _32811_/Q _32747_/Q _32683_/Q _21240_/X _21241_/X VGND VGND VPWR
+ VPWR _21427_/X sky130_fd_sc_hd__mux4_1
X_25195_ _25195_/A VGND VGND VPWR VPWR _33074_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24146_ _24146_/A VGND VGND VPWR VPWR _32610_/D sky130_fd_sc_hd__clkbuf_1
X_21358_ _35433_/Q _35369_/Q _35305_/Q _35241_/Q _21148_/X _21149_/X VGND VGND VPWR
+ VPWR _21358_/X sky130_fd_sc_hd__mux4_1
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20309_ _33677_/Q _33613_/Q _33549_/Q _33485_/Q _20206_/X _20207_/X VGND VGND VPWR
+ VPWR _20309_/X sky130_fd_sc_hd__mux4_1
XFILLER_162_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24077_ _24077_/A VGND VGND VPWR VPWR _32579_/D sky130_fd_sc_hd__clkbuf_1
X_28954_ _34788_/Q _27078_/X _28964_/S VGND VGND VPWR VPWR _28955_/A sky130_fd_sc_hd__mux2_1
X_21289_ _21285_/X _21288_/X _21045_/X VGND VGND VPWR VPWR _21297_/C sky130_fd_sc_hd__o21ba_1
XFILLER_150_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23028_ _23027_/X _32067_/Q _23040_/S VGND VGND VPWR VPWR _23029_/A sky130_fd_sc_hd__mux2_1
X_27905_ _27735_/X _34292_/Q _27923_/S VGND VGND VPWR VPWR _27906_/A sky130_fd_sc_hd__mux2_1
XTAP_5011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28885_ _28885_/A VGND VGND VPWR VPWR _34755_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27836_ _27836_/A VGND VGND VPWR VPWR _34260_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27767_ _27838_/S VGND VGND VPWR VPWR _27795_/S sky130_fd_sc_hd__buf_4
XTAP_4365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24979_ input54/X VGND VGND VPWR VPWR _24979_/X sky130_fd_sc_hd__buf_6
XTAP_4376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_434_CLK clkbuf_6_36__f_CLK/X VGND VGND VPWR VPWR _36146_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_79_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29506_ input53/X VGND VGND VPWR VPWR _29506_/X sky130_fd_sc_hd__clkbuf_4
XTAP_4387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17520_ _17520_/A _17520_/B _17520_/C _17520_/D VGND VGND VPWR VPWR _17521_/A sky130_fd_sc_hd__or4_1
XFILLER_45_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26718_ _33792_/Q _23429_/X _26732_/S VGND VGND VPWR VPWR _26719_/A sky130_fd_sc_hd__mux2_1
XTAP_4398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27698_ input10/X VGND VGND VPWR VPWR _27698_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17451_ _33917_/Q _33853_/Q _33789_/Q _36093_/Q _17377_/X _17378_/X VGND VGND VPWR
+ VPWR _17451_/X sky130_fd_sc_hd__mux4_1
X_29437_ _29437_/A VGND VGND VPWR VPWR _35000_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26649_ _26649_/A VGND VGND VPWR VPWR _33759_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16402_ _35679_/Q _32185_/Q _35551_/Q _35487_/Q _16258_/X _16259_/X VGND VGND VPWR
+ VPWR _16402_/X sky130_fd_sc_hd__mux4_1
XTAP_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29368_ _34978_/Q _29367_/X _29389_/S VGND VGND VPWR VPWR _29369_/A sky130_fd_sc_hd__mux2_1
X_17382_ _32635_/Q _32571_/Q _32507_/Q _35963_/Q _17276_/X _17060_/X VGND VGND VPWR
+ VPWR _17382_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19121_ _18800_/X _19119_/X _19120_/X _18803_/X VGND VGND VPWR VPWR _19121_/X sky130_fd_sc_hd__a22o_1
X_16333_ _35421_/Q _35357_/Q _35293_/Q _35229_/Q _16195_/X _16196_/X VGND VGND VPWR
+ VPWR _16333_/X sky130_fd_sc_hd__mux4_1
X_28319_ _28319_/A VGND VGND VPWR VPWR _34488_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29299_ _29326_/S VGND VGND VPWR VPWR _29318_/S sky130_fd_sc_hd__buf_4
XFILLER_199_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31330_ _31330_/A VGND VGND VPWR VPWR _35883_/D sky130_fd_sc_hd__clkbuf_1
X_19052_ _32873_/Q _32809_/Q _32745_/Q _32681_/Q _18940_/X _18941_/X VGND VGND VPWR
+ VPWR _19052_/X sky130_fd_sc_hd__mux4_1
X_16264_ _33051_/Q _32027_/Q _35803_/Q _35739_/Q _16067_/X _16069_/X VGND VGND VPWR
+ VPWR _16264_/X sky130_fd_sc_hd__mux4_1
XFILLER_158_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18003_ _34444_/Q _36172_/Q _34316_/Q _34252_/Q _17935_/X _17936_/X VGND VGND VPWR
+ VPWR _18003_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31261_ _27807_/X _35851_/Q _31273_/S VGND VGND VPWR VPWR _31262_/A sky130_fd_sc_hd__mux2_1
XFILLER_199_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16195_ _17850_/A VGND VGND VPWR VPWR _16195_/X sky130_fd_sc_hd__buf_6
XFILLER_86_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33000_ _35944_/CLK _33000_/D VGND VGND VPWR VPWR _33000_/Q sky130_fd_sc_hd__dfxtp_1
X_30212_ _35354_/Q _29342_/X _30222_/S VGND VGND VPWR VPWR _30213_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31192_ _27704_/X _35818_/Q _31210_/S VGND VGND VPWR VPWR _31193_/A sky130_fd_sc_hd__mux2_1
XFILLER_236_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19954_ _19954_/A _19954_/B _19954_/C _19954_/D VGND VGND VPWR VPWR _19955_/A sky130_fd_sc_hd__or4_4
X_30143_ _30143_/A VGND VGND VPWR VPWR _35321_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18905_ _33125_/Q _36005_/Q _32997_/Q _32933_/Q _18656_/X _18657_/X VGND VGND VPWR
+ VPWR _18905_/X sky130_fd_sc_hd__mux4_1
X_34951_ _36167_/CLK _34951_/D VGND VGND VPWR VPWR _34951_/Q sky130_fd_sc_hd__dfxtp_1
X_30074_ _30074_/A VGND VGND VPWR VPWR _35288_/D sky130_fd_sc_hd__clkbuf_1
X_19885_ _34944_/Q _34880_/Q _34816_/Q _34752_/Q _19813_/X _19814_/X VGND VGND VPWR
+ VPWR _19885_/X sky130_fd_sc_hd__mux4_1
XFILLER_136_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18836_ _18800_/X _18834_/X _18835_/X _18803_/X VGND VGND VPWR VPWR _18836_/X sky130_fd_sc_hd__a22o_1
X_33902_ _33902_/CLK _33902_/D VGND VGND VPWR VPWR _33902_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34882_ _36163_/CLK _34882_/D VGND VGND VPWR VPWR _34882_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1096 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33833_ _34153_/CLK _33833_/D VGND VGND VPWR VPWR _33833_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_6_43__f_CLK clkbuf_5_21_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_43__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_95_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18767_ _33889_/Q _33825_/Q _33761_/Q _36065_/Q _18618_/X _18619_/X VGND VGND VPWR
+ VPWR _18767_/X sky130_fd_sc_hd__mux4_1
X_15979_ input67/X input68/X VGND VGND VPWR VPWR _17765_/A sky130_fd_sc_hd__nor2b_4
XFILLER_110_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_212_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_425_CLK clkbuf_6_35__f_CLK/X VGND VGND VPWR VPWR _35828_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_82_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17718_ _35204_/Q _35140_/Q _35076_/Q _32260_/Q _17716_/X _17717_/X VGND VGND VPWR
+ VPWR _17718_/X sky130_fd_sc_hd__mux4_1
XFILLER_97_1443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_722 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33764_ _36070_/CLK _33764_/D VGND VGND VPWR VPWR _33764_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_1405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30976_ _30976_/A VGND VGND VPWR VPWR _35716_/D sky130_fd_sc_hd__clkbuf_1
X_18698_ _32095_/Q _32287_/Q _32351_/Q _35871_/Q _18521_/X _18662_/X VGND VGND VPWR
+ VPWR _18698_/X sky130_fd_sc_hd__mux4_1
XFILLER_82_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32715_ _32907_/CLK _32715_/D VGND VGND VPWR VPWR _32715_/Q sky130_fd_sc_hd__dfxtp_1
X_35503_ _35567_/CLK _35503_/D VGND VGND VPWR VPWR _35503_/Q sky130_fd_sc_hd__dfxtp_1
X_17649_ _17506_/X _17647_/X _17648_/X _17509_/X VGND VGND VPWR VPWR _17649_/X sky130_fd_sc_hd__a22o_1
XFILLER_91_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33695_ _35615_/CLK _33695_/D VGND VGND VPWR VPWR _33695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35434_ _35434_/CLK _35434_/D VGND VGND VPWR VPWR _35434_/Q sky130_fd_sc_hd__dfxtp_1
X_20660_ _22464_/A VGND VGND VPWR VPWR _20660_/X sky130_fd_sc_hd__buf_4
X_32646_ _35973_/CLK _32646_/D VGND VGND VPWR VPWR _32646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_991 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19319_ _19319_/A VGND VGND VPWR VPWR _32432_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35365_ _35365_/CLK _35365_/D VGND VGND VPWR VPWR _35365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20591_ _22510_/A VGND VGND VPWR VPWR _20591_/X sky130_fd_sc_hd__clkbuf_4
X_32577_ _35969_/CLK _32577_/D VGND VGND VPWR VPWR _32577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34316_ _36173_/CLK _34316_/D VGND VGND VPWR VPWR _34316_/Q sky130_fd_sc_hd__dfxtp_1
X_22330_ _22450_/A VGND VGND VPWR VPWR _22330_/X sky130_fd_sc_hd__buf_4
XFILLER_176_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31528_ _31528_/A VGND VGND VPWR VPWR _35977_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35296_ _36005_/CLK _35296_/D VGND VGND VPWR VPWR _35296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34247_ _34698_/CLK _34247_/D VGND VGND VPWR VPWR _34247_/Q sky130_fd_sc_hd__dfxtp_1
X_22261_ _22159_/X _22259_/X _22260_/X _22162_/X VGND VGND VPWR VPWR _22261_/X sky130_fd_sc_hd__a22o_1
X_31459_ _27701_/X _35945_/Q _31459_/S VGND VGND VPWR VPWR _31460_/A sky130_fd_sc_hd__mux2_1
X_24000_ _22915_/X _32543_/Q _24000_/S VGND VGND VPWR VPWR _24001_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21212_ _22400_/A VGND VGND VPWR VPWR _21212_/X sky130_fd_sc_hd__clkbuf_4
X_34178_ _34183_/CLK _34178_/D VGND VGND VPWR VPWR _34178_/Q sky130_fd_sc_hd__dfxtp_1
X_22192_ _22152_/X _22190_/X _22191_/X _22157_/X VGND VGND VPWR VPWR _22192_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21143_ _20961_/X _21141_/X _21142_/X _20965_/X VGND VGND VPWR VPWR _21143_/X sky130_fd_sc_hd__a22o_1
X_33129_ _36011_/CLK _33129_/D VGND VGND VPWR VPWR _33129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25951_ _24803_/X _33431_/Q _25967_/S VGND VGND VPWR VPWR _25952_/A sky130_fd_sc_hd__mux2_1
X_21074_ _32865_/Q _32801_/Q _32737_/Q _32673_/Q _20887_/X _20888_/X VGND VGND VPWR
+ VPWR _21074_/X sky130_fd_sc_hd__mux4_1
XFILLER_154_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20025_ _20025_/A VGND VGND VPWR VPWR _32452_/D sky130_fd_sc_hd__buf_2
X_24902_ input27/X VGND VGND VPWR VPWR _24902_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_63_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28670_ _28670_/A VGND VGND VPWR VPWR _34654_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_1294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25882_ _25882_/A VGND VGND VPWR VPWR _33398_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27621_ _34189_/Q _27205_/X _27629_/S VGND VGND VPWR VPWR _27622_/A sky130_fd_sc_hd__mux2_1
X_24833_ _24833_/A VGND VGND VPWR VPWR _32928_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_416_CLK clkbuf_6_32__f_CLK/X VGND VGND VPWR VPWR _35635_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_6_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27552_ _34156_/Q _27103_/X _27566_/S VGND VGND VPWR VPWR _27553_/A sky130_fd_sc_hd__mux2_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24764_ _24764_/A VGND VGND VPWR VPWR _32902_/D sky130_fd_sc_hd__clkbuf_1
X_21976_ _33403_/Q _33339_/Q _33275_/Q _33211_/Q _21727_/X _21728_/X VGND VGND VPWR
+ VPWR _21976_/X sky130_fd_sc_hd__mux4_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26503_ _24818_/X _33692_/Q _26509_/S VGND VGND VPWR VPWR _26504_/A sky130_fd_sc_hd__mux2_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23715_ _22897_/X _32345_/Q _23727_/S VGND VGND VPWR VPWR _23716_/A sky130_fd_sc_hd__mux2_1
X_20927_ _32861_/Q _32797_/Q _32733_/Q _32669_/Q _20887_/X _20888_/X VGND VGND VPWR
+ VPWR _20927_/X sky130_fd_sc_hd__mux4_1
XFILLER_25_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27483_ _27483_/A VGND VGND VPWR VPWR _34123_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24695_ _24695_/A VGND VGND VPWR VPWR _32869_/D sky130_fd_sc_hd__clkbuf_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_0_0_CLK clkbuf_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_7_0_CLK/A sky130_fd_sc_hd__clkbuf_8
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29222_ _34915_/Q _27075_/X _29234_/S VGND VGND VPWR VPWR _29223_/A sky130_fd_sc_hd__mux2_1
X_26434_ _33660_/Q _23414_/X _26436_/S VGND VGND VPWR VPWR _26435_/A sky130_fd_sc_hd__mux2_1
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20858_ _22399_/A VGND VGND VPWR VPWR _20858_/X sky130_fd_sc_hd__buf_6
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23646_ _22999_/X _32314_/Q _23652_/S VGND VGND VPWR VPWR _23647_/A sky130_fd_sc_hd__mux2_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29153_ _29153_/A VGND VGND VPWR VPWR _34882_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23577_ _22897_/X _32281_/Q _23589_/S VGND VGND VPWR VPWR _23578_/A sky130_fd_sc_hd__mux2_1
X_26365_ _33627_/Q _23246_/X _26373_/S VGND VGND VPWR VPWR _26366_/A sky130_fd_sc_hd__mux2_1
X_20789_ _32857_/Q _32793_/Q _32729_/Q _32665_/Q _20637_/X _20639_/X VGND VGND VPWR
+ VPWR _20789_/X sky130_fd_sc_hd__mux4_1
XFILLER_35_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28104_ _34387_/Q _27223_/X _28108_/S VGND VGND VPWR VPWR _28105_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22528_ _35466_/Q _35402_/Q _35338_/Q _35274_/Q _22207_/X _22208_/X VGND VGND VPWR
+ VPWR _22528_/X sky130_fd_sc_hd__mux4_1
X_25316_ _33131_/Q _23296_/X _25332_/S VGND VGND VPWR VPWR _25317_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26296_ _24914_/X _33595_/Q _26300_/S VGND VGND VPWR VPWR _26297_/A sky130_fd_sc_hd__mux2_1
X_29084_ _29084_/A VGND VGND VPWR VPWR _34849_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28035_ _34354_/Q _27121_/X _28037_/S VGND VGND VPWR VPWR _28036_/A sky130_fd_sc_hd__mux2_1
X_22459_ _22459_/A VGND VGND VPWR VPWR _22459_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_183_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25247_ _33099_/Q _23466_/X _25259_/S VGND VGND VPWR VPWR _25248_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25178_ _33066_/Q _23292_/X _25196_/S VGND VGND VPWR VPWR _25179_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24129_ _24129_/A VGND VGND VPWR VPWR _32602_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1074 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29986_ _35247_/Q _29407_/X _29994_/S VGND VGND VPWR VPWR _29987_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28937_ _34780_/Q _27053_/X _28943_/S VGND VGND VPWR VPWR _28938_/A sky130_fd_sc_hd__mux2_1
X_16951_ _34159_/Q _34095_/Q _34031_/Q _33967_/Q _16740_/X _16741_/X VGND VGND VPWR
+ VPWR _16951_/X sky130_fd_sc_hd__mux4_1
XFILLER_110_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19670_ _19666_/X _19669_/X _19465_/X VGND VGND VPWR VPWR _19671_/D sky130_fd_sc_hd__o21ba_1
X_28868_ _28868_/A VGND VGND VPWR VPWR _34747_/D sky130_fd_sc_hd__clkbuf_1
X_16882_ _16882_/A _16882_/B _16882_/C _16882_/D VGND VGND VPWR VPWR _16883_/A sky130_fd_sc_hd__or4_4
X_18621_ _18447_/X _18617_/X _18620_/X _18450_/X VGND VGND VPWR VPWR _18621_/X sky130_fd_sc_hd__a22o_1
XFILLER_49_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27819_ input53/X VGND VGND VPWR VPWR _27819_/X sky130_fd_sc_hd__clkbuf_4
XTAP_4151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28799_ _28799_/A VGND VGND VPWR VPWR _34714_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_407_CLK clkbuf_6_32__f_CLK/X VGND VGND VPWR VPWR _36082_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18552_ _33115_/Q _35995_/Q _32987_/Q _32923_/Q _18324_/X _18325_/X VGND VGND VPWR
+ VPWR _18552_/X sky130_fd_sc_hd__mux4_1
X_30830_ _35647_/Q input36/X _30846_/S VGND VGND VPWR VPWR _30831_/A sky130_fd_sc_hd__mux2_1
XTAP_4184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17503_ _17356_/X _17501_/X _17502_/X _17359_/X VGND VGND VPWR VPWR _17503_/X sky130_fd_sc_hd__a22o_1
XTAP_3472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18483_ _18447_/X _18481_/X _18482_/X _18450_/X VGND VGND VPWR VPWR _18483_/X sky130_fd_sc_hd__a22o_1
X_30761_ _30761_/A VGND VGND VPWR VPWR _35614_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1048 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32500_ _35956_/CLK _32500_/D VGND VGND VPWR VPWR _32500_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_233_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17434_ _17356_/X _17430_/X _17433_/X _17359_/X VGND VGND VPWR VPWR _17434_/X sky130_fd_sc_hd__a22o_1
X_33480_ _34121_/CLK _33480_/D VGND VGND VPWR VPWR _33480_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30692_ _30740_/S VGND VGND VPWR VPWR _30711_/S sky130_fd_sc_hd__buf_4
XFILLER_18_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32431_ _36072_/CLK _32431_/D VGND VGND VPWR VPWR _32431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17365_ _35194_/Q _35130_/Q _35066_/Q _32250_/Q _17363_/X _17364_/X VGND VGND VPWR
+ VPWR _17365_/X sky130_fd_sc_hd__mux4_1
XFILLER_242_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19104_ _19100_/X _19101_/X _19102_/X _19103_/X VGND VGND VPWR VPWR _19104_/X sky130_fd_sc_hd__a22o_1
X_35150_ _35731_/CLK _35150_/D VGND VGND VPWR VPWR _35150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16316_ _16140_/X _16314_/X _16315_/X _16145_/X VGND VGND VPWR VPWR _16316_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32362_ _35946_/CLK _32362_/D VGND VGND VPWR VPWR _32362_/Q sky130_fd_sc_hd__dfxtp_1
X_17296_ _17153_/X _17294_/X _17295_/X _17156_/X VGND VGND VPWR VPWR _17296_/X sky130_fd_sc_hd__a22o_1
XFILLER_105_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34101_ _34101_/CLK _34101_/D VGND VGND VPWR VPWR _34101_/Q sky130_fd_sc_hd__dfxtp_1
X_31313_ _31313_/A VGND VGND VPWR VPWR _35875_/D sky130_fd_sc_hd__clkbuf_1
X_19035_ _18752_/X _19033_/X _19034_/X _18757_/X VGND VGND VPWR VPWR _19035_/X sky130_fd_sc_hd__a22o_1
X_35081_ _35210_/CLK _35081_/D VGND VGND VPWR VPWR _35081_/Q sky130_fd_sc_hd__dfxtp_1
X_16247_ _33371_/Q _33307_/Q _33243_/Q _33179_/Q _16002_/X _16003_/X VGND VGND VPWR
+ VPWR _16247_/X sky130_fd_sc_hd__mux4_1
X_32293_ _35945_/CLK _32293_/D VGND VGND VPWR VPWR _32293_/Q sky130_fd_sc_hd__dfxtp_1
X_34032_ _35632_/CLK _34032_/D VGND VGND VPWR VPWR _34032_/Q sky130_fd_sc_hd__dfxtp_1
X_31244_ _27782_/X _35843_/Q _31252_/S VGND VGND VPWR VPWR _31245_/A sky130_fd_sc_hd__mux2_1
Xoutput104 _31980_/Q VGND VGND VPWR VPWR D1[22] sky130_fd_sc_hd__buf_2
X_16178_ _33625_/Q _33561_/Q _33497_/Q _33433_/Q _16141_/X _16142_/X VGND VGND VPWR
+ VPWR _16178_/X sky130_fd_sc_hd__mux4_1
XFILLER_142_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput115 _31990_/Q VGND VGND VPWR VPWR D1[32] sky130_fd_sc_hd__buf_2
XFILLER_99_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput126 _32000_/Q VGND VGND VPWR VPWR D1[42] sky130_fd_sc_hd__buf_2
XFILLER_47_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput137 _32010_/Q VGND VGND VPWR VPWR D1[52] sky130_fd_sc_hd__buf_2
Xoutput148 _32020_/Q VGND VGND VPWR VPWR D1[62] sky130_fd_sc_hd__buf_2
XFILLER_114_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput159 _36196_/Q VGND VGND VPWR VPWR D2[14] sky130_fd_sc_hd__buf_2
X_31175_ _27680_/X _35810_/Q _31189_/S VGND VGND VPWR VPWR _31176_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30126_ _30126_/A VGND VGND VPWR VPWR _35313_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_214_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19937_ _19932_/X _19936_/X _19793_/X _19794_/X VGND VGND VPWR VPWR _19954_/B sky130_fd_sc_hd__o211a_1
XFILLER_229_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35983_ _35983_/CLK _35983_/D VGND VGND VPWR VPWR _35983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30057_ _35281_/Q _29512_/X _30057_/S VGND VGND VPWR VPWR _30058_/A sky130_fd_sc_hd__mux2_1
X_19868_ _32128_/Q _32320_/Q _32384_/Q _35904_/Q _19580_/X _19721_/X VGND VGND VPWR
+ VPWR _19868_/X sky130_fd_sc_hd__mux4_1
XFILLER_25_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34934_ _36151_/CLK _34934_/D VGND VGND VPWR VPWR _34934_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_233_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18819_ _18815_/X _18818_/X _18745_/X VGND VGND VPWR VPWR _18829_/C sky130_fd_sc_hd__o21ba_1
X_19799_ _35646_/Q _35006_/Q _34366_/Q _33726_/Q _19797_/X _19798_/X VGND VGND VPWR
+ VPWR _19799_/X sky130_fd_sc_hd__mux4_1
XFILLER_23_1150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34865_ _35633_/CLK _34865_/D VGND VGND VPWR VPWR _34865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21830_ _22536_/A VGND VGND VPWR VPWR _21830_/X sky130_fd_sc_hd__buf_6
X_33816_ _36057_/CLK _33816_/D VGND VGND VPWR VPWR _33816_/Q sky130_fd_sc_hd__dfxtp_1
X_34796_ _34924_/CLK _34796_/D VGND VGND VPWR VPWR _34796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33747_ _35026_/CLK _33747_/D VGND VGND VPWR VPWR _33747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21761_ _21761_/A VGND VGND VPWR VPWR _21761_/X sky130_fd_sc_hd__buf_4
XFILLER_51_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30959_ _30959_/A VGND VGND VPWR VPWR _35708_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_212_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23500_ _23500_/A VGND VGND VPWR VPWR _32245_/D sky130_fd_sc_hd__clkbuf_1
X_20712_ _22450_/A VGND VGND VPWR VPWR _20712_/X sky130_fd_sc_hd__buf_6
XFILLER_52_966 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24480_ _24480_/A VGND VGND VPWR VPWR _32767_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33678_ _33934_/CLK _33678_/D VGND VGND VPWR VPWR _33678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21692_ _33651_/Q _33587_/Q _33523_/Q _33459_/Q _21447_/X _21448_/X VGND VGND VPWR
+ VPWR _21692_/X sky130_fd_sc_hd__mux4_1
XFILLER_11_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23431_ _23431_/A VGND VGND VPWR VPWR _32222_/D sky130_fd_sc_hd__clkbuf_1
X_35417_ _35801_/CLK _35417_/D VGND VGND VPWR VPWR _35417_/Q sky130_fd_sc_hd__dfxtp_1
X_20643_ input75/X VGND VGND VPWR VPWR _22446_/A sky130_fd_sc_hd__buf_6
X_32629_ _34485_/CLK _32629_/D VGND VGND VPWR VPWR _32629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26150_ _26150_/A VGND VGND VPWR VPWR _33525_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35348_ _35860_/CLK _35348_/D VGND VGND VPWR VPWR _35348_/Q sky130_fd_sc_hd__dfxtp_1
X_23362_ _32197_/Q _23292_/X _23385_/S VGND VGND VPWR VPWR _23363_/A sky130_fd_sc_hd__mux2_1
X_20574_ _34965_/Q _34901_/Q _34837_/Q _34773_/Q _18383_/X _18385_/X VGND VGND VPWR
+ VPWR _20574_/X sky130_fd_sc_hd__mux4_1
XFILLER_108_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22313_ _22309_/X _22310_/X _22311_/X _22312_/X VGND VGND VPWR VPWR _22313_/X sky130_fd_sc_hd__a22o_1
X_25101_ _24951_/X _33031_/Q _25101_/S VGND VGND VPWR VPWR _25102_/A sky130_fd_sc_hd__mux2_1
X_26081_ _26081_/A VGND VGND VPWR VPWR _33493_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_176_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35279_ _35599_/CLK _35279_/D VGND VGND VPWR VPWR _35279_/Q sky130_fd_sc_hd__dfxtp_1
X_23293_ _23565_/S VGND VGND VPWR VPWR _23424_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_194_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25032_ _24849_/X _32998_/Q _25038_/S VGND VGND VPWR VPWR _25033_/A sky130_fd_sc_hd__mux2_1
X_22244_ _22240_/X _22243_/X _22104_/X VGND VGND VPWR VPWR _22254_/C sky130_fd_sc_hd__o21ba_1
XFILLER_152_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29840_ _29930_/S VGND VGND VPWR VPWR _29859_/S sky130_fd_sc_hd__clkbuf_8
X_22175_ _35456_/Q _35392_/Q _35328_/Q _35264_/Q _21854_/X _21855_/X VGND VGND VPWR
+ VPWR _22175_/X sky130_fd_sc_hd__mux4_1
XFILLER_195_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21126_ _34914_/Q _34850_/Q _34786_/Q _34722_/Q _21054_/X _21055_/X VGND VGND VPWR
+ VPWR _21126_/X sky130_fd_sc_hd__mux4_1
X_29771_ _35145_/Q _29488_/X _29787_/S VGND VGND VPWR VPWR _29772_/A sky130_fd_sc_hd__mux2_1
XFILLER_132_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26983_ _27031_/S VGND VGND VPWR VPWR _27002_/S sky130_fd_sc_hd__buf_6
XFILLER_8_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28722_ _34679_/Q _27137_/X _28734_/S VGND VGND VPWR VPWR _28723_/A sky130_fd_sc_hd__mux2_1
X_25934_ _25934_/A VGND VGND VPWR VPWR _33423_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_1244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21057_ _21763_/A VGND VGND VPWR VPWR _21057_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_87_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20008_ _20004_/X _20005_/X _20006_/X _20007_/X VGND VGND VPWR VPWR _20008_/X sky130_fd_sc_hd__a22o_1
XFILLER_47_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28653_ _34646_/Q _27033_/X _28671_/S VGND VGND VPWR VPWR _28654_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_1015 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25865_ _25865_/A VGND VGND VPWR VPWR _33390_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27604_ _34181_/Q _27180_/X _27608_/S VGND VGND VPWR VPWR _27605_/A sky130_fd_sc_hd__mux2_1
X_24816_ _24815_/X _32923_/Q _24828_/S VGND VGND VPWR VPWR _24817_/A sky130_fd_sc_hd__mux2_1
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28584_ _27742_/X _34614_/Q _28598_/S VGND VGND VPWR VPWR _28585_/A sky130_fd_sc_hd__mux2_1
X_25796_ _24973_/X _33358_/Q _25802_/S VGND VGND VPWR VPWR _25797_/A sky130_fd_sc_hd__mux2_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27535_ _34148_/Q _27078_/X _27545_/S VGND VGND VPWR VPWR _27536_/A sky130_fd_sc_hd__mux2_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24747_ _23011_/X _32894_/Q _24765_/S VGND VGND VPWR VPWR _24748_/A sky130_fd_sc_hd__mux2_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21959_ _22469_/A VGND VGND VPWR VPWR _21959_/X sky130_fd_sc_hd__buf_4
XFILLER_128_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27466_ _27466_/A VGND VGND VPWR VPWR _34115_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24678_ _24678_/A VGND VGND VPWR VPWR _32861_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29205_ _34907_/Q _27050_/X _29213_/S VGND VGND VPWR VPWR _29206_/A sky130_fd_sc_hd__mux2_1
X_26417_ _26486_/S VGND VGND VPWR VPWR _26436_/S sky130_fd_sc_hd__buf_4
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23629_ _22974_/X _32306_/Q _23631_/S VGND VGND VPWR VPWR _23630_/A sky130_fd_sc_hd__mux2_1
X_27397_ _27397_/A VGND VGND VPWR VPWR _34082_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17150_ _17003_/X _17148_/X _17149_/X _17006_/X VGND VGND VPWR VPWR _17150_/X sky130_fd_sc_hd__a22o_1
X_29136_ _29136_/A VGND VGND VPWR VPWR _34874_/D sky130_fd_sc_hd__clkbuf_1
X_26348_ _24991_/X _33620_/Q _26350_/S VGND VGND VPWR VPWR _26349_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput17 DW[24] VGND VGND VPWR VPWR input17/X sky130_fd_sc_hd__buf_4
X_16101_ _17163_/A VGND VGND VPWR VPWR _16101_/X sky130_fd_sc_hd__clkbuf_4
Xinput28 DW[34] VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__clkbuf_4
XFILLER_13_1330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput39 DW[44] VGND VGND VPWR VPWR input39/X sky130_fd_sc_hd__buf_6
X_29067_ _29067_/A VGND VGND VPWR VPWR _34841_/D sky130_fd_sc_hd__clkbuf_1
X_17081_ _17003_/X _17077_/X _17080_/X _17006_/X VGND VGND VPWR VPWR _17081_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_6_7__f_CLK clkbuf_5_3_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_7__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_26279_ _24889_/X _33587_/Q _26279_/S VGND VGND VPWR VPWR _26280_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16032_ _17986_/A VGND VGND VPWR VPWR _16032_/X sky130_fd_sc_hd__buf_6
X_28018_ _28108_/S VGND VGND VPWR VPWR _28037_/S sky130_fd_sc_hd__buf_4
XFILLER_143_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17983_ _32652_/Q _32588_/Q _32524_/Q _35980_/Q _17982_/X _17766_/X VGND VGND VPWR
+ VPWR _17983_/X sky130_fd_sc_hd__mux4_1
XFILLER_2_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29969_ _35239_/Q _29382_/X _29973_/S VGND VGND VPWR VPWR _29970_/A sky130_fd_sc_hd__mux2_1
X_19722_ _32124_/Q _32316_/Q _32380_/Q _35900_/Q _19580_/X _19721_/X VGND VGND VPWR
+ VPWR _19722_/X sky130_fd_sc_hd__mux4_1
X_16934_ _16645_/X _16932_/X _16933_/X _16648_/X VGND VGND VPWR VPWR _16934_/X sky130_fd_sc_hd__a22o_1
X_32980_ _36052_/CLK _32980_/D VGND VGND VPWR VPWR _32980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31931_ _31931_/A VGND VGND VPWR VPWR _36168_/D sky130_fd_sc_hd__clkbuf_1
X_19653_ _35642_/Q _35002_/Q _34362_/Q _33722_/Q _19444_/X _19445_/X VGND VGND VPWR
+ VPWR _19653_/X sky130_fd_sc_hd__mux4_1
XFILLER_133_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16865_ _16861_/X _16864_/X _16787_/X _16788_/X VGND VGND VPWR VPWR _16882_/B sky130_fd_sc_hd__o211a_1
XFILLER_65_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18604_ _20016_/A VGND VGND VPWR VPWR _18604_/X sky130_fd_sc_hd__buf_6
X_34650_ _36125_/CLK _34650_/D VGND VGND VPWR VPWR _34650_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31862_ _23286_/X _36136_/Q _31864_/S VGND VGND VPWR VPWR _31863_/A sky130_fd_sc_hd__mux2_1
X_19584_ _19579_/X _19583_/X _19440_/X _19441_/X VGND VGND VPWR VPWR _19601_/B sky130_fd_sc_hd__o211a_1
X_16796_ _33066_/Q _32042_/Q _35818_/Q _35754_/Q _16725_/X _16726_/X VGND VGND VPWR
+ VPWR _16796_/X sky130_fd_sc_hd__mux4_1
X_33601_ _34180_/CLK _33601_/D VGND VGND VPWR VPWR _33601_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18535_ _34650_/Q _34586_/Q _34522_/Q _34458_/Q _18533_/X _18534_/X VGND VGND VPWR
+ VPWR _18535_/X sky130_fd_sc_hd__mux4_1
X_30813_ _35639_/Q input27/X _30825_/S VGND VGND VPWR VPWR _30814_/A sky130_fd_sc_hd__mux2_1
X_34581_ _34708_/CLK _34581_/D VGND VGND VPWR VPWR _34581_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31793_ _31793_/A VGND VGND VPWR VPWR _36103_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_179_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_916 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33532_ _36093_/CLK _33532_/D VGND VGND VPWR VPWR _33532_/Q sky130_fd_sc_hd__dfxtp_1
X_18466_ _18462_/X _18465_/X _18375_/X VGND VGND VPWR VPWR _18476_/C sky130_fd_sc_hd__o21ba_1
X_30744_ _35606_/Q input1/X _30762_/S VGND VGND VPWR VPWR _30745_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17417_ _33148_/Q _36028_/Q _33020_/Q _32956_/Q _17415_/X _17416_/X VGND VGND VPWR
+ VPWR _17417_/X sky130_fd_sc_hd__mux4_1
XFILLER_222_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33463_ _33911_/CLK _33463_/D VGND VGND VPWR VPWR _33463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_1170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18397_ _20074_/A VGND VGND VPWR VPWR _19461_/A sky130_fd_sc_hd__buf_12
X_30675_ _30675_/A VGND VGND VPWR VPWR _35573_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_222_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35202_ _35715_/CLK _35202_/D VGND VGND VPWR VPWR _35202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32414_ _33573_/CLK _32414_/D VGND VGND VPWR VPWR _32414_/Q sky130_fd_sc_hd__dfxtp_1
X_36182_ _36191_/CLK _36182_/D VGND VGND VPWR VPWR _36182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17348_ _32890_/Q _32826_/Q _32762_/Q _32698_/Q _17346_/X _17347_/X VGND VGND VPWR
+ VPWR _17348_/X sky130_fd_sc_hd__mux4_1
X_33394_ _36082_/CLK _33394_/D VGND VGND VPWR VPWR _33394_/Q sky130_fd_sc_hd__dfxtp_1
X_35133_ _35577_/CLK _35133_/D VGND VGND VPWR VPWR _35133_/Q sky130_fd_sc_hd__dfxtp_1
X_32345_ _35865_/CLK _32345_/D VGND VGND VPWR VPWR _32345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17279_ _17059_/X _17277_/X _17278_/X _17065_/X VGND VGND VPWR VPWR _17279_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19018_ _20215_/A VGND VGND VPWR VPWR _19018_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_106_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35064_ _36150_/CLK _35064_/D VGND VGND VPWR VPWR _35064_/Q sky130_fd_sc_hd__dfxtp_1
X_32276_ _35221_/CLK _32276_/D VGND VGND VPWR VPWR _32276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20290_ _20285_/X _20289_/X _20146_/X _20147_/X VGND VGND VPWR VPWR _20307_/B sky130_fd_sc_hd__o211a_1
XFILLER_161_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34015_ _36188_/CLK _34015_/D VGND VGND VPWR VPWR _34015_/Q sky130_fd_sc_hd__dfxtp_1
X_31227_ _27757_/X _35835_/Q _31231_/S VGND VGND VPWR VPWR _31228_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31158_ _27655_/X _35802_/Q _31168_/S VGND VGND VPWR VPWR _31159_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30109_ _30109_/A VGND VGND VPWR VPWR _35305_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23980_ _31418_/A _31553_/A VGND VGND VPWR VPWR _24113_/S sky130_fd_sc_hd__nand2_8
X_35966_ _36031_/CLK _35966_/D VGND VGND VPWR VPWR _35966_/Q sky130_fd_sc_hd__dfxtp_1
X_31089_ _35770_/Q input30/X _31095_/S VGND VGND VPWR VPWR _31090_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34917_ _34920_/CLK _34917_/D VGND VGND VPWR VPWR _34917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_1158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22931_ input6/X VGND VGND VPWR VPWR _22931_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_96_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_244_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35897_ _35961_/CLK _35897_/D VGND VGND VPWR VPWR _35897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_243_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25650_ _25650_/A VGND VGND VPWR VPWR _33288_/D sky130_fd_sc_hd__clkbuf_1
X_22862_ _22858_/X _22861_/X _22446_/A _22447_/A VGND VGND VPWR VPWR _22877_/B sky130_fd_sc_hd__o211a_1
X_34848_ _34915_/CLK _34848_/D VGND VGND VPWR VPWR _34848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24601_ _22996_/X _32825_/Q _24609_/S VGND VGND VPWR VPWR _24602_/A sky130_fd_sc_hd__mux2_1
X_21813_ _33142_/Q _36022_/Q _33014_/Q _32950_/Q _21662_/X _21663_/X VGND VGND VPWR
+ VPWR _21813_/X sky130_fd_sc_hd__mux4_1
X_22793_ _33939_/Q _33875_/Q _33811_/Q _36115_/Q _20662_/X _20664_/X VGND VGND VPWR
+ VPWR _22793_/X sky130_fd_sc_hd__mux4_1
X_25581_ _24855_/X _33256_/Q _25583_/S VGND VGND VPWR VPWR _25582_/A sky130_fd_sc_hd__mux2_1
X_34779_ _36121_/CLK _34779_/D VGND VGND VPWR VPWR _34779_/Q sky130_fd_sc_hd__dfxtp_1
X_27320_ _34046_/Q _27158_/X _27338_/S VGND VGND VPWR VPWR _27321_/A sky130_fd_sc_hd__mux2_1
X_24532_ _22894_/X _32792_/Q _24546_/S VGND VGND VPWR VPWR _24533_/A sky130_fd_sc_hd__mux2_1
XPHY_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21744_ _22598_/A VGND VGND VPWR VPWR _21744_/X sky130_fd_sc_hd__buf_6
XPHY_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27251_ _27251_/A VGND VGND VPWR VPWR _34013_/D sky130_fd_sc_hd__clkbuf_1
X_21675_ _35634_/Q _34994_/Q _34354_/Q _33714_/Q _21391_/X _21392_/X VGND VGND VPWR
+ VPWR _21675_/X sky130_fd_sc_hd__mux4_1
X_24463_ _24463_/A VGND VGND VPWR VPWR _32759_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_237_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26202_ _26202_/A VGND VGND VPWR VPWR _33550_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_225_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20626_ _33110_/Q _35990_/Q _32982_/Q _32918_/Q _20624_/X _20625_/X VGND VGND VPWR
+ VPWR _20626_/X sky130_fd_sc_hd__mux4_1
XFILLER_32_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23414_ input32/X VGND VGND VPWR VPWR _23414_/X sky130_fd_sc_hd__buf_4
X_27182_ _27182_/A VGND VGND VPWR VPWR _33989_/D sky130_fd_sc_hd__clkbuf_1
X_24394_ _24394_/A VGND VGND VPWR VPWR _32726_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26133_ _26133_/A VGND VGND VPWR VPWR _33517_/D sky130_fd_sc_hd__clkbuf_1
X_23345_ _32189_/Q _23268_/X _23359_/S VGND VGND VPWR VPWR _23346_/A sky130_fd_sc_hd__mux2_1
X_20557_ _33173_/Q _36053_/Q _33045_/Q _32981_/Q _18332_/X _19461_/A VGND VGND VPWR
+ VPWR _20557_/X sky130_fd_sc_hd__mux4_1
XFILLER_123_1377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26064_ _24970_/X _33485_/Q _26072_/S VGND VGND VPWR VPWR _26065_/A sky130_fd_sc_hd__mux2_1
X_23276_ _23276_/A VGND VGND VPWR VPWR _32164_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20488_ _20488_/A VGND VGND VPWR VPWR _32466_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_164_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22227_ _22159_/X _22225_/X _22226_/X _22162_/X VGND VGND VPWR VPWR _22227_/X sky130_fd_sc_hd__a22o_1
X_25015_ _24824_/X _32990_/Q _25017_/S VGND VGND VPWR VPWR _25016_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29823_ _29823_/A VGND VGND VPWR VPWR _35169_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22158_ _22152_/X _22155_/X _22156_/X _22157_/X VGND VGND VPWR VPWR _22158_/X sky130_fd_sc_hd__a22o_1
XTAP_6834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21109_ _32098_/Q _32290_/Q _32354_/Q _35874_/Q _20821_/X _20962_/X VGND VGND VPWR
+ VPWR _21109_/X sky130_fd_sc_hd__mux4_1
XTAP_6867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29754_ _35137_/Q _29463_/X _29766_/S VGND VGND VPWR VPWR _29755_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22089_ _22012_/X _22087_/X _22088_/X _22018_/X VGND VGND VPWR VPWR _22089_/X sky130_fd_sc_hd__a22o_1
X_26966_ _26966_/A VGND VGND VPWR VPWR _33909_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28705_ _34671_/Q _27112_/X _28713_/S VGND VGND VPWR VPWR _28706_/A sky130_fd_sc_hd__mux2_1
X_25917_ _25917_/A VGND VGND VPWR VPWR _33415_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29685_ _35104_/Q _29360_/X _29703_/S VGND VGND VPWR VPWR _29686_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26897_ _26897_/A VGND VGND VPWR VPWR _33877_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28636_ _27819_/X _34639_/Q _28640_/S VGND VGND VPWR VPWR _28637_/A sky130_fd_sc_hd__mux2_1
X_16650_ _17864_/A VGND VGND VPWR VPWR _16650_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_78_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25848_ _25848_/A VGND VGND VPWR VPWR _33382_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28567_ _27717_/X _34606_/Q _28577_/S VGND VGND VPWR VPWR _28568_/A sky130_fd_sc_hd__mux2_1
X_16581_ _16292_/X _16579_/X _16580_/X _16295_/X VGND VGND VPWR VPWR _16581_/X sky130_fd_sc_hd__a22o_1
X_25779_ _24948_/X _33350_/Q _25781_/S VGND VGND VPWR VPWR _25780_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18320_ _20282_/A VGND VGND VPWR VPWR _20166_/A sky130_fd_sc_hd__buf_12
X_27518_ _34140_/Q _27053_/X _27524_/S VGND VGND VPWR VPWR _27519_/A sky130_fd_sc_hd__mux2_1
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28498_ _28498_/A VGND VGND VPWR VPWR _34573_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18251_ _16018_/X _18249_/X _18250_/X _16027_/X VGND VGND VPWR VPWR _18251_/X sky130_fd_sc_hd__a22o_1
XFILLER_188_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27449_ _27449_/A VGND VGND VPWR VPWR _34107_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_230_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17202_ _33654_/Q _33590_/Q _33526_/Q _33462_/Q _17200_/X _17201_/X VGND VGND VPWR
+ VPWR _17202_/X sky130_fd_sc_hd__mux4_1
X_18182_ _16048_/X _18180_/X _18181_/X _16058_/X VGND VGND VPWR VPWR _18182_/X sky130_fd_sc_hd__a22o_1
X_30460_ _35472_/Q _29509_/X _30462_/S VGND VGND VPWR VPWR _30461_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_857 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17133_ _17126_/X _17131_/X _17132_/X VGND VGND VPWR VPWR _17167_/A sky130_fd_sc_hd__o21ba_1
X_29119_ _29119_/A VGND VGND VPWR VPWR _34866_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30391_ _35439_/Q _29407_/X _30399_/S VGND VGND VPWR VPWR _30392_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32130_ _35970_/CLK _32130_/D VGND VGND VPWR VPWR _32130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17064_ _33138_/Q _36018_/Q _33010_/Q _32946_/Q _17062_/X _17063_/X VGND VGND VPWR
+ VPWR _17064_/X sky130_fd_sc_hd__mux4_1
XFILLER_195_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16015_ _17838_/A VGND VGND VPWR VPWR _16015_/X sky130_fd_sc_hd__buf_4
X_32061_ _35453_/CLK _32061_/D VGND VGND VPWR VPWR _32061_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_1362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31012_ _31147_/A _31688_/A VGND VGND VPWR VPWR _31145_/S sky130_fd_sc_hd__nor2_8
XFILLER_112_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35820_ _35820_/CLK _35820_/D VGND VGND VPWR VPWR _35820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_215_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17966_ _34699_/Q _34635_/Q _34571_/Q _34507_/Q _17645_/X _17646_/X VGND VGND VPWR
+ VPWR _17966_/X sky130_fd_sc_hd__mux4_1
XFILLER_215_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16917_ _34158_/Q _34094_/Q _34030_/Q _33966_/Q _16740_/X _16741_/X VGND VGND VPWR
+ VPWR _16917_/X sky130_fd_sc_hd__mux4_1
X_19705_ _33660_/Q _33596_/Q _33532_/Q _33468_/Q _19500_/X _19501_/X VGND VGND VPWR
+ VPWR _19705_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32963_ _35779_/CLK _32963_/D VGND VGND VPWR VPWR _32963_/Q sky130_fd_sc_hd__dfxtp_1
X_35751_ _35814_/CLK _35751_/D VGND VGND VPWR VPWR _35751_/Q sky130_fd_sc_hd__dfxtp_1
X_17897_ _35209_/Q _35145_/Q _35081_/Q _32265_/Q _17716_/X _17717_/X VGND VGND VPWR
+ VPWR _17897_/X sky130_fd_sc_hd__mux4_1
XFILLER_22_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34702_ _35664_/CLK _34702_/D VGND VGND VPWR VPWR _34702_/Q sky130_fd_sc_hd__dfxtp_1
X_31914_ _31914_/A VGND VGND VPWR VPWR _36160_/D sky130_fd_sc_hd__clkbuf_1
X_19636_ _34170_/Q _34106_/Q _34042_/Q _33978_/Q _19393_/X _19394_/X VGND VGND VPWR
+ VPWR _19636_/X sky130_fd_sc_hd__mux4_1
X_16848_ _17907_/A VGND VGND VPWR VPWR _16848_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_65_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32894_ _32894_/CLK _32894_/D VGND VGND VPWR VPWR _32894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35682_ _36135_/CLK _35682_/D VGND VGND VPWR VPWR _35682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34633_ _34633_/CLK _34633_/D VGND VGND VPWR VPWR _34633_/Q sky130_fd_sc_hd__dfxtp_1
X_31845_ _31956_/S VGND VGND VPWR VPWR _31864_/S sky130_fd_sc_hd__buf_4
X_19567_ _19567_/A _19567_/B _19567_/C _19567_/D VGND VGND VPWR VPWR _19568_/A sky130_fd_sc_hd__or4_1
XFILLER_92_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16779_ _17838_/A VGND VGND VPWR VPWR _16779_/X sky130_fd_sc_hd__buf_2
XFILLER_81_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18518_ _32602_/Q _32538_/Q _32474_/Q _35930_/Q _18517_/X _20017_/A VGND VGND VPWR
+ VPWR _18518_/X sky130_fd_sc_hd__mux4_1
XFILLER_230_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34564_ _34693_/CLK _34564_/D VGND VGND VPWR VPWR _34564_/Q sky130_fd_sc_hd__dfxtp_1
X_31776_ _36095_/Q input36/X _31792_/S VGND VGND VPWR VPWR _31777_/A sky130_fd_sc_hd__mux2_1
X_19498_ _19498_/A VGND VGND VPWR VPWR _32437_/D sky130_fd_sc_hd__buf_2
XFILLER_59_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30727_ _30727_/A VGND VGND VPWR VPWR _35598_/D sky130_fd_sc_hd__clkbuf_1
X_18449_ _33880_/Q _33816_/Q _33752_/Q _36056_/Q _18412_/X _18413_/X VGND VGND VPWR
+ VPWR _18449_/X sky130_fd_sc_hd__mux4_1
X_33515_ _33895_/CLK _33515_/D VGND VGND VPWR VPWR _33515_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34495_ _35071_/CLK _34495_/D VGND VGND VPWR VPWR _34495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36234_ _36235_/CLK _36234_/D VGND VGND VPWR VPWR _36234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33446_ _34146_/CLK _33446_/D VGND VGND VPWR VPWR _33446_/Q sky130_fd_sc_hd__dfxtp_1
X_21460_ _33132_/Q _36012_/Q _33004_/Q _32940_/Q _21309_/X _21310_/X VGND VGND VPWR
+ VPWR _21460_/X sky130_fd_sc_hd__mux4_1
XFILLER_222_1243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30658_ _30658_/A VGND VGND VPWR VPWR _35565_/D sky130_fd_sc_hd__clkbuf_1
X_20411_ _19458_/A _20409_/X _20410_/X _19463_/A VGND VGND VPWR VPWR _20411_/X sky130_fd_sc_hd__a22o_1
X_36165_ _36165_/CLK _36165_/D VGND VGND VPWR VPWR _36165_/Q sky130_fd_sc_hd__dfxtp_1
X_33377_ _36066_/CLK _33377_/D VGND VGND VPWR VPWR _33377_/Q sky130_fd_sc_hd__dfxtp_1
X_21391_ _22598_/A VGND VGND VPWR VPWR _21391_/X sky130_fd_sc_hd__buf_6
X_30589_ _35533_/Q _29500_/X _30597_/S VGND VGND VPWR VPWR _30590_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23130_ _23130_/A VGND VGND VPWR VPWR _32104_/D sky130_fd_sc_hd__clkbuf_1
X_20342_ _33422_/Q _33358_/Q _33294_/Q _33230_/Q _20133_/X _20134_/X VGND VGND VPWR
+ VPWR _20342_/X sky130_fd_sc_hd__mux4_1
X_32328_ _35976_/CLK _32328_/D VGND VGND VPWR VPWR _32328_/Q sky130_fd_sc_hd__dfxtp_1
X_35116_ _35564_/CLK _35116_/D VGND VGND VPWR VPWR _35116_/Q sky130_fd_sc_hd__dfxtp_1
X_36096_ _36096_/CLK _36096_/D VGND VGND VPWR VPWR _36096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23061_ input52/X VGND VGND VPWR VPWR _23061_/X sky130_fd_sc_hd__buf_2
X_35047_ _35367_/CLK _35047_/D VGND VGND VPWR VPWR _35047_/Q sky130_fd_sc_hd__dfxtp_1
X_32259_ _34691_/CLK _32259_/D VGND VGND VPWR VPWR _32259_/Q sky130_fd_sc_hd__dfxtp_1
X_20273_ _20273_/A _20273_/B _20273_/C _20273_/D VGND VGND VPWR VPWR _20274_/A sky130_fd_sc_hd__or4_1
XTAP_6108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22012_ _22505_/A VGND VGND VPWR VPWR _22012_/X sky130_fd_sc_hd__clkbuf_4
XTAP_6119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26820_ _26820_/A VGND VGND VPWR VPWR _33840_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1069 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26751_ _33808_/Q _23481_/X _26753_/S VGND VGND VPWR VPWR _26752_/A sky130_fd_sc_hd__mux2_1
XTAP_4728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23963_ _23061_/X _32526_/Q _23969_/S VGND VGND VPWR VPWR _23964_/A sky130_fd_sc_hd__mux2_1
X_35949_ _35949_/CLK _35949_/D VGND VGND VPWR VPWR _35949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25702_ _24834_/X _33313_/Q _25718_/S VGND VGND VPWR VPWR _25703_/A sky130_fd_sc_hd__mux2_1
XFILLER_229_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29470_ _35011_/Q _29469_/X _29482_/S VGND VGND VPWR VPWR _29471_/A sky130_fd_sc_hd__mux2_1
X_22914_ _22914_/A VGND VGND VPWR VPWR _32030_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26682_ _33775_/Q _23316_/X _26690_/S VGND VGND VPWR VPWR _26683_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23894_ _22959_/X _32493_/Q _23906_/S VGND VGND VPWR VPWR _23895_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28421_ _27701_/X _34537_/Q _28421_/S VGND VGND VPWR VPWR _28422_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25633_ _25633_/A VGND VGND VPWR VPWR _33280_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22845_ _20660_/X _22843_/X _22844_/X _20672_/X VGND VGND VPWR VPWR _22845_/X sky130_fd_sc_hd__a22o_1
XFILLER_227_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28352_ _27797_/X _34504_/Q _28370_/S VGND VGND VPWR VPWR _28353_/A sky130_fd_sc_hd__mux2_1
X_25564_ _25675_/S VGND VGND VPWR VPWR _25583_/S sky130_fd_sc_hd__buf_4
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22776_ _35474_/Q _35410_/Q _35346_/Q _35282_/Q _22560_/X _22561_/X VGND VGND VPWR
+ VPWR _22776_/X sky130_fd_sc_hd__mux4_1
XFILLER_13_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27303_ _34038_/Q _27134_/X _27317_/S VGND VGND VPWR VPWR _27304_/A sky130_fd_sc_hd__mux2_1
XFILLER_223_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24515_ _24515_/A VGND VGND VPWR VPWR _32784_/D sky130_fd_sc_hd__clkbuf_1
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21727_ _22433_/A VGND VGND VPWR VPWR _21727_/X sky130_fd_sc_hd__buf_4
XFILLER_33_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28283_ _28283_/A VGND VGND VPWR VPWR _34471_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25495_ _24927_/X _33215_/Q _25511_/S VGND VGND VPWR VPWR _25496_/A sky130_fd_sc_hd__mux2_1
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27234_ _30607_/B _31688_/B VGND VGND VPWR VPWR _27367_/S sky130_fd_sc_hd__nor2_8
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21658_ _21654_/X _21657_/X _21379_/X VGND VGND VPWR VPWR _21690_/A sky130_fd_sc_hd__o21ba_1
XFILLER_40_777 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24446_ _24446_/A VGND VGND VPWR VPWR _32751_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27165_ input37/X VGND VGND VPWR VPWR _27165_/X sky130_fd_sc_hd__clkbuf_4
X_20609_ _22560_/A VGND VGND VPWR VPWR _20609_/X sky130_fd_sc_hd__buf_6
XFILLER_240_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24377_ _23064_/X _32719_/Q _24381_/S VGND VGND VPWR VPWR _24378_/A sky130_fd_sc_hd__mux2_1
X_21589_ _32624_/Q _32560_/Q _32496_/Q _35952_/Q _21523_/X _21307_/X VGND VGND VPWR
+ VPWR _21589_/X sky130_fd_sc_hd__mux4_1
XFILLER_197_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26116_ _26116_/A VGND VGND VPWR VPWR _33509_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23328_ _23328_/A VGND VGND VPWR VPWR _32181_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27096_ input13/X VGND VGND VPWR VPWR _27096_/X sky130_fd_sc_hd__buf_2
XFILLER_125_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26047_ _24945_/X _33477_/Q _26051_/S VGND VGND VPWR VPWR _26048_/A sky130_fd_sc_hd__mux2_1
X_23259_ _32159_/Q _23258_/X _23259_/S VGND VGND VPWR VPWR _23260_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17820_ _17816_/X _17819_/X _17504_/X VGND VGND VPWR VPWR _17828_/C sky130_fd_sc_hd__o21ba_1
XTAP_6653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29806_ _29806_/A VGND VGND VPWR VPWR _35161_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27998_ _34336_/Q _27065_/X _28016_/S VGND VGND VPWR VPWR _27999_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_1191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17751_ _17506_/X _17749_/X _17750_/X _17509_/X VGND VGND VPWR VPWR _17751_/X sky130_fd_sc_hd__a22o_1
XFILLER_48_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26949_ _26949_/A VGND VGND VPWR VPWR _33901_/D sky130_fd_sc_hd__clkbuf_1
X_29737_ _35129_/Q _29438_/X _29745_/S VGND VGND VPWR VPWR _29738_/A sky130_fd_sc_hd__mux2_1
XTAP_5974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_844 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16702_ _33384_/Q _33320_/Q _33256_/Q _33192_/Q _16421_/X _16422_/X VGND VGND VPWR
+ VPWR _16702_/X sky130_fd_sc_hd__mux4_1
XFILLER_207_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29668_ _35096_/Q _29336_/X _29682_/S VGND VGND VPWR VPWR _29669_/A sky130_fd_sc_hd__mux2_1
X_17682_ _34435_/Q _36163_/Q _34307_/Q _34243_/Q _17582_/X _17583_/X VGND VGND VPWR
+ VPWR _17682_/X sky130_fd_sc_hd__mux4_1
XFILLER_75_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19421_ _19417_/X _19420_/X _19112_/X VGND VGND VPWR VPWR _19422_/D sky130_fd_sc_hd__o21ba_1
X_28619_ _27794_/X _34631_/Q _28619_/S VGND VGND VPWR VPWR _28620_/A sky130_fd_sc_hd__mux2_1
X_16633_ _33894_/Q _33830_/Q _33766_/Q _36070_/Q _16318_/X _16319_/X VGND VGND VPWR
+ VPWR _16633_/X sky130_fd_sc_hd__mux4_1
XFILLER_223_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29599_ _29599_/A VGND VGND VPWR VPWR _35063_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_222_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19352_ _33650_/Q _33586_/Q _33522_/Q _33458_/Q _19147_/X _19148_/X VGND VGND VPWR
+ VPWR _19352_/X sky130_fd_sc_hd__mux4_1
X_31630_ _27754_/X _36026_/Q _31636_/S VGND VGND VPWR VPWR _31631_/A sky130_fd_sc_hd__mux2_1
XFILLER_216_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16564_ _34148_/Q _34084_/Q _34020_/Q _33956_/Q _16387_/X _16388_/X VGND VGND VPWR
+ VPWR _16564_/X sky130_fd_sc_hd__mux4_1
XFILLER_91_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18303_ _20100_/A VGND VGND VPWR VPWR _18303_/X sky130_fd_sc_hd__buf_4
XFILLER_91_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31561_ _27652_/X _35993_/Q _31573_/S VGND VGND VPWR VPWR _31562_/A sky130_fd_sc_hd__mux2_1
X_19283_ _34160_/Q _34096_/Q _34032_/Q _33968_/Q _19040_/X _19041_/X VGND VGND VPWR
+ VPWR _19283_/X sky130_fd_sc_hd__mux4_1
XFILLER_245_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16495_ _17907_/A VGND VGND VPWR VPWR _16495_/X sky130_fd_sc_hd__buf_4
X_33300_ _36180_/CLK _33300_/D VGND VGND VPWR VPWR _33300_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18234_ _35668_/Q _35028_/Q _34388_/Q _33748_/Q _16112_/X _16113_/X VGND VGND VPWR
+ VPWR _18234_/X sky130_fd_sc_hd__mux4_1
X_30512_ _30512_/A VGND VGND VPWR VPWR _35496_/D sky130_fd_sc_hd__clkbuf_1
X_34280_ _34914_/CLK _34280_/D VGND VGND VPWR VPWR _34280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31492_ _31492_/A VGND VGND VPWR VPWR _35960_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33231_ _34186_/CLK _33231_/D VGND VGND VPWR VPWR _33231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18165_ _18161_/X _18164_/X _17838_/A VGND VGND VPWR VPWR _18187_/A sky130_fd_sc_hd__o21ba_1
X_30443_ _30470_/S VGND VGND VPWR VPWR _30462_/S sky130_fd_sc_hd__buf_4
XFILLER_191_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17116_ _35187_/Q _35123_/Q _35059_/Q _32220_/Q _17010_/X _17011_/X VGND VGND VPWR
+ VPWR _17116_/X sky130_fd_sc_hd__mux4_1
X_33162_ _36040_/CLK _33162_/D VGND VGND VPWR VPWR _33162_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18096_ _18092_/X _18095_/X _17871_/X VGND VGND VPWR VPWR _18097_/D sky130_fd_sc_hd__o21ba_1
XFILLER_176_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30374_ _35431_/Q _29382_/X _30378_/S VGND VGND VPWR VPWR _30375_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32113_ _35953_/CLK _32113_/D VGND VGND VPWR VPWR _32113_/Q sky130_fd_sc_hd__dfxtp_1
X_17047_ _34929_/Q _34865_/Q _34801_/Q _34737_/Q _16807_/X _16808_/X VGND VGND VPWR
+ VPWR _17047_/X sky130_fd_sc_hd__mux4_1
XFILLER_239_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33093_ _35843_/CLK _33093_/D VGND VGND VPWR VPWR _33093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32044_ _35820_/CLK _32044_/D VGND VGND VPWR VPWR _32044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18998_ _18998_/A VGND VGND VPWR VPWR _32423_/D sky130_fd_sc_hd__clkbuf_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35803_ _36059_/CLK _35803_/D VGND VGND VPWR VPWR _35803_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17949_ _17945_/X _17948_/X _17838_/X VGND VGND VPWR VPWR _17973_/A sky130_fd_sc_hd__o21ba_2
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33995_ _34187_/CLK _33995_/D VGND VGND VPWR VPWR _33995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_245_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35734_ _36118_/CLK _35734_/D VGND VGND VPWR VPWR _35734_/Q sky130_fd_sc_hd__dfxtp_1
X_20960_ _20953_/X _20955_/X _20958_/X _20959_/X VGND VGND VPWR VPWR _20960_/X sky130_fd_sc_hd__a22o_1
XFILLER_226_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32946_ _36019_/CLK _32946_/D VGND VGND VPWR VPWR _32946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19619_ _35705_/Q _32214_/Q _35577_/Q _35513_/Q _19617_/X _19618_/X VGND VGND VPWR
+ VPWR _19619_/X sky130_fd_sc_hd__mux4_2
XFILLER_226_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35665_ _35728_/CLK _35665_/D VGND VGND VPWR VPWR _35665_/Q sky130_fd_sc_hd__dfxtp_1
X_20891_ _20885_/X _20890_/X _20644_/X _20646_/X VGND VGND VPWR VPWR _20912_/B sky130_fd_sc_hd__o211a_1
X_32877_ _32877_/CLK _32877_/D VGND VGND VPWR VPWR _32877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22630_ _34701_/Q _34637_/Q _34573_/Q _34509_/Q _22598_/X _22599_/X VGND VGND VPWR
+ VPWR _22630_/X sky130_fd_sc_hd__mux4_1
X_34616_ _35193_/CLK _34616_/D VGND VGND VPWR VPWR _34616_/Q sky130_fd_sc_hd__dfxtp_1
X_31828_ _31828_/A VGND VGND VPWR VPWR _36119_/D sky130_fd_sc_hd__clkbuf_1
X_35596_ _35596_/CLK _35596_/D VGND VGND VPWR VPWR _35596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_722 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22561_ _22561_/A VGND VGND VPWR VPWR _22561_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_94_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31759_ _36087_/Q input27/X _31771_/S VGND VGND VPWR VPWR _31760_/A sky130_fd_sc_hd__mux2_1
X_34547_ _34611_/CLK _34547_/D VGND VGND VPWR VPWR _34547_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_834 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24300_ _22949_/X _32682_/Q _24318_/S VGND VGND VPWR VPWR _24301_/A sky130_fd_sc_hd__mux2_1
X_21512_ _21405_/X _21510_/X _21511_/X _21410_/X VGND VGND VPWR VPWR _21512_/X sky130_fd_sc_hd__a22o_1
X_25280_ _33114_/Q _23243_/X _25290_/S VGND VGND VPWR VPWR _25281_/A sky130_fd_sc_hd__mux2_1
X_22492_ _35465_/Q _35401_/Q _35337_/Q _35273_/Q _22207_/X _22208_/X VGND VGND VPWR
+ VPWR _22492_/X sky130_fd_sc_hd__mux4_1
XFILLER_21_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34478_ _36142_/CLK _34478_/D VGND VGND VPWR VPWR _34478_/Q sky130_fd_sc_hd__dfxtp_1
X_36217_ _36219_/CLK _36217_/D VGND VGND VPWR VPWR _36217_/Q sky130_fd_sc_hd__dfxtp_1
X_24231_ _32651_/Q _23466_/X _24243_/S VGND VGND VPWR VPWR _24232_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21443_ _21439_/X _21442_/X _21412_/X VGND VGND VPWR VPWR _21444_/D sky130_fd_sc_hd__o21ba_1
X_33429_ _36180_/CLK _33429_/D VGND VGND VPWR VPWR _33429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24162_ _32618_/Q _23292_/X _24180_/S VGND VGND VPWR VPWR _24163_/A sky130_fd_sc_hd__mux2_1
XFILLER_175_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21374_ _22433_/A VGND VGND VPWR VPWR _21374_/X sky130_fd_sc_hd__buf_4
X_36148_ _36149_/CLK _36148_/D VGND VGND VPWR VPWR _36148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20325_ _20004_/X _20323_/X _20324_/X _20007_/X VGND VGND VPWR VPWR _20325_/X sky130_fd_sc_hd__a22o_1
X_23113_ _22918_/X _32096_/Q _23131_/S VGND VGND VPWR VPWR _23114_/A sky130_fd_sc_hd__mux2_1
X_24093_ _23052_/X _32587_/Q _24105_/S VGND VGND VPWR VPWR _24094_/A sky130_fd_sc_hd__mux2_1
X_28970_ _28970_/A VGND VGND VPWR VPWR _34795_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36079_ _36079_/CLK _36079_/D VGND VGND VPWR VPWR _36079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23044_ _23042_/X _32072_/Q _23071_/S VGND VGND VPWR VPWR _23045_/A sky130_fd_sc_hd__mux2_1
X_27921_ _27760_/X _34300_/Q _27923_/S VGND VGND VPWR VPWR _27922_/A sky130_fd_sc_hd__mux2_1
X_20256_ _20252_/X _20255_/X _20146_/X _20147_/X VGND VGND VPWR VPWR _20273_/B sky130_fd_sc_hd__o211a_1
XFILLER_135_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27852_ _27658_/X _34267_/Q _27860_/S VGND VGND VPWR VPWR _27853_/A sky130_fd_sc_hd__mux2_1
XTAP_5215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20187_ _20073_/X _20185_/X _20186_/X _20077_/X VGND VGND VPWR VPWR _20187_/X sky130_fd_sc_hd__a22o_1
XTAP_5226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26803_ _26803_/A VGND VGND VPWR VPWR _33832_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27783_ _27782_/X _34243_/Q _27795_/S VGND VGND VPWR VPWR _27784_/A sky130_fd_sc_hd__mux2_1
XTAP_4525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24995_ _24994_/X _32981_/Q _24995_/S VGND VGND VPWR VPWR _24996_/A sky130_fd_sc_hd__mux2_1
XTAP_4536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29522_ _35028_/Q _29521_/X _29525_/S VGND VGND VPWR VPWR _29523_/A sky130_fd_sc_hd__mux2_1
XTAP_4547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26734_ _26761_/S VGND VGND VPWR VPWR _26753_/S sky130_fd_sc_hd__buf_4
XTAP_4558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23946_ _23036_/X _32518_/Q _23948_/S VGND VGND VPWR VPWR _23947_/A sky130_fd_sc_hd__mux2_1
XTAP_3824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29453_ input35/X VGND VGND VPWR VPWR _29453_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_6_0_CLK clkbuf_5_7_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_6_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_205_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26665_ _33767_/Q _23283_/X _26669_/S VGND VGND VPWR VPWR _26666_/A sky130_fd_sc_hd__mux2_1
XFILLER_245_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23877_ _22934_/X _32485_/Q _23885_/S VGND VGND VPWR VPWR _23878_/A sky130_fd_sc_hd__mux2_1
X_28404_ _28404_/A VGND VGND VPWR VPWR _34528_/D sky130_fd_sc_hd__clkbuf_1
X_25616_ _25616_/A VGND VGND VPWR VPWR _33272_/D sky130_fd_sc_hd__clkbuf_1
X_22828_ _21753_/A _22826_/X _22827_/X _21756_/A VGND VGND VPWR VPWR _22828_/X sky130_fd_sc_hd__a22o_1
X_29384_ _29384_/A VGND VGND VPWR VPWR _34983_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26596_ _24954_/X _33736_/Q _26614_/S VGND VGND VPWR VPWR _26597_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_1222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28335_ _27773_/X _34496_/Q _28349_/S VGND VGND VPWR VPWR _28336_/A sky130_fd_sc_hd__mux2_1
X_25547_ _25547_/A VGND VGND VPWR VPWR _33239_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22759_ _33682_/Q _33618_/Q _33554_/Q _33490_/Q _22506_/X _22507_/X VGND VGND VPWR
+ VPWR _22759_/X sky130_fd_sc_hd__mux4_1
XFILLER_198_874 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28266_ _28266_/A VGND VGND VPWR VPWR _34463_/D sky130_fd_sc_hd__clkbuf_1
X_16280_ _33884_/Q _33820_/Q _33756_/Q _36060_/Q _16112_/X _16113_/X VGND VGND VPWR
+ VPWR _16280_/X sky130_fd_sc_hd__mux4_1
X_25478_ _24902_/X _33207_/Q _25490_/S VGND VGND VPWR VPWR _25479_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27217_ input55/X VGND VGND VPWR VPWR _27217_/X sky130_fd_sc_hd__buf_4
X_24429_ _24429_/A VGND VGND VPWR VPWR _32743_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28197_ _28197_/A VGND VGND VPWR VPWR _34430_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27148_ _27148_/A VGND VGND VPWR VPWR _33978_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19970_ _20099_/A VGND VGND VPWR VPWR _19970_/X sky130_fd_sc_hd__buf_4
XFILLER_153_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27079_ _33956_/Q _27078_/X _27094_/S VGND VGND VPWR VPWR _27080_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1018 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18921_ _35173_/Q _35109_/Q _35045_/Q _32165_/Q _18604_/X _18605_/X VGND VGND VPWR
+ VPWR _18921_/X sky130_fd_sc_hd__mux4_1
XTAP_7140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30090_ _35296_/Q _29360_/X _30108_/S VGND VGND VPWR VPWR _30091_/A sky130_fd_sc_hd__mux2_1
XFILLER_134_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18852_ _18597_/X _18850_/X _18851_/X _18600_/X VGND VGND VPWR VPWR _18852_/X sky130_fd_sc_hd__a22o_1
XTAP_6450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17803_ _33415_/Q _33351_/Q _33287_/Q _33223_/Q _17480_/X _17481_/X VGND VGND VPWR
+ VPWR _17803_/X sky130_fd_sc_hd__mux4_1
XTAP_6494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18783_ _18779_/X _18782_/X _18745_/X VGND VGND VPWR VPWR _18791_/C sky130_fd_sc_hd__o21ba_1
XFILLER_79_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15995_ _17800_/A VGND VGND VPWR VPWR _15995_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_95_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17734_ _17728_/X _17733_/X _17485_/X VGND VGND VPWR VPWR _17756_/A sky130_fd_sc_hd__o21ba_1
XTAP_5782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32800_ _35871_/CLK _32800_/D VGND VGND VPWR VPWR _32800_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30992_ _35724_/Q input50/X _31002_/S VGND VGND VPWR VPWR _30993_/A sky130_fd_sc_hd__mux2_1
X_33780_ _36085_/CLK _33780_/D VGND VGND VPWR VPWR _33780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_236_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32731_ _35995_/CLK _32731_/D VGND VGND VPWR VPWR _32731_/Q sky130_fd_sc_hd__dfxtp_1
X_17665_ _17412_/X _17663_/X _17664_/X _17418_/X VGND VGND VPWR VPWR _17665_/X sky130_fd_sc_hd__a22o_1
XFILLER_91_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16616_ _35429_/Q _35365_/Q _35301_/Q _35237_/Q _16548_/X _16549_/X VGND VGND VPWR
+ VPWR _16616_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19404_ _32115_/Q _32307_/Q _32371_/Q _35891_/Q _19227_/X _19368_/X VGND VGND VPWR
+ VPWR _19404_/X sky130_fd_sc_hd__mux4_1
X_32662_ _32856_/CLK _32662_/D VGND VGND VPWR VPWR _32662_/Q sky130_fd_sc_hd__dfxtp_1
X_35450_ _35451_/CLK _35450_/D VGND VGND VPWR VPWR _35450_/Q sky130_fd_sc_hd__dfxtp_1
X_17596_ _17592_/X _17595_/X _17485_/X VGND VGND VPWR VPWR _17620_/A sky130_fd_sc_hd__o21ba_1
XFILLER_189_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34401_ _36128_/CLK _34401_/D VGND VGND VPWR VPWR _34401_/Q sky130_fd_sc_hd__dfxtp_1
X_31613_ _27729_/X _36018_/Q _31615_/S VGND VGND VPWR VPWR _31614_/A sky130_fd_sc_hd__mux2_1
XFILLER_206_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16547_ _16292_/X _16545_/X _16546_/X _16295_/X VGND VGND VPWR VPWR _16547_/X sky130_fd_sc_hd__a22o_1
X_19335_ _19331_/X _19334_/X _19087_/X _19088_/X VGND VGND VPWR VPWR _19350_/B sky130_fd_sc_hd__o211a_1
X_32593_ _35982_/CLK _32593_/D VGND VGND VPWR VPWR _32593_/Q sky130_fd_sc_hd__dfxtp_1
X_35381_ _35446_/CLK _35381_/D VGND VGND VPWR VPWR _35381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34332_ _36060_/CLK _34332_/D VGND VGND VPWR VPWR _34332_/Q sky130_fd_sc_hd__dfxtp_1
X_31544_ _31544_/A VGND VGND VPWR VPWR _35985_/D sky130_fd_sc_hd__clkbuf_1
X_19266_ _35695_/Q _32203_/Q _35567_/Q _35503_/Q _19264_/X _19265_/X VGND VGND VPWR
+ VPWR _19266_/X sky130_fd_sc_hd__mux4_1
X_16478_ _35617_/Q _34977_/Q _34337_/Q _33697_/Q _16438_/X _16439_/X VGND VGND VPWR
+ VPWR _16478_/X sky130_fd_sc_hd__mux4_2
XFILLER_108_1467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18217_ _18217_/A _18217_/B _18217_/C _18217_/D VGND VGND VPWR VPWR _18218_/A sky130_fd_sc_hd__or4_4
X_34263_ _34585_/CLK _34263_/D VGND VGND VPWR VPWR _34263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19197_ _19193_/X _19196_/X _19087_/X _19088_/X VGND VGND VPWR VPWR _19214_/B sky130_fd_sc_hd__o211a_1
X_31475_ _31475_/A VGND VGND VPWR VPWR _35952_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33214_ _33921_/CLK _33214_/D VGND VGND VPWR VPWR _33214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36002_ _36002_/CLK _36002_/D VGND VGND VPWR VPWR _36002_/Q sky130_fd_sc_hd__dfxtp_1
X_18148_ _16001_/X _18146_/X _18147_/X _16007_/X VGND VGND VPWR VPWR _18148_/X sky130_fd_sc_hd__a22o_1
X_30426_ _30426_/A VGND VGND VPWR VPWR _35455_/D sky130_fd_sc_hd__clkbuf_1
X_34194_ _34897_/CLK _34194_/D VGND VGND VPWR VPWR _34194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33145_ _36025_/CLK _33145_/D VGND VGND VPWR VPWR _33145_/Q sky130_fd_sc_hd__dfxtp_1
X_30357_ _35423_/Q _29357_/X _30357_/S VGND VGND VPWR VPWR _30358_/A sky130_fd_sc_hd__mux2_1
X_18079_ _32143_/Q _32335_/Q _32399_/Q _35919_/Q _17986_/X _17774_/X VGND VGND VPWR
+ VPWR _18079_/X sky130_fd_sc_hd__mux4_1
XFILLER_160_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20110_ _32135_/Q _32327_/Q _32391_/Q _35911_/Q _19933_/X _20074_/X VGND VGND VPWR
+ VPWR _20110_/X sky130_fd_sc_hd__mux4_1
X_33076_ _35698_/CLK _33076_/D VGND VGND VPWR VPWR _33076_/Q sky130_fd_sc_hd__dfxtp_1
X_21090_ _21086_/X _21089_/X _21059_/X VGND VGND VPWR VPWR _21091_/D sky130_fd_sc_hd__o21ba_1
XFILLER_125_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30288_ _35390_/Q _29453_/X _30306_/S VGND VGND VPWR VPWR _30289_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32027_ _34007_/CLK _32027_/D VGND VGND VPWR VPWR _32027_/Q sky130_fd_sc_hd__dfxtp_1
X_20041_ _20037_/X _20040_/X _19793_/X _19794_/X VGND VGND VPWR VPWR _20056_/B sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_140_CLK clkbuf_6_22__f_CLK/X VGND VGND VPWR VPWR _35993_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1039 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23800_ _23800_/A VGND VGND VPWR VPWR _32385_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24780_ _23061_/X _32910_/Q _24786_/S VGND VGND VPWR VPWR _24781_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33978_ _35320_/CLK _33978_/D VGND VGND VPWR VPWR _33978_/Q sky130_fd_sc_hd__dfxtp_1
X_21992_ _35451_/Q _35387_/Q _35323_/Q _35259_/Q _21854_/X _21855_/X VGND VGND VPWR
+ VPWR _21992_/X sky130_fd_sc_hd__mux4_1
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35717_ _35717_/CLK _35717_/D VGND VGND VPWR VPWR _35717_/Q sky130_fd_sc_hd__dfxtp_1
X_23731_ _23731_/A VGND VGND VPWR VPWR _32352_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20943_ _20939_/X _20942_/X _20704_/X VGND VGND VPWR VPWR _20944_/D sky130_fd_sc_hd__o21ba_1
X_32929_ _36003_/CLK _32929_/D VGND VGND VPWR VPWR _32929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26450_ _26450_/A VGND VGND VPWR VPWR _33667_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35648_ _35648_/CLK _35648_/D VGND VGND VPWR VPWR _35648_/Q sky130_fd_sc_hd__dfxtp_1
X_23662_ _23662_/A VGND VGND VPWR VPWR _32321_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20874_ _20874_/A _20874_/B _20874_/C _20874_/D VGND VGND VPWR VPWR _20875_/A sky130_fd_sc_hd__or4_2
XFILLER_53_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25401_ _33172_/Q _23495_/X _25403_/S VGND VGND VPWR VPWR _25402_/A sky130_fd_sc_hd__mux2_1
X_22613_ _33933_/Q _33869_/Q _33805_/Q _36109_/Q _22330_/X _22331_/X VGND VGND VPWR
+ VPWR _22613_/X sky130_fd_sc_hd__mux4_1
XFILLER_228_1282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26381_ _26381_/A VGND VGND VPWR VPWR _33634_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23593_ _23593_/A VGND VGND VPWR VPWR _32288_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35579_ _35709_/CLK _35579_/D VGND VGND VPWR VPWR _35579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28120_ _27655_/X _34394_/Q _28130_/S VGND VGND VPWR VPWR _28121_/A sky130_fd_sc_hd__mux2_1
X_25332_ _33139_/Q _23384_/X _25332_/S VGND VGND VPWR VPWR _25333_/A sky130_fd_sc_hd__mux2_1
X_22544_ _34187_/Q _34123_/Q _34059_/Q _33995_/Q _22399_/X _22400_/X VGND VGND VPWR
+ VPWR _22544_/X sky130_fd_sc_hd__mux4_1
XFILLER_194_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28051_ _28051_/A VGND VGND VPWR VPWR _34361_/D sky130_fd_sc_hd__clkbuf_1
X_25263_ _33107_/Q _23492_/X _25267_/S VGND VGND VPWR VPWR _25264_/A sky130_fd_sc_hd__mux2_1
X_22475_ _33673_/Q _33609_/Q _33545_/Q _33481_/Q _22153_/X _22154_/X VGND VGND VPWR
+ VPWR _22475_/X sky130_fd_sc_hd__mux4_1
XFILLER_210_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27002_ _33927_/Q _23450_/X _27002_/S VGND VGND VPWR VPWR _27003_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24214_ _32643_/Q _23438_/X _24222_/S VGND VGND VPWR VPWR _24215_/A sky130_fd_sc_hd__mux2_1
XFILLER_136_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21426_ _32107_/Q _32299_/Q _32363_/Q _35883_/Q _21174_/X _21315_/X VGND VGND VPWR
+ VPWR _21426_/X sky130_fd_sc_hd__mux4_1
X_25194_ _33074_/Q _23381_/X _25196_/S VGND VGND VPWR VPWR _25195_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_955 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24145_ _32610_/Q _23268_/X _24159_/S VGND VGND VPWR VPWR _24146_/A sky130_fd_sc_hd__mux2_1
X_21357_ _21245_/X _21355_/X _21356_/X _21248_/X VGND VGND VPWR VPWR _21357_/X sky130_fd_sc_hd__a22o_1
XFILLER_163_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20308_ _20308_/A VGND VGND VPWR VPWR _32460_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_123_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24076_ _23027_/X _32579_/Q _24084_/S VGND VGND VPWR VPWR _24077_/A sky130_fd_sc_hd__mux2_1
X_28953_ _28953_/A VGND VGND VPWR VPWR _34787_/D sky130_fd_sc_hd__clkbuf_1
X_21288_ _21250_/X _21286_/X _21287_/X _21253_/X VGND VGND VPWR VPWR _21288_/X sky130_fd_sc_hd__a22o_1
XFILLER_235_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20239_ _20164_/X _20237_/X _20238_/X _20169_/X VGND VGND VPWR VPWR _20239_/X sky130_fd_sc_hd__a22o_1
X_23027_ input40/X VGND VGND VPWR VPWR _23027_/X sky130_fd_sc_hd__buf_2
X_27904_ _27973_/S VGND VGND VPWR VPWR _27923_/S sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_131_CLK clkbuf_6_23__f_CLK/X VGND VGND VPWR VPWR _34904_/CLK sky130_fd_sc_hd__clkbuf_16
X_28884_ _34755_/Q _27174_/X _28892_/S VGND VGND VPWR VPWR _28885_/A sky130_fd_sc_hd__mux2_1
XTAP_5001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27835_ _27834_/X _34260_/Q _27838_/S VGND VGND VPWR VPWR _27836_/A sky130_fd_sc_hd__mux2_1
XTAP_4300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27766_ input35/X VGND VGND VPWR VPWR _27766_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24978_ _24978_/A VGND VGND VPWR VPWR _32975_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29505_ _29505_/A VGND VGND VPWR VPWR _35022_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26717_ _26717_/A VGND VGND VPWR VPWR _33791_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23929_ _23977_/S VGND VGND VPWR VPWR _23948_/S sky130_fd_sc_hd__buf_4
XFILLER_206_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27697_ _27697_/A VGND VGND VPWR VPWR _34215_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17450_ _33405_/Q _33341_/Q _33277_/Q _33213_/Q _17127_/X _17128_/X VGND VGND VPWR
+ VPWR _17450_/X sky130_fd_sc_hd__mux4_1
X_29436_ _35000_/Q _29435_/X _29451_/S VGND VGND VPWR VPWR _29437_/A sky130_fd_sc_hd__mux2_1
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26648_ _33759_/Q _23258_/X _26648_/S VGND VGND VPWR VPWR _26649_/A sky130_fd_sc_hd__mux2_1
XTAP_3698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16401_ _16397_/X _16400_/X _16044_/X _16046_/X VGND VGND VPWR VPWR _16416_/B sky130_fd_sc_hd__o211a_1
XTAP_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17381_ _17375_/X _17380_/X _17132_/X VGND VGND VPWR VPWR _17403_/A sky130_fd_sc_hd__o21ba_1
X_29367_ input4/X VGND VGND VPWR VPWR _29367_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_198_CLK clkbuf_6_49__f_CLK/X VGND VGND VPWR VPWR _35596_/CLK sky130_fd_sc_hd__clkbuf_16
X_26579_ _24930_/X _33728_/Q _26593_/S VGND VGND VPWR VPWR _26580_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19120_ _33899_/Q _33835_/Q _33771_/Q _36075_/Q _18971_/X _18972_/X VGND VGND VPWR
+ VPWR _19120_/X sky130_fd_sc_hd__mux4_1
X_16332_ _16292_/X _16330_/X _16331_/X _16295_/X VGND VGND VPWR VPWR _16332_/X sky130_fd_sc_hd__a22o_1
X_28318_ _27748_/X _34488_/Q _28328_/S VGND VGND VPWR VPWR _28319_/A sky130_fd_sc_hd__mux2_1
X_29298_ _29298_/A VGND VGND VPWR VPWR _34951_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_203_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19051_ _32105_/Q _32297_/Q _32361_/Q _35881_/Q _18874_/X _19015_/X VGND VGND VPWR
+ VPWR _19051_/X sky130_fd_sc_hd__mux4_1
X_28249_ _27646_/X _34455_/Q _28265_/S VGND VGND VPWR VPWR _28250_/A sky130_fd_sc_hd__mux2_1
X_16263_ _35419_/Q _35355_/Q _35291_/Q _35227_/Q _16195_/X _16196_/X VGND VGND VPWR
+ VPWR _16263_/X sky130_fd_sc_hd__mux4_1
XFILLER_16_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18002_ _17859_/X _18000_/X _18001_/X _17862_/X VGND VGND VPWR VPWR _18002_/X sky130_fd_sc_hd__a22o_1
XFILLER_187_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31260_ _31260_/A VGND VGND VPWR VPWR _35850_/D sky130_fd_sc_hd__clkbuf_1
X_16194_ _16048_/X _16192_/X _16193_/X _16058_/X VGND VGND VPWR VPWR _16194_/X sky130_fd_sc_hd__a22o_1
XFILLER_126_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30211_ _30211_/A VGND VGND VPWR VPWR _35353_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_370_CLK clkbuf_6_43__f_CLK/X VGND VGND VPWR VPWR _36153_/CLK sky130_fd_sc_hd__clkbuf_16
X_31191_ _31281_/S VGND VGND VPWR VPWR _31210_/S sky130_fd_sc_hd__buf_4
XFILLER_99_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30142_ _35321_/Q _29438_/X _30150_/S VGND VGND VPWR VPWR _30143_/A sky130_fd_sc_hd__mux2_1
X_19953_ _19949_/X _19952_/X _19818_/X VGND VGND VPWR VPWR _19954_/D sky130_fd_sc_hd__o21ba_1
XFILLER_141_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18904_ _32613_/Q _32549_/Q _32485_/Q _35941_/Q _18870_/X _18654_/X VGND VGND VPWR
+ VPWR _18904_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_122_CLK clkbuf_6_21__f_CLK/X VGND VGND VPWR VPWR _36125_/CLK sky130_fd_sc_hd__clkbuf_16
X_30073_ _35288_/Q _29336_/X _30087_/S VGND VGND VPWR VPWR _30074_/A sky130_fd_sc_hd__mux2_1
X_34950_ _36165_/CLK _34950_/D VGND VGND VPWR VPWR _34950_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19884_ _34432_/Q _36160_/Q _34304_/Q _34240_/Q _19882_/X _19883_/X VGND VGND VPWR
+ VPWR _19884_/X sky130_fd_sc_hd__mux4_1
XFILLER_132_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33901_ _34093_/CLK _33901_/D VGND VGND VPWR VPWR _33901_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_1359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18835_ _33891_/Q _33827_/Q _33763_/Q _36067_/Q _18618_/X _18619_/X VGND VGND VPWR
+ VPWR _18835_/X sky130_fd_sc_hd__mux4_1
XTAP_6280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34881_ _36104_/CLK _34881_/D VGND VGND VPWR VPWR _34881_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33832_ _33897_/CLK _33832_/D VGND VGND VPWR VPWR _33832_/Q sky130_fd_sc_hd__dfxtp_1
X_18766_ _33377_/Q _33313_/Q _33249_/Q _33185_/Q _18721_/X _18722_/X VGND VGND VPWR
+ VPWR _18766_/X sky130_fd_sc_hd__mux4_1
XTAP_5590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_780 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17717_ _17717_/A VGND VGND VPWR VPWR _17717_/X sky130_fd_sc_hd__buf_4
X_30975_ _35716_/Q input41/X _30981_/S VGND VGND VPWR VPWR _30976_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33763_ _33827_/CLK _33763_/D VGND VGND VPWR VPWR _33763_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18697_ _18653_/X _18695_/X _18696_/X _18659_/X VGND VGND VPWR VPWR _18697_/X sky130_fd_sc_hd__a22o_1
XFILLER_36_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35502_ _35566_/CLK _35502_/D VGND VGND VPWR VPWR _35502_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32714_ _32906_/CLK _32714_/D VGND VGND VPWR VPWR _32714_/Q sky130_fd_sc_hd__dfxtp_1
X_17648_ _35202_/Q _35138_/Q _35074_/Q _32258_/Q _17363_/X _17364_/X VGND VGND VPWR
+ VPWR _17648_/X sky130_fd_sc_hd__mux4_1
X_33694_ _35615_/CLK _33694_/D VGND VGND VPWR VPWR _33694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_212_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35433_ _35433_/CLK _35433_/D VGND VGND VPWR VPWR _35433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17579_ _34688_/Q _34624_/Q _34560_/Q _34496_/Q _17292_/X _17293_/X VGND VGND VPWR
+ VPWR _17579_/X sky130_fd_sc_hd__mux4_1
X_32645_ _36038_/CLK _32645_/D VGND VGND VPWR VPWR _32645_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_189_CLK clkbuf_6_48__f_CLK/X VGND VGND VPWR VPWR _35983_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_195_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19318_ _19318_/A _19318_/B _19318_/C _19318_/D VGND VGND VPWR VPWR _19319_/A sky130_fd_sc_hd__or4_4
XFILLER_188_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20590_ _22371_/A VGND VGND VPWR VPWR _22510_/A sky130_fd_sc_hd__buf_12
X_32576_ _36031_/CLK _32576_/D VGND VGND VPWR VPWR _32576_/Q sky130_fd_sc_hd__dfxtp_1
X_35364_ _35817_/CLK _35364_/D VGND VGND VPWR VPWR _35364_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_984 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34315_ _36173_/CLK _34315_/D VGND VGND VPWR VPWR _34315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31527_ _27801_/X _35977_/Q _31543_/S VGND VGND VPWR VPWR _31528_/A sky130_fd_sc_hd__mux2_1
X_19249_ _19249_/A VGND VGND VPWR VPWR _32430_/D sky130_fd_sc_hd__clkbuf_1
X_35295_ _35743_/CLK _35295_/D VGND VGND VPWR VPWR _35295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22260_ _33923_/Q _33859_/Q _33795_/Q _36099_/Q _21977_/X _21978_/X VGND VGND VPWR
+ VPWR _22260_/X sky130_fd_sc_hd__mux4_1
X_34246_ _36165_/CLK _34246_/D VGND VGND VPWR VPWR _34246_/Q sky130_fd_sc_hd__dfxtp_1
X_31458_ _31458_/A VGND VGND VPWR VPWR _35944_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21211_ _22399_/A VGND VGND VPWR VPWR _21211_/X sky130_fd_sc_hd__buf_4
X_30409_ _30409_/A VGND VGND VPWR VPWR _35447_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_247_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22191_ _34177_/Q _34113_/Q _34049_/Q _33985_/Q _22046_/X _22047_/X VGND VGND VPWR
+ VPWR _22191_/X sky130_fd_sc_hd__mux4_1
X_34177_ _34177_/CLK _34177_/D VGND VGND VPWR VPWR _34177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31389_ _31416_/S VGND VGND VPWR VPWR _31408_/S sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_361_CLK clkbuf_6_46__f_CLK/X VGND VGND VPWR VPWR _36026_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_160_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21142_ _32867_/Q _32803_/Q _32739_/Q _32675_/Q _20887_/X _20888_/X VGND VGND VPWR
+ VPWR _21142_/X sky130_fd_sc_hd__mux4_1
XFILLER_104_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_958 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33128_ _36011_/CLK _33128_/D VGND VGND VPWR VPWR _33128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_113_CLK clkbuf_6_20__f_CLK/X VGND VGND VPWR VPWR _35482_/CLK sky130_fd_sc_hd__clkbuf_16
X_25950_ _25950_/A VGND VGND VPWR VPWR _33430_/D sky130_fd_sc_hd__clkbuf_1
X_21073_ _32097_/Q _32289_/Q _32353_/Q _35873_/Q _20821_/X _20962_/X VGND VGND VPWR
+ VPWR _21073_/X sky130_fd_sc_hd__mux4_1
X_33059_ _35684_/CLK _33059_/D VGND VGND VPWR VPWR _33059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20024_ _20024_/A _20024_/B _20024_/C _20024_/D VGND VGND VPWR VPWR _20025_/A sky130_fd_sc_hd__or4_2
XFILLER_8_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24901_ _24901_/A VGND VGND VPWR VPWR _32950_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25881_ _24899_/X _33398_/Q _25895_/S VGND VGND VPWR VPWR _25882_/A sky130_fd_sc_hd__mux2_1
X_27620_ _27620_/A VGND VGND VPWR VPWR _34188_/D sky130_fd_sc_hd__clkbuf_1
X_24832_ _24830_/X _32928_/Q _24859_/S VGND VGND VPWR VPWR _24833_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27551_ _27551_/A VGND VGND VPWR VPWR _34155_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24763_ _23036_/X _32902_/Q _24765_/S VGND VGND VPWR VPWR _24764_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21975_ _21799_/X _21973_/X _21974_/X _21804_/X VGND VGND VPWR VPWR _21975_/X sky130_fd_sc_hd__a22o_1
XFILLER_55_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26502_ _26502_/A VGND VGND VPWR VPWR _33691_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23714_ _23714_/A VGND VGND VPWR VPWR _32344_/D sky130_fd_sc_hd__clkbuf_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27482_ _34123_/Q _27199_/X _27494_/S VGND VGND VPWR VPWR _27483_/A sky130_fd_sc_hd__mux2_1
X_20926_ _32093_/Q _32285_/Q _32349_/Q _35869_/Q _20821_/X _22467_/A VGND VGND VPWR
+ VPWR _20926_/X sky130_fd_sc_hd__mux4_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24694_ _22934_/X _32869_/Q _24702_/S VGND VGND VPWR VPWR _24695_/A sky130_fd_sc_hd__mux2_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29221_ _29221_/A VGND VGND VPWR VPWR _34914_/D sky130_fd_sc_hd__clkbuf_1
X_26433_ _26433_/A VGND VGND VPWR VPWR _33659_/D sky130_fd_sc_hd__clkbuf_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23645_ _23645_/A VGND VGND VPWR VPWR _32313_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_242_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20857_ _20853_/X _20856_/X _20644_/X _20646_/X VGND VGND VPWR VPWR _20874_/B sky130_fd_sc_hd__o211a_1
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29152_ _34882_/Q _27171_/X _29162_/S VGND VGND VPWR VPWR _29153_/A sky130_fd_sc_hd__mux2_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26364_ _26364_/A VGND VGND VPWR VPWR _33626_/D sky130_fd_sc_hd__clkbuf_1
X_23576_ _23576_/A VGND VGND VPWR VPWR _32280_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20788_ _32089_/Q _32281_/Q _32345_/Q _35865_/Q _20632_/X _22467_/A VGND VGND VPWR
+ VPWR _20788_/X sky130_fd_sc_hd__mux4_1
XFILLER_74_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28103_ _28103_/A VGND VGND VPWR VPWR _34386_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25315_ _25315_/A VGND VGND VPWR VPWR _33130_/D sky130_fd_sc_hd__clkbuf_1
X_22527_ _22304_/X _22525_/X _22526_/X _22307_/X VGND VGND VPWR VPWR _22527_/X sky130_fd_sc_hd__a22o_1
XFILLER_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29083_ _34849_/Q _27069_/X _29099_/S VGND VGND VPWR VPWR _29084_/A sky130_fd_sc_hd__mux2_1
X_26295_ _26295_/A VGND VGND VPWR VPWR _33594_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28034_ _28034_/A VGND VGND VPWR VPWR _34353_/D sky130_fd_sc_hd__clkbuf_1
X_25246_ _25246_/A VGND VGND VPWR VPWR _33098_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22458_ _22453_/X _22456_/X _22457_/X VGND VGND VPWR VPWR _22473_/C sky130_fd_sc_hd__o21ba_1
XFILLER_170_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21409_ _34922_/Q _34858_/Q _34794_/Q _34730_/Q _21407_/X _21408_/X VGND VGND VPWR
+ VPWR _21409_/X sky130_fd_sc_hd__mux4_1
XFILLER_68_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25177_ _25267_/S VGND VGND VPWR VPWR _25196_/S sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_352_CLK clkbuf_6_47__f_CLK/X VGND VGND VPWR VPWR _36029_/CLK sky130_fd_sc_hd__clkbuf_16
X_22389_ _34694_/Q _34630_/Q _34566_/Q _34502_/Q _22245_/X _22246_/X VGND VGND VPWR
+ VPWR _22389_/X sky130_fd_sc_hd__mux4_1
XFILLER_136_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24128_ _32602_/Q _23243_/X _24138_/S VGND VGND VPWR VPWR _24129_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29985_ _29985_/A VGND VGND VPWR VPWR _35246_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28936_ _28936_/A VGND VGND VPWR VPWR _34779_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_104_CLK clkbuf_leaf_99_CLK/A VGND VGND VPWR VPWR _36057_/CLK sky130_fd_sc_hd__clkbuf_16
X_16950_ _33647_/Q _33583_/Q _33519_/Q _33455_/Q _16847_/X _16848_/X VGND VGND VPWR
+ VPWR _16950_/X sky130_fd_sc_hd__mux4_1
X_24059_ _23002_/X _32571_/Q _24063_/S VGND VGND VPWR VPWR _24060_/A sky130_fd_sc_hd__mux2_1
XFILLER_238_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16881_ _16875_/X _16880_/X _16812_/X VGND VGND VPWR VPWR _16882_/D sky130_fd_sc_hd__o21ba_1
XFILLER_131_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28867_ _34747_/Q _27149_/X _28871_/S VGND VGND VPWR VPWR _28868_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18620_ _33885_/Q _33821_/Q _33757_/Q _36061_/Q _18618_/X _18619_/X VGND VGND VPWR
+ VPWR _18620_/X sky130_fd_sc_hd__mux4_1
X_27818_ _27818_/A VGND VGND VPWR VPWR _34254_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28798_ _34714_/Q _27047_/X _28808_/S VGND VGND VPWR VPWR _28799_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18551_ _32603_/Q _32539_/Q _32475_/Q _35931_/Q _18517_/X _20017_/A VGND VGND VPWR
+ VPWR _18551_/X sky130_fd_sc_hd__mux4_1
XTAP_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27749_ _27748_/X _34232_/Q _27764_/S VGND VGND VPWR VPWR _27750_/A sky130_fd_sc_hd__mux2_1
XTAP_4196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17502_ _33086_/Q _32062_/Q _35838_/Q _35774_/Q _17431_/X _17432_/X VGND VGND VPWR
+ VPWR _17502_/X sky130_fd_sc_hd__mux4_1
XTAP_3473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18482_ _33881_/Q _33817_/Q _33753_/Q _36057_/Q _18412_/X _18413_/X VGND VGND VPWR
+ VPWR _18482_/X sky130_fd_sc_hd__mux4_1
X_30760_ _35614_/Q input63/X _30762_/S VGND VGND VPWR VPWR _30761_/A sky130_fd_sc_hd__mux2_1
XTAP_3484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_923 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ _33084_/Q _32060_/Q _35836_/Q _35772_/Q _17431_/X _17432_/X VGND VGND VPWR
+ VPWR _17433_/X sky130_fd_sc_hd__mux4_1
X_29419_ input22/X VGND VGND VPWR VPWR _29419_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30691_ _30691_/A VGND VGND VPWR VPWR _35581_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32430_ _33897_/CLK _32430_/D VGND VGND VPWR VPWR _32430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17364_ _17717_/A VGND VGND VPWR VPWR _17364_/X sky130_fd_sc_hd__buf_6
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16315_ _34141_/Q _34077_/Q _34013_/Q _33949_/Q _16009_/X _16011_/X VGND VGND VPWR
+ VPWR _16315_/X sky130_fd_sc_hd__mux4_1
XFILLER_14_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19103_ _19456_/A VGND VGND VPWR VPWR _19103_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_201_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32361_ _35947_/CLK _32361_/D VGND VGND VPWR VPWR _32361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17295_ _35192_/Q _35128_/Q _35064_/Q _32248_/Q _17010_/X _17011_/X VGND VGND VPWR
+ VPWR _17295_/X sky130_fd_sc_hd__mux4_1
XFILLER_12_1000 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34100_ _34100_/CLK _34100_/D VGND VGND VPWR VPWR _34100_/Q sky130_fd_sc_hd__dfxtp_1
X_19034_ _34920_/Q _34856_/Q _34792_/Q _34728_/Q _18754_/X _18755_/X VGND VGND VPWR
+ VPWR _19034_/X sky130_fd_sc_hd__mux4_1
X_31312_ _27683_/X _35875_/Q _31324_/S VGND VGND VPWR VPWR _31313_/A sky130_fd_sc_hd__mux2_1
X_35080_ _35212_/CLK _35080_/D VGND VGND VPWR VPWR _35080_/Q sky130_fd_sc_hd__dfxtp_1
X_16246_ _16140_/X _16244_/X _16245_/X _16145_/X VGND VGND VPWR VPWR _16246_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32292_ _32356_/CLK _32292_/D VGND VGND VPWR VPWR _32292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34031_ _34991_/CLK _34031_/D VGND VGND VPWR VPWR _34031_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31243_ _31243_/A VGND VGND VPWR VPWR _35842_/D sky130_fd_sc_hd__clkbuf_1
X_16177_ _16177_/A VGND VGND VPWR VPWR _31960_/D sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_343_CLK clkbuf_6_45__f_CLK/X VGND VGND VPWR VPWR _32895_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_127_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput105 _31981_/Q VGND VGND VPWR VPWR D1[23] sky130_fd_sc_hd__buf_2
Xoutput116 _31991_/Q VGND VGND VPWR VPWR D1[33] sky130_fd_sc_hd__buf_2
XFILLER_182_891 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput127 _32001_/Q VGND VGND VPWR VPWR D1[43] sky130_fd_sc_hd__buf_2
XFILLER_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput138 _32011_/Q VGND VGND VPWR VPWR D1[53] sky130_fd_sc_hd__buf_2
XFILLER_217_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31174_ _31174_/A VGND VGND VPWR VPWR _35809_/D sky130_fd_sc_hd__clkbuf_1
Xoutput149 _32021_/Q VGND VGND VPWR VPWR D1[63] sky130_fd_sc_hd__buf_2
XFILLER_47_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30125_ _35313_/Q _29413_/X _30129_/S VGND VGND VPWR VPWR _30126_/A sky130_fd_sc_hd__mux2_1
X_19936_ _19720_/X _19934_/X _19935_/X _19724_/X VGND VGND VPWR VPWR _19936_/X sky130_fd_sc_hd__a22o_1
XFILLER_218_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35982_ _35982_/CLK _35982_/D VGND VGND VPWR VPWR _35982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_218_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30056_ _30056_/A VGND VGND VPWR VPWR _35280_/D sky130_fd_sc_hd__clkbuf_1
X_34933_ _35126_/CLK _34933_/D VGND VGND VPWR VPWR _34933_/Q sky130_fd_sc_hd__dfxtp_1
X_19867_ _19712_/X _19865_/X _19866_/X _19718_/X VGND VGND VPWR VPWR _19867_/X sky130_fd_sc_hd__a22o_1
XFILLER_229_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18818_ _18597_/X _18816_/X _18817_/X _18600_/X VGND VGND VPWR VPWR _18818_/X sky130_fd_sc_hd__a22o_1
XFILLER_7_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34864_ _35439_/CLK _34864_/D VGND VGND VPWR VPWR _34864_/Q sky130_fd_sc_hd__dfxtp_1
X_19798_ _20151_/A VGND VGND VPWR VPWR _19798_/X sky130_fd_sc_hd__buf_4
XFILLER_23_1162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33815_ _34007_/CLK _33815_/D VGND VGND VPWR VPWR _33815_/Q sky130_fd_sc_hd__dfxtp_1
X_18749_ _35168_/Q _35104_/Q _35040_/Q _32160_/Q _18604_/X _18605_/X VGND VGND VPWR
+ VPWR _18749_/X sky130_fd_sc_hd__mux4_1
XFILLER_110_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34795_ _34924_/CLK _34795_/D VGND VGND VPWR VPWR _34795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33746_ _35026_/CLK _33746_/D VGND VGND VPWR VPWR _33746_/Q sky130_fd_sc_hd__dfxtp_1
X_21760_ _22466_/A VGND VGND VPWR VPWR _21760_/X sky130_fd_sc_hd__buf_4
XFILLER_52_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30958_ _35708_/Q input32/X _30960_/S VGND VGND VPWR VPWR _30959_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20711_ _33367_/Q _33303_/Q _33239_/Q _33175_/Q _20602_/X _20603_/X VGND VGND VPWR
+ VPWR _20711_/X sky130_fd_sc_hd__mux4_1
XFILLER_180_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33677_ _34441_/CLK _33677_/D VGND VGND VPWR VPWR _33677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21691_ _21691_/A VGND VGND VPWR VPWR _36210_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_211_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30889_ _35675_/Q input56/X _30897_/S VGND VGND VPWR VPWR _30890_/A sky130_fd_sc_hd__mux2_1
X_35416_ _35799_/CLK _35416_/D VGND VGND VPWR VPWR _35416_/Q sky130_fd_sc_hd__dfxtp_1
X_23430_ _32222_/Q _23429_/X _23451_/S VGND VGND VPWR VPWR _23431_/A sky130_fd_sc_hd__mux2_1
XFILLER_225_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20642_ _20630_/X _20635_/X _20640_/X _20641_/X VGND VGND VPWR VPWR _20642_/X sky130_fd_sc_hd__a22o_1
X_32628_ _36021_/CLK _32628_/D VGND VGND VPWR VPWR _32628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20573_ _34453_/Q _36181_/Q _34325_/Q _34261_/Q _18367_/X _18369_/X VGND VGND VPWR
+ VPWR _20573_/X sky130_fd_sc_hd__mux4_1
X_35347_ _35666_/CLK _35347_/D VGND VGND VPWR VPWR _35347_/Q sky130_fd_sc_hd__dfxtp_1
X_23361_ _23499_/S VGND VGND VPWR VPWR _23385_/S sky130_fd_sc_hd__buf_6
X_32559_ _35952_/CLK _32559_/D VGND VGND VPWR VPWR _32559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25100_ _25100_/A VGND VGND VPWR VPWR _33030_/D sky130_fd_sc_hd__clkbuf_1
X_22312_ _22469_/A VGND VGND VPWR VPWR _22312_/X sky130_fd_sc_hd__clkbuf_4
X_26080_ _24994_/X _33493_/Q _26080_/S VGND VGND VPWR VPWR _26081_/A sky130_fd_sc_hd__mux2_1
X_35278_ _35599_/CLK _35278_/D VGND VGND VPWR VPWR _35278_/Q sky130_fd_sc_hd__dfxtp_1
X_23292_ input13/X VGND VGND VPWR VPWR _23292_/X sky130_fd_sc_hd__buf_4
XFILLER_164_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25031_ _25031_/A VGND VGND VPWR VPWR _32997_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22243_ _21956_/X _22241_/X _22242_/X _21959_/X VGND VGND VPWR VPWR _22243_/X sky130_fd_sc_hd__a22o_1
X_34229_ _35187_/CLK _34229_/D VGND VGND VPWR VPWR _34229_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_334_CLK clkbuf_6_44__f_CLK/X VGND VGND VPWR VPWR _36025_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_192_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22174_ _21951_/X _22172_/X _22173_/X _21954_/X VGND VGND VPWR VPWR _22174_/X sky130_fd_sc_hd__a22o_1
XFILLER_127_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21125_ _34402_/Q _36130_/Q _34274_/Q _34210_/Q _21123_/X _21124_/X VGND VGND VPWR
+ VPWR _21125_/X sky130_fd_sc_hd__mux4_1
XFILLER_105_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29770_ _29770_/A VGND VGND VPWR VPWR _35144_/D sky130_fd_sc_hd__clkbuf_1
X_26982_ _26982_/A VGND VGND VPWR VPWR _33917_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25933_ _24976_/X _33423_/Q _25937_/S VGND VGND VPWR VPWR _25934_/A sky130_fd_sc_hd__mux2_1
X_28721_ _28721_/A VGND VGND VPWR VPWR _34678_/D sky130_fd_sc_hd__clkbuf_1
X_21056_ _34912_/Q _34848_/Q _34784_/Q _34720_/Q _21054_/X _21055_/X VGND VGND VPWR
+ VPWR _21056_/X sky130_fd_sc_hd__mux4_2
XFILLER_120_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20007_ _20162_/A VGND VGND VPWR VPWR _20007_/X sky130_fd_sc_hd__clkbuf_4
X_28652_ _28784_/S VGND VGND VPWR VPWR _28671_/S sky130_fd_sc_hd__buf_4
XFILLER_87_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25864_ _24874_/X _33390_/Q _25874_/S VGND VGND VPWR VPWR _25865_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27603_ _27603_/A VGND VGND VPWR VPWR _34180_/D sky130_fd_sc_hd__clkbuf_1
X_24815_ input56/X VGND VGND VPWR VPWR _24815_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_228_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28583_ _28583_/A VGND VGND VPWR VPWR _34613_/D sky130_fd_sc_hd__clkbuf_1
X_25795_ _25795_/A VGND VGND VPWR VPWR _33357_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_189_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27534_ _27534_/A VGND VGND VPWR VPWR _34147_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24746_ _24794_/S VGND VGND VPWR VPWR _24765_/S sky130_fd_sc_hd__buf_4
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21958_ _33082_/Q _32058_/Q _35834_/Q _35770_/Q _21678_/X _21679_/X VGND VGND VPWR
+ VPWR _21958_/X sky130_fd_sc_hd__mux4_1
XFILLER_226_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27465_ _34115_/Q _27174_/X _27473_/S VGND VGND VPWR VPWR _27466_/A sky130_fd_sc_hd__mux2_1
X_20909_ _34908_/Q _34844_/Q _34780_/Q _34716_/Q _20696_/X _20698_/X VGND VGND VPWR
+ VPWR _20909_/X sky130_fd_sc_hd__mux4_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24677_ _22909_/X _32861_/Q _24681_/S VGND VGND VPWR VPWR _24678_/A sky130_fd_sc_hd__mux2_1
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21889_ _33080_/Q _32056_/Q _35832_/Q _35768_/Q _21678_/X _21679_/X VGND VGND VPWR
+ VPWR _21889_/X sky130_fd_sc_hd__mux4_1
XFILLER_202_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29204_ _29204_/A VGND VGND VPWR VPWR _34906_/D sky130_fd_sc_hd__clkbuf_1
X_26416_ _26416_/A VGND VGND VPWR VPWR _33651_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23628_ _23628_/A VGND VGND VPWR VPWR _32305_/D sky130_fd_sc_hd__clkbuf_1
X_27396_ _34082_/Q _27072_/X _27410_/S VGND VGND VPWR VPWR _27397_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_243_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29135_ _34874_/Q _27146_/X _29141_/S VGND VGND VPWR VPWR _29136_/A sky130_fd_sc_hd__mux2_1
X_26347_ _26347_/A VGND VGND VPWR VPWR _33619_/D sky130_fd_sc_hd__clkbuf_1
X_23559_ _32274_/Q _23487_/X _23565_/S VGND VGND VPWR VPWR _23560_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16100_ _17777_/A VGND VGND VPWR VPWR _17163_/A sky130_fd_sc_hd__buf_12
Xinput18 DW[25] VGND VGND VPWR VPWR input18/X sky130_fd_sc_hd__buf_4
XFILLER_35_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29066_ _34841_/Q _27044_/X _29078_/S VGND VGND VPWR VPWR _29067_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput29 DW[35] VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__buf_4
X_17080_ _33074_/Q _32050_/Q _35826_/Q _35762_/Q _17078_/X _17079_/X VGND VGND VPWR
+ VPWR _17080_/X sky130_fd_sc_hd__mux4_1
XFILLER_182_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26278_ _26278_/A VGND VGND VPWR VPWR _33586_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16031_ _16061_/A VGND VGND VPWR VPWR _17986_/A sky130_fd_sc_hd__buf_8
XFILLER_143_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28017_ _28017_/A VGND VGND VPWR VPWR _34345_/D sky130_fd_sc_hd__clkbuf_1
X_25229_ _25229_/A VGND VGND VPWR VPWR _33090_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_325_CLK clkbuf_6_39__f_CLK/X VGND VGND VPWR VPWR _32901_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_109_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17982_ _17982_/A VGND VGND VPWR VPWR _17982_/X sky130_fd_sc_hd__buf_6
XFILLER_111_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29968_ _29968_/A VGND VGND VPWR VPWR _35238_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_991 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19721_ _20074_/A VGND VGND VPWR VPWR _19721_/X sky130_fd_sc_hd__clkbuf_4
X_28919_ _34772_/Q _27226_/X _28921_/S VGND VGND VPWR VPWR _28920_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16933_ _35630_/Q _34990_/Q _34350_/Q _33710_/Q _16791_/X _16792_/X VGND VGND VPWR
+ VPWR _16933_/X sky130_fd_sc_hd__mux4_1
X_29899_ _35206_/Q _29478_/X _29901_/S VGND VGND VPWR VPWR _29900_/A sky130_fd_sc_hd__mux2_1
XFILLER_237_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31930_ _23453_/X _36168_/Q _31948_/S VGND VGND VPWR VPWR _31931_/A sky130_fd_sc_hd__mux2_1
X_19652_ _35706_/Q _32215_/Q _35578_/Q _35514_/Q _19617_/X _19618_/X VGND VGND VPWR
+ VPWR _19652_/X sky130_fd_sc_hd__mux4_1
X_16864_ _16714_/X _16862_/X _16863_/X _16718_/X VGND VGND VPWR VPWR _16864_/X sky130_fd_sc_hd__a22o_1
X_18603_ _34652_/Q _34588_/Q _34524_/Q _34460_/Q _18533_/X _18534_/X VGND VGND VPWR
+ VPWR _18603_/X sky130_fd_sc_hd__mux4_1
XFILLER_20_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16795_ _35434_/Q _35370_/Q _35306_/Q _35242_/Q _16548_/X _16549_/X VGND VGND VPWR
+ VPWR _16795_/X sky130_fd_sc_hd__mux4_1
X_31861_ _31861_/A VGND VGND VPWR VPWR _36135_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19583_ _19367_/X _19581_/X _19582_/X _19371_/X VGND VGND VPWR VPWR _19583_/X sky130_fd_sc_hd__a22o_1
XFILLER_234_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33600_ _34180_/CLK _33600_/D VGND VGND VPWR VPWR _33600_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_248_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18534_ _20299_/A VGND VGND VPWR VPWR _18534_/X sky130_fd_sc_hd__buf_6
X_30812_ _30812_/A VGND VGND VPWR VPWR _35638_/D sky130_fd_sc_hd__clkbuf_1
X_34580_ _34708_/CLK _34580_/D VGND VGND VPWR VPWR _34580_/Q sky130_fd_sc_hd__dfxtp_1
X_31792_ _36103_/Q input44/X _31792_/S VGND VGND VPWR VPWR _31793_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33531_ _33531_/CLK _33531_/D VGND VGND VPWR VPWR _33531_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18465_ _18360_/X _18463_/X _18464_/X _18372_/X VGND VGND VPWR VPWR _18465_/X sky130_fd_sc_hd__a22o_1
X_30743_ _30875_/S VGND VGND VPWR VPWR _30762_/S sky130_fd_sc_hd__clkbuf_8
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17416_ _17774_/A VGND VGND VPWR VPWR _17416_/X sky130_fd_sc_hd__buf_4
X_18396_ _20166_/A VGND VGND VPWR VPWR _18396_/X sky130_fd_sc_hd__buf_4
X_33462_ _33911_/CLK _33462_/D VGND VGND VPWR VPWR _33462_/Q sky130_fd_sc_hd__dfxtp_1
X_30674_ _35573_/Q _29426_/X _30690_/S VGND VGND VPWR VPWR _30675_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35201_ _35715_/CLK _35201_/D VGND VGND VPWR VPWR _35201_/Q sky130_fd_sc_hd__dfxtp_1
X_17347_ _17834_/A VGND VGND VPWR VPWR _17347_/X sky130_fd_sc_hd__clkbuf_4
X_32413_ _33573_/CLK _32413_/D VGND VGND VPWR VPWR _32413_/Q sky130_fd_sc_hd__dfxtp_1
X_36181_ _36181_/CLK _36181_/D VGND VGND VPWR VPWR _36181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33393_ _33393_/CLK _33393_/D VGND VGND VPWR VPWR _33393_/Q sky130_fd_sc_hd__dfxtp_1
X_35132_ _35577_/CLK _35132_/D VGND VGND VPWR VPWR _35132_/Q sky130_fd_sc_hd__dfxtp_1
X_32344_ _35863_/CLK _32344_/D VGND VGND VPWR VPWR _32344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17278_ _33144_/Q _36024_/Q _33016_/Q _32952_/Q _17062_/X _17063_/X VGND VGND VPWR
+ VPWR _17278_/X sky130_fd_sc_hd__mux4_1
XFILLER_179_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16229_ _35418_/Q _35354_/Q _35290_/Q _35226_/Q _16195_/X _16196_/X VGND VGND VPWR
+ VPWR _16229_/X sky130_fd_sc_hd__mux4_1
X_19017_ _32872_/Q _32808_/Q _32744_/Q _32680_/Q _18940_/X _18941_/X VGND VGND VPWR
+ VPWR _19017_/X sky130_fd_sc_hd__mux4_1
X_32275_ _36114_/CLK _32275_/D VGND VGND VPWR VPWR _32275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_316_CLK clkbuf_6_48__f_CLK/X VGND VGND VPWR VPWR _35916_/CLK sky130_fd_sc_hd__clkbuf_16
X_35063_ _35191_/CLK _35063_/D VGND VGND VPWR VPWR _35063_/Q sky130_fd_sc_hd__dfxtp_1
X_34014_ _36188_/CLK _34014_/D VGND VGND VPWR VPWR _34014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31226_ _31226_/A VGND VGND VPWR VPWR _35834_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31157_ _31157_/A VGND VGND VPWR VPWR _35801_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30108_ _35305_/Q _29388_/X _30108_/S VGND VGND VPWR VPWR _30109_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19919_ _19915_/X _19918_/X _19818_/X VGND VGND VPWR VPWR _19920_/D sky130_fd_sc_hd__o21ba_1
X_31088_ _31088_/A VGND VGND VPWR VPWR _35769_/D sky130_fd_sc_hd__clkbuf_1
X_35965_ _35965_/CLK _35965_/D VGND VGND VPWR VPWR _35965_/Q sky130_fd_sc_hd__dfxtp_1
X_30039_ _35272_/Q _29484_/X _30057_/S VGND VGND VPWR VPWR _30040_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34916_ _34918_/CLK _34916_/D VGND VGND VPWR VPWR _34916_/Q sky130_fd_sc_hd__dfxtp_1
X_22930_ _22930_/A VGND VGND VPWR VPWR _32035_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35896_ _35961_/CLK _35896_/D VGND VGND VPWR VPWR _35896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34847_ _34911_/CLK _34847_/D VGND VGND VPWR VPWR _34847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22861_ _21758_/A _22859_/X _22860_/X _21763_/A VGND VGND VPWR VPWR _22861_/X sky130_fd_sc_hd__a22o_1
XFILLER_84_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24600_ _24600_/A VGND VGND VPWR VPWR _32824_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21812_ _32630_/Q _32566_/Q _32502_/Q _35958_/Q _21523_/X _21660_/X VGND VGND VPWR
+ VPWR _21812_/X sky130_fd_sc_hd__mux4_1
X_25580_ _25580_/A VGND VGND VPWR VPWR _33255_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1075 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34778_ _36245_/CLK _34778_/D VGND VGND VPWR VPWR _34778_/Q sky130_fd_sc_hd__dfxtp_1
X_22792_ _33427_/Q _33363_/Q _33299_/Q _33235_/Q _20637_/X _20639_/X VGND VGND VPWR
+ VPWR _22792_/X sky130_fd_sc_hd__mux4_1
XFILLER_243_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24531_ _24531_/A VGND VGND VPWR VPWR _32791_/D sky130_fd_sc_hd__clkbuf_1
XPHY_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33729_ _36099_/CLK _33729_/D VGND VGND VPWR VPWR _33729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21743_ _35700_/Q _32208_/Q _35572_/Q _35508_/Q _21564_/X _21565_/X VGND VGND VPWR
+ VPWR _21743_/X sky130_fd_sc_hd__mux4_1
XPHY_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27250_ _34013_/Q _27056_/X _27254_/S VGND VGND VPWR VPWR _27251_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24462_ _22990_/X _32759_/Q _24474_/S VGND VGND VPWR VPWR _24463_/A sky130_fd_sc_hd__mux2_1
XFILLER_212_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21674_ _35698_/Q _32206_/Q _35570_/Q _35506_/Q _21564_/X _21565_/X VGND VGND VPWR
+ VPWR _21674_/X sky130_fd_sc_hd__mux4_1
X_26201_ _24973_/X _33550_/Q _26207_/S VGND VGND VPWR VPWR _26202_/A sky130_fd_sc_hd__mux2_1
XFILLER_212_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23413_ _23413_/A VGND VGND VPWR VPWR _32216_/D sky130_fd_sc_hd__clkbuf_1
X_27181_ _33989_/Q _27180_/X _27187_/S VGND VGND VPWR VPWR _27182_/A sky130_fd_sc_hd__mux2_1
X_20625_ _22507_/A VGND VGND VPWR VPWR _20625_/X sky130_fd_sc_hd__buf_4
X_24393_ _22879_/X _32726_/Q _24411_/S VGND VGND VPWR VPWR _24394_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26132_ _24871_/X _33517_/Q _26144_/S VGND VGND VPWR VPWR _26133_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23344_ _23344_/A VGND VGND VPWR VPWR _32188_/D sky130_fd_sc_hd__clkbuf_1
X_20556_ _32661_/Q _32597_/Q _32533_/Q _35989_/Q _20282_/X _19177_/A VGND VGND VPWR
+ VPWR _20556_/X sky130_fd_sc_hd__mux4_1
XFILLER_192_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26063_ _26063_/A VGND VGND VPWR VPWR _33484_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_307_CLK clkbuf_6_50__f_CLK/X VGND VGND VPWR VPWR _36039_/CLK sky130_fd_sc_hd__clkbuf_16
X_23275_ _32164_/Q _23274_/X _23290_/S VGND VGND VPWR VPWR _23276_/A sky130_fd_sc_hd__mux2_1
X_20487_ _20487_/A _20487_/B _20487_/C _20487_/D VGND VGND VPWR VPWR _20488_/A sky130_fd_sc_hd__or4_1
XFILLER_118_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25014_ _25014_/A VGND VGND VPWR VPWR _32989_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22226_ _33922_/Q _33858_/Q _33794_/Q _36098_/Q _21977_/X _21978_/X VGND VGND VPWR
+ VPWR _22226_/X sky130_fd_sc_hd__mux4_1
XFILLER_65_1026 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29822_ _35169_/Q _29364_/X _29838_/S VGND VGND VPWR VPWR _29823_/A sky130_fd_sc_hd__mux2_1
XTAP_6824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22157_ _22510_/A VGND VGND VPWR VPWR _22157_/X sky130_fd_sc_hd__clkbuf_4
XTAP_6835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21108_ _20953_/X _21106_/X _21107_/X _20959_/X VGND VGND VPWR VPWR _21108_/X sky130_fd_sc_hd__a22o_1
XTAP_6868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29753_ _29753_/A VGND VGND VPWR VPWR _35136_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_219_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22088_ _33150_/Q _36030_/Q _33022_/Q _32958_/Q _22015_/X _22016_/X VGND VGND VPWR
+ VPWR _22088_/X sky130_fd_sc_hd__mux4_1
X_26965_ _33909_/Q _23393_/X _26981_/S VGND VGND VPWR VPWR _26966_/A sky130_fd_sc_hd__mux2_1
XTAP_6879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28704_ _28704_/A VGND VGND VPWR VPWR _34670_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_247_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25916_ _24951_/X _33415_/Q _25916_/S VGND VGND VPWR VPWR _25917_/A sky130_fd_sc_hd__mux2_1
X_21039_ _22599_/A VGND VGND VPWR VPWR _21039_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_101_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26896_ _33877_/Q _23498_/X _26896_/S VGND VGND VPWR VPWR _26897_/A sky130_fd_sc_hd__mux2_1
XFILLER_208_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29684_ _29795_/S VGND VGND VPWR VPWR _29703_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_235_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28635_ _28635_/A VGND VGND VPWR VPWR _34638_/D sky130_fd_sc_hd__clkbuf_1
X_25847_ _24849_/X _33382_/Q _25853_/S VGND VGND VPWR VPWR _25848_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16580_ _35620_/Q _34980_/Q _34340_/Q _33700_/Q _16438_/X _16439_/X VGND VGND VPWR
+ VPWR _16580_/X sky130_fd_sc_hd__mux4_1
X_25778_ _25778_/A VGND VGND VPWR VPWR _33349_/D sky130_fd_sc_hd__clkbuf_1
X_28566_ _28566_/A VGND VGND VPWR VPWR _34605_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27517_ _27517_/A VGND VGND VPWR VPWR _34139_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24729_ _24729_/A VGND VGND VPWR VPWR _32885_/D sky130_fd_sc_hd__clkbuf_1
X_28497_ _27813_/X _34573_/Q _28505_/S VGND VGND VPWR VPWR _28498_/A sky130_fd_sc_hd__mux2_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18250_ _34197_/Q _34133_/Q _34069_/Q _34005_/Q _16049_/X _16050_/X VGND VGND VPWR
+ VPWR _18250_/X sky130_fd_sc_hd__mux4_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27448_ _34107_/Q _27149_/X _27452_/S VGND VGND VPWR VPWR _27449_/A sky130_fd_sc_hd__mux2_1
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_1100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _17907_/A VGND VGND VPWR VPWR _17201_/X sky130_fd_sc_hd__buf_4
XFILLER_42_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18181_ _35218_/Q _35154_/Q _35090_/Q _32274_/Q _16092_/X _16094_/X VGND VGND VPWR
+ VPWR _18181_/X sky130_fd_sc_hd__mux4_1
XFILLER_54_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27379_ _34074_/Q _27047_/X _27389_/S VGND VGND VPWR VPWR _27380_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_1472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_994 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17132_ _17838_/A VGND VGND VPWR VPWR _17132_/X sky130_fd_sc_hd__buf_2
X_29118_ _34866_/Q _27121_/X _29120_/S VGND VGND VPWR VPWR _29119_/A sky130_fd_sc_hd__mux2_1
XFILLER_200_1008 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30390_ _30390_/A VGND VGND VPWR VPWR _35438_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29049_ _29049_/A VGND VGND VPWR VPWR _34833_/D sky130_fd_sc_hd__clkbuf_1
X_17063_ _17774_/A VGND VGND VPWR VPWR _17063_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_239_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16014_ input69/X input70/X VGND VGND VPWR VPWR _17838_/A sky130_fd_sc_hd__or2b_4
XFILLER_109_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32060_ _32575_/CLK _32060_/D VGND VGND VPWR VPWR _32060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31011_ _31011_/A VGND VGND VPWR VPWR _35733_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17965_ _17959_/X _17964_/X _17857_/X VGND VGND VPWR VPWR _17973_/C sky130_fd_sc_hd__o21ba_1
XFILLER_112_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19704_ _19704_/A VGND VGND VPWR VPWR _32443_/D sky130_fd_sc_hd__clkbuf_4
X_16916_ _33646_/Q _33582_/Q _33518_/Q _33454_/Q _16847_/X _16848_/X VGND VGND VPWR
+ VPWR _16916_/X sky130_fd_sc_hd__mux4_1
XFILLER_61_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35750_ _35817_/CLK _35750_/D VGND VGND VPWR VPWR _35750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32962_ _36034_/CLK _32962_/D VGND VGND VPWR VPWR _32962_/Q sky130_fd_sc_hd__dfxtp_1
X_17896_ _34697_/Q _34633_/Q _34569_/Q _34505_/Q _17645_/X _17646_/X VGND VGND VPWR
+ VPWR _17896_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34701_ _35213_/CLK _34701_/D VGND VGND VPWR VPWR _34701_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31913_ _23429_/X _36160_/Q _31927_/S VGND VGND VPWR VPWR _31914_/A sky130_fd_sc_hd__mux2_1
X_19635_ _33658_/Q _33594_/Q _33530_/Q _33466_/Q _19500_/X _19501_/X VGND VGND VPWR
+ VPWR _19635_/X sky130_fd_sc_hd__mux4_1
XFILLER_65_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16847_ _17906_/A VGND VGND VPWR VPWR _16847_/X sky130_fd_sc_hd__buf_4
X_35681_ _35747_/CLK _35681_/D VGND VGND VPWR VPWR _35681_/Q sky130_fd_sc_hd__dfxtp_1
X_32893_ _32896_/CLK _32893_/D VGND VGND VPWR VPWR _32893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_1132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34632_ _36113_/CLK _34632_/D VGND VGND VPWR VPWR _34632_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31844_ _31844_/A VGND VGND VPWR VPWR _36127_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19566_ _19562_/X _19565_/X _19465_/X VGND VGND VPWR VPWR _19567_/D sky130_fd_sc_hd__o21ba_1
XFILLER_129_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16778_ _16500_/X _16776_/X _16777_/X _16503_/X VGND VGND VPWR VPWR _16778_/X sky130_fd_sc_hd__a22o_1
XFILLER_225_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18517_ _20282_/A VGND VGND VPWR VPWR _18517_/X sky130_fd_sc_hd__buf_6
X_34563_ _36164_/CLK _34563_/D VGND VGND VPWR VPWR _34563_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31775_ _31775_/A VGND VGND VPWR VPWR _36094_/D sky130_fd_sc_hd__clkbuf_1
X_19497_ _19497_/A _19497_/B _19497_/C _19497_/D VGND VGND VPWR VPWR _19498_/A sky130_fd_sc_hd__or4_1
XFILLER_230_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33514_ _35690_/CLK _33514_/D VGND VGND VPWR VPWR _33514_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30726_ _35598_/Q _29503_/X _30732_/S VGND VGND VPWR VPWR _30727_/A sky130_fd_sc_hd__mux2_1
X_18448_ _33368_/Q _33304_/Q _33240_/Q _33176_/Q _18302_/X _18303_/X VGND VGND VPWR
+ VPWR _18448_/X sky130_fd_sc_hd__mux4_1
XFILLER_22_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34494_ _36101_/CLK _34494_/D VGND VGND VPWR VPWR _34494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36233_ _36235_/CLK _36233_/D VGND VGND VPWR VPWR _36233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33445_ _34151_/CLK _33445_/D VGND VGND VPWR VPWR _33445_/Q sky130_fd_sc_hd__dfxtp_1
X_18379_ _20235_/A VGND VGND VPWR VPWR _18379_/X sky130_fd_sc_hd__buf_6
X_30657_ _35565_/Q _29401_/X _30669_/S VGND VGND VPWR VPWR _30658_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_93_CLK clkbuf_leaf_96_CLK/A VGND VGND VPWR VPWR _36191_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_222_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20410_ _32912_/Q _32848_/Q _32784_/Q _32720_/Q _18284_/X _18287_/X VGND VGND VPWR
+ VPWR _20410_/X sky130_fd_sc_hd__mux4_1
X_36164_ _36164_/CLK _36164_/D VGND VGND VPWR VPWR _36164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21390_ _35690_/Q _32197_/Q _35562_/Q _35498_/Q _21211_/X _21212_/X VGND VGND VPWR
+ VPWR _21390_/X sky130_fd_sc_hd__mux4_1
X_30588_ _30588_/A VGND VGND VPWR VPWR _35532_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_179_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33376_ _36066_/CLK _33376_/D VGND VGND VPWR VPWR _33376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_912 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35115_ _35434_/CLK _35115_/D VGND VGND VPWR VPWR _35115_/Q sky130_fd_sc_hd__dfxtp_1
X_20341_ _20205_/X _20339_/X _20340_/X _20210_/X VGND VGND VPWR VPWR _20341_/X sky130_fd_sc_hd__a22o_1
X_32327_ _35976_/CLK _32327_/D VGND VGND VPWR VPWR _32327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36095_ _36095_/CLK _36095_/D VGND VGND VPWR VPWR _36095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1018 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20272_ _20268_/X _20271_/X _20171_/X VGND VGND VPWR VPWR _20273_/D sky130_fd_sc_hd__o21ba_1
XFILLER_179_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23060_ _23060_/A VGND VGND VPWR VPWR _32077_/D sky130_fd_sc_hd__clkbuf_1
X_35046_ _35625_/CLK _35046_/D VGND VGND VPWR VPWR _35046_/Q sky130_fd_sc_hd__dfxtp_1
X_32258_ _34626_/CLK _32258_/D VGND VGND VPWR VPWR _32258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22011_ _22007_/X _22010_/X _21732_/X VGND VGND VPWR VPWR _22043_/A sky130_fd_sc_hd__o21ba_2
XFILLER_68_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31209_ _31209_/A VGND VGND VPWR VPWR _35826_/D sky130_fd_sc_hd__clkbuf_1
X_32189_ _36135_/CLK _32189_/D VGND VGND VPWR VPWR _32189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_1319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1070 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26750_ _26750_/A VGND VGND VPWR VPWR _33807_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_1384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23962_ _23962_/A VGND VGND VPWR VPWR _32525_/D sky130_fd_sc_hd__clkbuf_1
X_35948_ _35949_/CLK _35948_/D VGND VGND VPWR VPWR _35948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25701_ _25701_/A VGND VGND VPWR VPWR _33312_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_245_935 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22913_ _22912_/X _32030_/Q _22916_/S VGND VGND VPWR VPWR _22914_/A sky130_fd_sc_hd__mux2_1
XFILLER_57_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26681_ _26681_/A VGND VGND VPWR VPWR _33774_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23893_ _23893_/A VGND VGND VPWR VPWR _32492_/D sky130_fd_sc_hd__clkbuf_1
X_35879_ _35941_/CLK _35879_/D VGND VGND VPWR VPWR _35879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25632_ _24930_/X _33280_/Q _25646_/S VGND VGND VPWR VPWR _25633_/A sky130_fd_sc_hd__mux2_1
X_28420_ _28420_/A VGND VGND VPWR VPWR _34536_/D sky130_fd_sc_hd__clkbuf_1
X_22844_ _34964_/Q _34900_/Q _34836_/Q _34772_/Q _20683_/X _20685_/X VGND VGND VPWR
+ VPWR _22844_/X sky130_fd_sc_hd__mux4_1
XFILLER_16_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28351_ _28378_/S VGND VGND VPWR VPWR _28370_/S sky130_fd_sc_hd__buf_4
X_25563_ _25563_/A VGND VGND VPWR VPWR _33247_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22775_ _20581_/X _22773_/X _22774_/X _20591_/X VGND VGND VPWR VPWR _22775_/X sky130_fd_sc_hd__a22o_1
XFILLER_140_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27302_ _27302_/A VGND VGND VPWR VPWR _34037_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24514_ _23067_/X _32784_/Q _24516_/S VGND VGND VPWR VPWR _24515_/A sky130_fd_sc_hd__mux2_1
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21726_ _21446_/X _21724_/X _21725_/X _21451_/X VGND VGND VPWR VPWR _21726_/X sky130_fd_sc_hd__a22o_1
X_28282_ _27695_/X _34471_/Q _28286_/S VGND VGND VPWR VPWR _28283_/A sky130_fd_sc_hd__mux2_1
XFILLER_227_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25494_ _25494_/A VGND VGND VPWR VPWR _33214_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27233_ _27233_/A VGND VGND VPWR VPWR _30607_/B sky130_fd_sc_hd__buf_6
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24445_ _22965_/X _32751_/Q _24453_/S VGND VGND VPWR VPWR _24446_/A sky130_fd_sc_hd__mux2_1
X_21657_ _21453_/X _21655_/X _21656_/X _21456_/X VGND VGND VPWR VPWR _21657_/X sky130_fd_sc_hd__a22o_1
XFILLER_71_1041 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_84_CLK clkbuf_leaf_88_CLK/A VGND VGND VPWR VPWR _35999_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_8_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20608_ _20661_/A VGND VGND VPWR VPWR _22560_/A sky130_fd_sc_hd__buf_12
X_27164_ _27164_/A VGND VGND VPWR VPWR _33983_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_240_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24376_ _24376_/A VGND VGND VPWR VPWR _32718_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21588_ _21584_/X _21587_/X _21379_/X VGND VGND VPWR VPWR _21618_/A sky130_fd_sc_hd__o21ba_1
XFILLER_149_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26115_ _24846_/X _33509_/Q _26123_/S VGND VGND VPWR VPWR _26116_/A sky130_fd_sc_hd__mux2_1
X_23327_ _32181_/Q _23246_/X _23335_/S VGND VGND VPWR VPWR _23328_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20539_ _20535_/X _20538_/X _20157_/A VGND VGND VPWR VPWR _20547_/C sky130_fd_sc_hd__o21ba_1
X_27095_ _27095_/A VGND VGND VPWR VPWR _33961_/D sky130_fd_sc_hd__clkbuf_1
X_26046_ _26046_/A VGND VGND VPWR VPWR _33476_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23258_ input64/X VGND VGND VPWR VPWR _23258_/X sky130_fd_sc_hd__buf_4
XFILLER_165_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22209_ _35457_/Q _35393_/Q _35329_/Q _35265_/Q _22207_/X _22208_/X VGND VGND VPWR
+ VPWR _22209_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23189_ _23189_/A VGND VGND VPWR VPWR _32132_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29805_ _35161_/Q _29339_/X _29817_/S VGND VGND VPWR VPWR _29806_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27997_ _28108_/S VGND VGND VPWR VPWR _28016_/S sky130_fd_sc_hd__buf_4
XFILLER_43_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17750_ _35205_/Q _35141_/Q _35077_/Q _32261_/Q _17716_/X _17717_/X VGND VGND VPWR
+ VPWR _17750_/X sky130_fd_sc_hd__mux4_1
X_29736_ _29736_/A VGND VGND VPWR VPWR _35128_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26948_ _33901_/Q _23302_/X _26960_/S VGND VGND VPWR VPWR _26949_/A sky130_fd_sc_hd__mux2_1
XTAP_5964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16701_ _16493_/X _16699_/X _16700_/X _16498_/X VGND VGND VPWR VPWR _16701_/X sky130_fd_sc_hd__a22o_1
XFILLER_47_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29667_ _29667_/A VGND VGND VPWR VPWR _35095_/D sky130_fd_sc_hd__clkbuf_1
X_17681_ _17506_/X _17679_/X _17680_/X _17509_/X VGND VGND VPWR VPWR _17681_/X sky130_fd_sc_hd__a22o_1
X_26879_ _26879_/A VGND VGND VPWR VPWR _33868_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_968 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19420_ _19105_/X _19418_/X _19419_/X _19110_/X VGND VGND VPWR VPWR _19420_/X sky130_fd_sc_hd__a22o_1
X_28618_ _28618_/A VGND VGND VPWR VPWR _34630_/D sky130_fd_sc_hd__clkbuf_1
X_16632_ _33382_/Q _33318_/Q _33254_/Q _33190_/Q _16421_/X _16422_/X VGND VGND VPWR
+ VPWR _16632_/X sky130_fd_sc_hd__mux4_1
XFILLER_63_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29598_ _35063_/Q _29432_/X _29610_/S VGND VGND VPWR VPWR _29599_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19351_ _19351_/A VGND VGND VPWR VPWR _32433_/D sky130_fd_sc_hd__clkbuf_1
X_16563_ _33636_/Q _33572_/Q _33508_/Q _33444_/Q _16494_/X _16495_/X VGND VGND VPWR
+ VPWR _16563_/X sky130_fd_sc_hd__mux4_1
X_28549_ _28549_/A VGND VGND VPWR VPWR _34597_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_245_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18302_ _20099_/A VGND VGND VPWR VPWR _18302_/X sky130_fd_sc_hd__buf_4
XFILLER_206_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31560_ _31560_/A VGND VGND VPWR VPWR _35992_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16494_ _17906_/A VGND VGND VPWR VPWR _16494_/X sky130_fd_sc_hd__buf_6
X_19282_ _33648_/Q _33584_/Q _33520_/Q _33456_/Q _19147_/X _19148_/X VGND VGND VPWR
+ VPWR _19282_/X sky130_fd_sc_hd__mux4_1
XFILLER_43_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18233_ _35732_/Q _32244_/Q _35604_/Q _35540_/Q _15993_/X _15995_/X VGND VGND VPWR
+ VPWR _18233_/X sky130_fd_sc_hd__mux4_1
XFILLER_15_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30511_ _35496_/Q _29385_/X _30513_/S VGND VGND VPWR VPWR _30512_/A sky130_fd_sc_hd__mux2_1
X_31491_ _27748_/X _35960_/Q _31501_/S VGND VGND VPWR VPWR _31492_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_75_CLK clkbuf_leaf_77_CLK/A VGND VGND VPWR VPWR _35861_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_15_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33230_ _33425_/CLK _33230_/D VGND VGND VPWR VPWR _33230_/Q sky130_fd_sc_hd__dfxtp_1
X_30442_ _30442_/A VGND VGND VPWR VPWR _35463_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18164_ _17912_/X _18162_/X _18163_/X _17915_/X VGND VGND VPWR VPWR _18164_/X sky130_fd_sc_hd__a22o_1
XFILLER_157_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_912 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17115_ _34675_/Q _34611_/Q _34547_/Q _34483_/Q _16939_/X _16940_/X VGND VGND VPWR
+ VPWR _17115_/X sky130_fd_sc_hd__mux4_1
X_18095_ _17864_/X _18093_/X _18094_/X _17869_/X VGND VGND VPWR VPWR _18095_/X sky130_fd_sc_hd__a22o_1
X_33161_ _36044_/CLK _33161_/D VGND VGND VPWR VPWR _33161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30373_ _30373_/A VGND VGND VPWR VPWR _35430_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17046_ _34417_/Q _36145_/Q _34289_/Q _34225_/Q _16876_/X _16877_/X VGND VGND VPWR
+ VPWR _17046_/X sky130_fd_sc_hd__mux4_1
X_32112_ _35952_/CLK _32112_/D VGND VGND VPWR VPWR _32112_/Q sky130_fd_sc_hd__dfxtp_1
X_33092_ _35779_/CLK _33092_/D VGND VGND VPWR VPWR _33092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_861 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32043_ _35820_/CLK _32043_/D VGND VGND VPWR VPWR _32043_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18997_ _18997_/A _18997_/B _18997_/C _18997_/D VGND VGND VPWR VPWR _18998_/A sky130_fd_sc_hd__or4_2
XFILLER_97_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35802_ _35802_/CLK _35802_/D VGND VGND VPWR VPWR _35802_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17948_ _17912_/X _17946_/X _17947_/X _17915_/X VGND VGND VPWR VPWR _17948_/X sky130_fd_sc_hd__a22o_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_992 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33994_ _34187_/CLK _33994_/D VGND VGND VPWR VPWR _33994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_245_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35733_ _35733_/CLK _35733_/D VGND VGND VPWR VPWR _35733_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32945_ _36016_/CLK _32945_/D VGND VGND VPWR VPWR _32945_/Q sky130_fd_sc_hd__dfxtp_1
X_17879_ _33929_/Q _33865_/Q _33801_/Q _36105_/Q _17730_/X _17731_/X VGND VGND VPWR
+ VPWR _17879_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_1434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_6_26__f_CLK clkbuf_5_13_0_CLK/X VGND VGND VPWR VPWR clkbuf_leaf_65_CLK/A sky130_fd_sc_hd__clkbuf_16
X_19618_ _20100_/A VGND VGND VPWR VPWR _19618_/X sky130_fd_sc_hd__buf_4
X_35664_ _35664_/CLK _35664_/D VGND VGND VPWR VPWR _35664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20890_ _20630_/X _20886_/X _20889_/X _20641_/X VGND VGND VPWR VPWR _20890_/X sky130_fd_sc_hd__a22o_1
X_32876_ _32913_/CLK _32876_/D VGND VGND VPWR VPWR _32876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1019 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34615_ _35191_/CLK _34615_/D VGND VGND VPWR VPWR _34615_/Q sky130_fd_sc_hd__dfxtp_1
X_31827_ _23234_/X _36119_/Q _31843_/S VGND VGND VPWR VPWR _31828_/A sky130_fd_sc_hd__mux2_1
X_19549_ _19367_/X _19547_/X _19548_/X _19371_/X VGND VGND VPWR VPWR _19549_/X sky130_fd_sc_hd__a22o_1
X_35595_ _35596_/CLK _35595_/D VGND VGND VPWR VPWR _35595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22560_ _22560_/A VGND VGND VPWR VPWR _22560_/X sky130_fd_sc_hd__buf_4
X_34546_ _35056_/CLK _34546_/D VGND VGND VPWR VPWR _34546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31758_ _31758_/A VGND VGND VPWR VPWR _36086_/D sky130_fd_sc_hd__clkbuf_1
X_21511_ _34925_/Q _34861_/Q _34797_/Q _34733_/Q _21407_/X _21408_/X VGND VGND VPWR
+ VPWR _21511_/X sky130_fd_sc_hd__mux4_1
XFILLER_210_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30709_ _35590_/Q _29478_/X _30711_/S VGND VGND VPWR VPWR _30710_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22491_ _22304_/X _22489_/X _22490_/X _22307_/X VGND VGND VPWR VPWR _22491_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34477_ _35181_/CLK _34477_/D VGND VGND VPWR VPWR _34477_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_66_CLK clkbuf_leaf_73_CLK/A VGND VGND VPWR VPWR _35988_/CLK sky130_fd_sc_hd__clkbuf_16
X_31689_ _31821_/S VGND VGND VPWR VPWR _31708_/S sky130_fd_sc_hd__buf_6
XFILLER_107_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36216_ _36219_/CLK _36216_/D VGND VGND VPWR VPWR _36216_/Q sky130_fd_sc_hd__dfxtp_1
X_24230_ _24230_/A VGND VGND VPWR VPWR _32650_/D sky130_fd_sc_hd__clkbuf_1
X_33428_ _36180_/CLK _33428_/D VGND VGND VPWR VPWR _33428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21442_ _21405_/X _21440_/X _21441_/X _21410_/X VGND VGND VPWR VPWR _21442_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36147_ _36147_/CLK _36147_/D VGND VGND VPWR VPWR _36147_/Q sky130_fd_sc_hd__dfxtp_1
X_24161_ _24251_/S VGND VGND VPWR VPWR _24180_/S sky130_fd_sc_hd__buf_4
X_33359_ _33425_/CLK _33359_/D VGND VGND VPWR VPWR _33359_/Q sky130_fd_sc_hd__dfxtp_1
X_21373_ _21093_/X _21371_/X _21372_/X _21098_/X VGND VGND VPWR VPWR _21373_/X sky130_fd_sc_hd__a22o_1
XFILLER_134_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23112_ _23223_/S VGND VGND VPWR VPWR _23131_/S sky130_fd_sc_hd__buf_4
XFILLER_194_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20324_ _35661_/Q _35021_/Q _34381_/Q _33741_/Q _20150_/X _20151_/X VGND VGND VPWR
+ VPWR _20324_/X sky130_fd_sc_hd__mux4_1
X_24092_ _24092_/A VGND VGND VPWR VPWR _32586_/D sky130_fd_sc_hd__clkbuf_1
X_36078_ _36079_/CLK _36078_/D VGND VGND VPWR VPWR _36078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35029_ _35669_/CLK _35029_/D VGND VGND VPWR VPWR _35029_/Q sky130_fd_sc_hd__dfxtp_1
X_23043_ _23083_/S VGND VGND VPWR VPWR _23071_/S sky130_fd_sc_hd__buf_4
XFILLER_150_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27920_ _27920_/A VGND VGND VPWR VPWR _34299_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20255_ _20073_/X _20253_/X _20254_/X _20077_/X VGND VGND VPWR VPWR _20255_/X sky130_fd_sc_hd__a22o_1
XFILLER_103_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27851_ _27851_/A VGND VGND VPWR VPWR _34266_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20186_ _32905_/Q _32841_/Q _32777_/Q _32713_/Q _19999_/X _20000_/X VGND VGND VPWR
+ VPWR _20186_/X sky130_fd_sc_hd__mux4_1
XTAP_5216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26802_ _33832_/Q _23286_/X _26804_/S VGND VGND VPWR VPWR _26803_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24994_ input60/X VGND VGND VPWR VPWR _24994_/X sky130_fd_sc_hd__clkbuf_4
X_27782_ input40/X VGND VGND VPWR VPWR _27782_/X sky130_fd_sc_hd__clkbuf_4
XTAP_4515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29521_ input59/X VGND VGND VPWR VPWR _29521_/X sky130_fd_sc_hd__buf_2
XTAP_4548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26733_ _26733_/A VGND VGND VPWR VPWR _33799_/D sky130_fd_sc_hd__clkbuf_1
X_23945_ _23945_/A VGND VGND VPWR VPWR _32517_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_1466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26664_ _26664_/A VGND VGND VPWR VPWR _33766_/D sky130_fd_sc_hd__clkbuf_1
X_29452_ _29452_/A VGND VGND VPWR VPWR _35005_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23876_ _23876_/A VGND VGND VPWR VPWR _32484_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25615_ _24905_/X _33272_/Q _25625_/S VGND VGND VPWR VPWR _25616_/A sky130_fd_sc_hd__mux2_1
X_28403_ _27673_/X _34528_/Q _28421_/S VGND VGND VPWR VPWR _28404_/A sky130_fd_sc_hd__mux2_1
X_22827_ _33172_/Q _36052_/Q _33044_/Q _32980_/Q _20632_/X _21761_/A VGND VGND VPWR
+ VPWR _22827_/X sky130_fd_sc_hd__mux4_1
XFILLER_60_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26595_ _26622_/S VGND VGND VPWR VPWR _26614_/S sky130_fd_sc_hd__buf_4
X_29383_ _34983_/Q _29382_/X _29389_/S VGND VGND VPWR VPWR _29384_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28334_ _28334_/A VGND VGND VPWR VPWR _34495_/D sky130_fd_sc_hd__clkbuf_1
X_25546_ _24803_/X _33239_/Q _25562_/S VGND VGND VPWR VPWR _25547_/A sky130_fd_sc_hd__mux2_1
X_22758_ _22758_/A VGND VGND VPWR VPWR _36241_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_756 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28265_ _27670_/X _34463_/Q _28265_/S VGND VGND VPWR VPWR _28266_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_1286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21709_ _35635_/Q _34995_/Q _34355_/Q _33715_/Q _21391_/X _21392_/X VGND VGND VPWR
+ VPWR _21709_/X sky130_fd_sc_hd__mux4_1
XFILLER_200_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25477_ _25477_/A VGND VGND VPWR VPWR _33206_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22689_ _22685_/X _22688_/X _22457_/X VGND VGND VPWR VPWR _22697_/C sky130_fd_sc_hd__o21ba_1
XFILLER_8_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_57_CLK clkbuf_leaf_57_CLK/A VGND VGND VPWR VPWR _32873_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_9_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27216_ _27216_/A VGND VGND VPWR VPWR _34000_/D sky130_fd_sc_hd__clkbuf_1
X_24428_ _22940_/X _32743_/Q _24432_/S VGND VGND VPWR VPWR _24429_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28196_ _27766_/X _34430_/Q _28214_/S VGND VGND VPWR VPWR _28197_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27147_ _33978_/Q _27146_/X _27156_/S VGND VGND VPWR VPWR _27148_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24359_ _24359_/A VGND VGND VPWR VPWR _32710_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27078_ input6/X VGND VGND VPWR VPWR _27078_/X sky130_fd_sc_hd__buf_4
XFILLER_197_1095 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26029_ _26029_/A VGND VGND VPWR VPWR _33468_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18920_ _34661_/Q _34597_/Q _34533_/Q _34469_/Q _18886_/X _18887_/X VGND VGND VPWR
+ VPWR _18920_/X sky130_fd_sc_hd__mux4_1
XTAP_7130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18851_ _33059_/Q _32035_/Q _35811_/Q _35747_/Q _18672_/X _18673_/X VGND VGND VPWR
+ VPWR _18851_/X sky130_fd_sc_hd__mux4_1
XTAP_6440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17802_ _17552_/X _17798_/X _17801_/X _17557_/X VGND VGND VPWR VPWR _17802_/X sky130_fd_sc_hd__a22o_1
XTAP_6473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18782_ _18597_/X _18780_/X _18781_/X _18600_/X VGND VGND VPWR VPWR _18782_/X sky130_fd_sc_hd__a22o_1
X_15994_ _16063_/A VGND VGND VPWR VPWR _17800_/A sky130_fd_sc_hd__buf_12
XFILLER_227_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17733_ _17559_/X _17729_/X _17732_/X _17562_/X VGND VGND VPWR VPWR _17733_/X sky130_fd_sc_hd__a22o_1
XTAP_5783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29719_ _29719_/A VGND VGND VPWR VPWR _35120_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30991_ _30991_/A VGND VGND VPWR VPWR _35723_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_984 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32730_ _35994_/CLK _32730_/D VGND VGND VPWR VPWR _32730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_932 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17664_ _33155_/Q _36035_/Q _33027_/Q _32963_/Q _17415_/X _17416_/X VGND VGND VPWR
+ VPWR _17664_/X sky130_fd_sc_hd__mux4_1
XFILLER_247_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19403_ _19359_/X _19401_/X _19402_/X _19365_/X VGND VGND VPWR VPWR _19403_/X sky130_fd_sc_hd__a22o_1
XFILLER_91_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16615_ _16292_/X _16613_/X _16614_/X _16295_/X VGND VGND VPWR VPWR _16615_/X sky130_fd_sc_hd__a22o_1
XFILLER_223_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32661_ _36053_/CLK _32661_/D VGND VGND VPWR VPWR _32661_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17595_ _17559_/X _17593_/X _17594_/X _17562_/X VGND VGND VPWR VPWR _17595_/X sky130_fd_sc_hd__a22o_1
XFILLER_245_1030 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34400_ _34593_/CLK _34400_/D VGND VGND VPWR VPWR _34400_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31612_ _31612_/A VGND VGND VPWR VPWR _36017_/D sky130_fd_sc_hd__clkbuf_1
X_19334_ _19014_/X _19332_/X _19333_/X _19018_/X VGND VGND VPWR VPWR _19334_/X sky130_fd_sc_hd__a22o_1
X_35380_ _35698_/CLK _35380_/D VGND VGND VPWR VPWR _35380_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16546_ _35619_/Q _34979_/Q _34339_/Q _33699_/Q _16438_/X _16439_/X VGND VGND VPWR
+ VPWR _16546_/X sky130_fd_sc_hd__mux4_1
X_32592_ _35982_/CLK _32592_/D VGND VGND VPWR VPWR _32592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34331_ _34331_/CLK _34331_/D VGND VGND VPWR VPWR _34331_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_245_1096 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31543_ _27825_/X _35985_/Q _31543_/S VGND VGND VPWR VPWR _31544_/A sky130_fd_sc_hd__mux2_1
X_19265_ _20100_/A VGND VGND VPWR VPWR _19265_/X sky130_fd_sc_hd__clkbuf_4
X_16477_ _35681_/Q _32188_/Q _35553_/Q _35489_/Q _16258_/X _16259_/X VGND VGND VPWR
+ VPWR _16477_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_48_CLK clkbuf_leaf_49_CLK/A VGND VGND VPWR VPWR _35944_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_203_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18216_ _18212_/X _18215_/X _17871_/A VGND VGND VPWR VPWR _18217_/D sky130_fd_sc_hd__o21ba_1
X_34262_ _34647_/CLK _34262_/D VGND VGND VPWR VPWR _34262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31474_ _27723_/X _35952_/Q _31480_/S VGND VGND VPWR VPWR _31475_/A sky130_fd_sc_hd__mux2_1
X_19196_ _19014_/X _19194_/X _19195_/X _19018_/X VGND VGND VPWR VPWR _19196_/X sky130_fd_sc_hd__a22o_1
XFILLER_223_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36001_ _36003_/CLK _36001_/D VGND VGND VPWR VPWR _36001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33213_ _33531_/CLK _33213_/D VGND VGND VPWR VPWR _33213_/Q sky130_fd_sc_hd__dfxtp_1
X_18147_ _33105_/Q _32081_/Q _35857_/Q _35793_/Q _16079_/X _16080_/X VGND VGND VPWR
+ VPWR _18147_/X sky130_fd_sc_hd__mux4_1
X_30425_ _35455_/Q _29457_/X _30441_/S VGND VGND VPWR VPWR _30426_/A sky130_fd_sc_hd__mux2_1
X_34193_ _34193_/CLK _34193_/D VGND VGND VPWR VPWR _34193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_1067 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33144_ _36025_/CLK _33144_/D VGND VGND VPWR VPWR _33144_/Q sky130_fd_sc_hd__dfxtp_1
X_18078_ _17765_/X _18076_/X _18077_/X _17771_/X VGND VGND VPWR VPWR _18078_/X sky130_fd_sc_hd__a22o_1
X_30356_ _30356_/A VGND VGND VPWR VPWR _35422_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_176_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17029_ _32625_/Q _32561_/Q _32497_/Q _35953_/Q _16923_/X _16707_/X VGND VGND VPWR
+ VPWR _17029_/X sky130_fd_sc_hd__mux4_1
XFILLER_217_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30287_ _30335_/S VGND VGND VPWR VPWR _30306_/S sky130_fd_sc_hd__buf_6
X_33075_ _35187_/CLK _33075_/D VGND VGND VPWR VPWR _33075_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20040_ _19720_/X _20038_/X _20039_/X _19724_/X VGND VGND VPWR VPWR _20040_/X sky130_fd_sc_hd__a22o_1
X_32026_ _34007_/CLK _32026_/D VGND VGND VPWR VPWR _32026_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_962 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33977_ _35641_/CLK _33977_/D VGND VGND VPWR VPWR _33977_/Q sky130_fd_sc_hd__dfxtp_1
X_21991_ _21951_/X _21989_/X _21990_/X _21954_/X VGND VGND VPWR VPWR _21991_/X sky130_fd_sc_hd__a22o_1
XFILLER_6_1276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35716_ _35716_/CLK _35716_/D VGND VGND VPWR VPWR _35716_/Q sky130_fd_sc_hd__dfxtp_1
X_23730_ _22918_/X _32352_/Q _23748_/S VGND VGND VPWR VPWR _23731_/A sky130_fd_sc_hd__mux2_1
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20942_ _20691_/X _20940_/X _20941_/X _20701_/X VGND VGND VPWR VPWR _20942_/X sky130_fd_sc_hd__a22o_1
X_32928_ _36003_/CLK _32928_/D VGND VGND VPWR VPWR _32928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35647_ _36096_/CLK _35647_/D VGND VGND VPWR VPWR _35647_/Q sky130_fd_sc_hd__dfxtp_1
X_23661_ _23021_/X _32321_/Q _23673_/S VGND VGND VPWR VPWR _23662_/A sky130_fd_sc_hd__mux2_1
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20873_ _20869_/X _20872_/X _20704_/X VGND VGND VPWR VPWR _20874_/D sky130_fd_sc_hd__o21ba_1
X_32859_ _35668_/CLK _32859_/D VGND VGND VPWR VPWR _32859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25400_ _25400_/A VGND VGND VPWR VPWR _33171_/D sky130_fd_sc_hd__clkbuf_1
X_22612_ _33421_/Q _33357_/Q _33293_/Q _33229_/Q _22433_/X _22434_/X VGND VGND VPWR
+ VPWR _22612_/X sky130_fd_sc_hd__mux4_1
XFILLER_228_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26380_ _33634_/Q _23268_/X _26394_/S VGND VGND VPWR VPWR _26381_/A sky130_fd_sc_hd__mux2_1
X_23592_ _22918_/X _32288_/Q _23610_/S VGND VGND VPWR VPWR _23593_/A sky130_fd_sc_hd__mux2_1
X_35578_ _35581_/CLK _35578_/D VGND VGND VPWR VPWR _35578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25331_ _25331_/A VGND VGND VPWR VPWR _33138_/D sky130_fd_sc_hd__clkbuf_1
X_22543_ _33675_/Q _33611_/Q _33547_/Q _33483_/Q _22506_/X _22507_/X VGND VGND VPWR
+ VPWR _22543_/X sky130_fd_sc_hd__mux4_1
X_34529_ _35297_/CLK _34529_/D VGND VGND VPWR VPWR _34529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_39_CLK clkbuf_6_7__f_CLK/X VGND VGND VPWR VPWR _35939_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_202_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28050_ _34361_/Q _27143_/X _28058_/S VGND VGND VPWR VPWR _28051_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25262_ _25262_/A VGND VGND VPWR VPWR _33106_/D sky130_fd_sc_hd__clkbuf_1
X_22474_ _22474_/A VGND VGND VPWR VPWR _36232_/D sky130_fd_sc_hd__clkbuf_1
X_27001_ _27001_/A VGND VGND VPWR VPWR _33926_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24213_ _24213_/A VGND VGND VPWR VPWR _32642_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21425_ _21306_/X _21423_/X _21424_/X _21312_/X VGND VGND VPWR VPWR _21425_/X sky130_fd_sc_hd__a22o_1
XFILLER_212_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25193_ _25193_/A VGND VGND VPWR VPWR _33073_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24144_ _24144_/A VGND VGND VPWR VPWR _32609_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21356_ _35625_/Q _34985_/Q _34345_/Q _33705_/Q _21038_/X _21039_/X VGND VGND VPWR
+ VPWR _21356_/X sky130_fd_sc_hd__mux4_1
XFILLER_120_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20307_ _20307_/A _20307_/B _20307_/C _20307_/D VGND VGND VPWR VPWR _20308_/A sky130_fd_sc_hd__or4_1
X_24075_ _24075_/A VGND VGND VPWR VPWR _32578_/D sky130_fd_sc_hd__clkbuf_1
X_28952_ _34787_/Q _27075_/X _28964_/S VGND VGND VPWR VPWR _28953_/A sky130_fd_sc_hd__mux2_1
X_21287_ _33063_/Q _32039_/Q _35815_/Q _35751_/Q _20972_/X _20973_/X VGND VGND VPWR
+ VPWR _21287_/X sky130_fd_sc_hd__mux4_1
XFILLER_104_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_831 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23026_ _23026_/A VGND VGND VPWR VPWR _32066_/D sky130_fd_sc_hd__clkbuf_1
X_27903_ _27903_/A VGND VGND VPWR VPWR _34291_/D sky130_fd_sc_hd__clkbuf_1
X_20238_ _34954_/Q _34890_/Q _34826_/Q _34762_/Q _20166_/X _20167_/X VGND VGND VPWR
+ VPWR _20238_/X sky130_fd_sc_hd__mux4_1
X_28883_ _28883_/A VGND VGND VPWR VPWR _34754_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1052 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27834_ input59/X VGND VGND VPWR VPWR _27834_/X sky130_fd_sc_hd__clkbuf_4
XTAP_5035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20169_ _20169_/A VGND VGND VPWR VPWR _20169_/X sky130_fd_sc_hd__clkbuf_4
XTAP_5046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27765_ _27765_/A VGND VGND VPWR VPWR _34237_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24977_ _24976_/X _32975_/Q _24983_/S VGND VGND VPWR VPWR _24978_/A sky130_fd_sc_hd__mux2_1
XTAP_4356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29504_ _35022_/Q _29503_/X _29513_/S VGND VGND VPWR VPWR _29505_/A sky130_fd_sc_hd__mux2_1
XTAP_3633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26716_ _33791_/Q _23426_/X _26732_/S VGND VGND VPWR VPWR _26717_/A sky130_fd_sc_hd__mux2_1
XTAP_4389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23928_ _23928_/A VGND VGND VPWR VPWR _32509_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27696_ _27695_/X _34215_/Q _27702_/S VGND VGND VPWR VPWR _27697_/A sky130_fd_sc_hd__mux2_1
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29435_ input28/X VGND VGND VPWR VPWR _29435_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23859_ _23859_/A VGND VGND VPWR VPWR _32476_/D sky130_fd_sc_hd__clkbuf_1
X_26647_ _26647_/A VGND VGND VPWR VPWR _33758_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16400_ _16361_/X _16398_/X _16399_/X _16365_/X VGND VGND VPWR VPWR _16400_/X sky130_fd_sc_hd__a22o_1
XTAP_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17380_ _17206_/X _17376_/X _17379_/X _17209_/X VGND VGND VPWR VPWR _17380_/X sky130_fd_sc_hd__a22o_1
X_29366_ _29366_/A VGND VGND VPWR VPWR _34977_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26578_ _26578_/A VGND VGND VPWR VPWR _33727_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_242_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16331_ _35613_/Q _34973_/Q _34333_/Q _33693_/Q _16053_/X _16055_/X VGND VGND VPWR
+ VPWR _16331_/X sky130_fd_sc_hd__mux4_1
XFILLER_111_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28317_ _28317_/A VGND VGND VPWR VPWR _34487_/D sky130_fd_sc_hd__clkbuf_1
X_25529_ _25529_/A VGND VGND VPWR VPWR _33231_/D sky130_fd_sc_hd__clkbuf_1
X_29297_ _34951_/Q _27186_/X _29297_/S VGND VGND VPWR VPWR _29298_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16262_ _16048_/X _16260_/X _16261_/X _16058_/X VGND VGND VPWR VPWR _16262_/X sky130_fd_sc_hd__a22o_1
X_19050_ _19006_/X _19048_/X _19049_/X _19012_/X VGND VGND VPWR VPWR _19050_/X sky130_fd_sc_hd__a22o_1
X_28248_ _28248_/A VGND VGND VPWR VPWR _34454_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18001_ _35212_/Q _35148_/Q _35084_/Q _32268_/Q _17716_/X _17717_/X VGND VGND VPWR
+ VPWR _18001_/X sky130_fd_sc_hd__mux4_1
XFILLER_199_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_923 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16193_ _35609_/Q _34969_/Q _34329_/Q _33689_/Q _16053_/X _16055_/X VGND VGND VPWR
+ VPWR _16193_/X sky130_fd_sc_hd__mux4_1
XFILLER_103_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28179_ _27742_/X _34422_/Q _28193_/S VGND VGND VPWR VPWR _28180_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30210_ _35353_/Q _29339_/X _30222_/S VGND VGND VPWR VPWR _30211_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31190_ _31190_/A VGND VGND VPWR VPWR _35817_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30141_ _30141_/A VGND VGND VPWR VPWR _35320_/D sky130_fd_sc_hd__clkbuf_1
X_19952_ _19811_/X _19950_/X _19951_/X _19816_/X VGND VGND VPWR VPWR _19952_/X sky130_fd_sc_hd__a22o_1
XFILLER_5_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18903_ _18899_/X _18902_/X _18726_/X VGND VGND VPWR VPWR _18927_/A sky130_fd_sc_hd__o21ba_1
X_30072_ _30072_/A VGND VGND VPWR VPWR _35287_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_206_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19883_ _20236_/A VGND VGND VPWR VPWR _19883_/X sky130_fd_sc_hd__buf_4
XFILLER_171_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33900_ _34093_/CLK _33900_/D VGND VGND VPWR VPWR _33900_/Q sky130_fd_sc_hd__dfxtp_1
X_18834_ _33379_/Q _33315_/Q _33251_/Q _33187_/Q _18721_/X _18722_/X VGND VGND VPWR
+ VPWR _18834_/X sky130_fd_sc_hd__mux4_1
X_34880_ _34945_/CLK _34880_/D VGND VGND VPWR VPWR _34880_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33831_ _33897_/CLK _33831_/D VGND VGND VPWR VPWR _33831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18765_ _18440_/X _18763_/X _18764_/X _18445_/X VGND VGND VPWR VPWR _18765_/X sky130_fd_sc_hd__a22o_1
XTAP_5580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_222_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17716_ _17716_/A VGND VGND VPWR VPWR _17716_/X sky130_fd_sc_hd__clkbuf_8
X_33762_ _36066_/CLK _33762_/D VGND VGND VPWR VPWR _33762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_247_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30974_ _30974_/A VGND VGND VPWR VPWR _35715_/D sky130_fd_sc_hd__clkbuf_1
X_18696_ _33119_/Q _35999_/Q _32991_/Q _32927_/Q _18656_/X _18657_/X VGND VGND VPWR
+ VPWR _18696_/X sky130_fd_sc_hd__mux4_1
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35501_ _35693_/CLK _35501_/D VGND VGND VPWR VPWR _35501_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32713_ _32907_/CLK _32713_/D VGND VGND VPWR VPWR _32713_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17647_ _34690_/Q _34626_/Q _34562_/Q _34498_/Q _17645_/X _17646_/X VGND VGND VPWR
+ VPWR _17647_/X sky130_fd_sc_hd__mux4_1
XFILLER_224_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33693_ _35613_/CLK _33693_/D VGND VGND VPWR VPWR _33693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35432_ _35434_/CLK _35432_/D VGND VGND VPWR VPWR _35432_/Q sky130_fd_sc_hd__dfxtp_1
X_32644_ _36038_/CLK _32644_/D VGND VGND VPWR VPWR _32644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_1180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17578_ _17574_/X _17577_/X _17504_/X VGND VGND VPWR VPWR _17588_/C sky130_fd_sc_hd__o21ba_1
XFILLER_205_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19317_ _19313_/X _19316_/X _19112_/X VGND VGND VPWR VPWR _19318_/D sky130_fd_sc_hd__o21ba_1
XFILLER_182_1172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35363_ _35814_/CLK _35363_/D VGND VGND VPWR VPWR _35363_/Q sky130_fd_sc_hd__dfxtp_1
X_16529_ _16529_/A _16529_/B _16529_/C _16529_/D VGND VGND VPWR VPWR _16530_/A sky130_fd_sc_hd__or4_2
X_32575_ _32575_/CLK _32575_/D VGND VGND VPWR VPWR _32575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34314_ _36173_/CLK _34314_/D VGND VGND VPWR VPWR _34314_/Q sky130_fd_sc_hd__dfxtp_1
X_31526_ _31526_/A VGND VGND VPWR VPWR _35976_/D sky130_fd_sc_hd__clkbuf_1
X_19248_ _19248_/A _19248_/B _19248_/C _19248_/D VGND VGND VPWR VPWR _19249_/A sky130_fd_sc_hd__or4_4
XFILLER_220_996 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35294_ _35743_/CLK _35294_/D VGND VGND VPWR VPWR _35294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34245_ _36165_/CLK _34245_/D VGND VGND VPWR VPWR _34245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19179_ _34924_/Q _34860_/Q _34796_/Q _34732_/Q _19107_/X _19108_/X VGND VGND VPWR
+ VPWR _19179_/X sky130_fd_sc_hd__mux4_1
X_31457_ _27698_/X _35944_/Q _31459_/S VGND VGND VPWR VPWR _31458_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21210_ _21206_/X _21209_/X _21034_/X _21035_/X VGND VGND VPWR VPWR _21227_/B sky130_fd_sc_hd__o211a_1
X_30408_ _35447_/Q _29432_/X _30420_/S VGND VGND VPWR VPWR _30409_/A sky130_fd_sc_hd__mux2_1
X_22190_ _33665_/Q _33601_/Q _33537_/Q _33473_/Q _22153_/X _22154_/X VGND VGND VPWR
+ VPWR _22190_/X sky130_fd_sc_hd__mux4_1
X_34176_ _36159_/CLK _34176_/D VGND VGND VPWR VPWR _34176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31388_ _31388_/A VGND VGND VPWR VPWR _35911_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_5_5_0_CLK clkbuf_5_7_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_5_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_219_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33127_ _35943_/CLK _33127_/D VGND VGND VPWR VPWR _33127_/Q sky130_fd_sc_hd__dfxtp_1
X_21141_ _32099_/Q _32291_/Q _32355_/Q _35875_/Q _20821_/X _20962_/X VGND VGND VPWR
+ VPWR _21141_/X sky130_fd_sc_hd__mux4_1
X_30339_ _35414_/Q _29328_/X _30357_/S VGND VGND VPWR VPWR _30340_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21072_ _20953_/X _21070_/X _21071_/X _20959_/X VGND VGND VPWR VPWR _21072_/X sky130_fd_sc_hd__a22o_1
XFILLER_116_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33058_ _35812_/CLK _33058_/D VGND VGND VPWR VPWR _33058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20023_ _20019_/X _20022_/X _19818_/X VGND VGND VPWR VPWR _20024_/D sky130_fd_sc_hd__o21ba_1
X_24900_ _24899_/X _32950_/Q _24921_/S VGND VGND VPWR VPWR _24901_/A sky130_fd_sc_hd__mux2_1
X_32009_ _36209_/CLK _32009_/D VGND VGND VPWR VPWR _32009_/Q sky130_fd_sc_hd__dfxtp_1
X_25880_ _25880_/A VGND VGND VPWR VPWR _33397_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_246_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_1422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24831_ _24995_/S VGND VGND VPWR VPWR _24859_/S sky130_fd_sc_hd__buf_4
XFILLER_80_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24762_ _24762_/A VGND VGND VPWR VPWR _32901_/D sky130_fd_sc_hd__clkbuf_1
X_27550_ _34155_/Q _27100_/X _27566_/S VGND VGND VPWR VPWR _27551_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21974_ _34171_/Q _34107_/Q _34043_/Q _33979_/Q _21693_/X _21694_/X VGND VGND VPWR
+ VPWR _21974_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23713_ _22894_/X _32344_/Q _23727_/S VGND VGND VPWR VPWR _23714_/A sky130_fd_sc_hd__mux2_1
X_26501_ _24815_/X _33691_/Q _26509_/S VGND VGND VPWR VPWR _26502_/A sky130_fd_sc_hd__mux2_1
X_27481_ _27481_/A VGND VGND VPWR VPWR _34122_/D sky130_fd_sc_hd__clkbuf_1
X_20925_ _20618_/X _20923_/X _20924_/X _20627_/X VGND VGND VPWR VPWR _20925_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24693_ _24693_/A VGND VGND VPWR VPWR _32868_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29220_ _34914_/Q _27072_/X _29234_/S VGND VGND VPWR VPWR _29221_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26432_ _33659_/Q _23411_/X _26436_/S VGND VGND VPWR VPWR _26433_/A sky130_fd_sc_hd__mux2_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23644_ _22996_/X _32313_/Q _23652_/S VGND VGND VPWR VPWR _23645_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20856_ _20630_/X _20854_/X _20855_/X _20641_/X VGND VGND VPWR VPWR _20856_/X sky130_fd_sc_hd__a22o_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29151_ _29151_/A VGND VGND VPWR VPWR _34881_/D sky130_fd_sc_hd__clkbuf_1
X_26363_ _33626_/Q _23243_/X _26373_/S VGND VGND VPWR VPWR _26364_/A sky130_fd_sc_hd__mux2_1
X_23575_ _22894_/X _32280_/Q _23589_/S VGND VGND VPWR VPWR _23576_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20787_ _20618_/X _20785_/X _20786_/X _20627_/X VGND VGND VPWR VPWR _20787_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28102_ _34386_/Q _27220_/X _28108_/S VGND VGND VPWR VPWR _28103_/A sky130_fd_sc_hd__mux2_1
X_25314_ _33130_/Q _23292_/X _25332_/S VGND VGND VPWR VPWR _25315_/A sky130_fd_sc_hd__mux2_1
X_22526_ _35658_/Q _35018_/Q _34378_/Q _33738_/Q _22450_/X _22451_/X VGND VGND VPWR
+ VPWR _22526_/X sky130_fd_sc_hd__mux4_1
XFILLER_22_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26294_ _24911_/X _33594_/Q _26300_/S VGND VGND VPWR VPWR _26295_/A sky130_fd_sc_hd__mux2_1
X_29082_ _29082_/A VGND VGND VPWR VPWR _34848_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_241_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25245_ _33098_/Q _23463_/X _25259_/S VGND VGND VPWR VPWR _25246_/A sky130_fd_sc_hd__mux2_1
X_28033_ _34353_/Q _27118_/X _28037_/S VGND VGND VPWR VPWR _28034_/A sky130_fd_sc_hd__mux2_1
XFILLER_202_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22457_ _22457_/A VGND VGND VPWR VPWR _22457_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21408_ _21761_/A VGND VGND VPWR VPWR _21408_/X sky130_fd_sc_hd__clkbuf_4
X_25176_ _25176_/A VGND VGND VPWR VPWR _33065_/D sky130_fd_sc_hd__clkbuf_1
X_22388_ _22382_/X _22387_/X _22104_/X VGND VGND VPWR VPWR _22396_/C sky130_fd_sc_hd__o21ba_1
XFILLER_157_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24127_ _24127_/A VGND VGND VPWR VPWR _32601_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21339_ _33641_/Q _33577_/Q _33513_/Q _33449_/Q _21094_/X _21095_/X VGND VGND VPWR
+ VPWR _21339_/X sky130_fd_sc_hd__mux4_1
X_29984_ _35246_/Q _29404_/X _29994_/S VGND VGND VPWR VPWR _29985_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28935_ _34779_/Q _27050_/X _28943_/S VGND VGND VPWR VPWR _28936_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24058_ _24058_/A VGND VGND VPWR VPWR _32570_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23009_ _23008_/X _32061_/Q _23009_/S VGND VGND VPWR VPWR _23010_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28866_ _28866_/A VGND VGND VPWR VPWR _34746_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16880_ _16805_/X _16878_/X _16879_/X _16810_/X VGND VGND VPWR VPWR _16880_/X sky130_fd_sc_hd__a22o_1
XFILLER_77_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27817_ _27816_/X _34254_/Q _27826_/S VGND VGND VPWR VPWR _27818_/A sky130_fd_sc_hd__mux2_1
XTAP_4120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28797_ _28797_/A VGND VGND VPWR VPWR _34713_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18550_ _18546_/X _18549_/X _18315_/X VGND VGND VPWR VPWR _18574_/A sky130_fd_sc_hd__o21ba_1
XTAP_4164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27748_ input28/X VGND VGND VPWR VPWR _27748_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17501_ _35454_/Q _35390_/Q _35326_/Q _35262_/Q _17254_/X _17255_/X VGND VGND VPWR
+ VPWR _17501_/X sky130_fd_sc_hd__mux4_1
XFILLER_73_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_233_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18481_ _33369_/Q _33305_/Q _33241_/Q _33177_/Q _18302_/X _18303_/X VGND VGND VPWR
+ VPWR _18481_/X sky130_fd_sc_hd__mux4_1
XTAP_3474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27679_ _27679_/A VGND VGND VPWR VPWR _34209_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_935 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29418_ _29418_/A VGND VGND VPWR VPWR _34994_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17432_ _17936_/A VGND VGND VPWR VPWR _17432_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_221_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30690_ _35581_/Q _29450_/X _30690_/S VGND VGND VPWR VPWR _30691_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_1410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29349_ _34972_/Q _29348_/X _29358_/S VGND VGND VPWR VPWR _29350_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17363_ _17716_/A VGND VGND VPWR VPWR _17363_/X sky130_fd_sc_hd__buf_6
XFILLER_159_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19102_ _35178_/Q _35114_/Q _35050_/Q _32170_/Q _18957_/X _18958_/X VGND VGND VPWR
+ VPWR _19102_/X sky130_fd_sc_hd__mux4_1
XFILLER_92_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16314_ _33629_/Q _33565_/Q _33501_/Q _33437_/Q _16141_/X _16142_/X VGND VGND VPWR
+ VPWR _16314_/X sky130_fd_sc_hd__mux4_1
XFILLER_140_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32360_ _32873_/CLK _32360_/D VGND VGND VPWR VPWR _32360_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17294_ _34680_/Q _34616_/Q _34552_/Q _34488_/Q _17292_/X _17293_/X VGND VGND VPWR
+ VPWR _17294_/X sky130_fd_sc_hd__mux4_1
X_31311_ _31311_/A VGND VGND VPWR VPWR _35874_/D sky130_fd_sc_hd__clkbuf_1
X_19033_ _34408_/Q _36136_/Q _34280_/Q _34216_/Q _18823_/X _18824_/X VGND VGND VPWR
+ VPWR _19033_/X sky130_fd_sc_hd__mux4_1
X_16245_ _34139_/Q _34075_/Q _34011_/Q _33947_/Q _16009_/X _16011_/X VGND VGND VPWR
+ VPWR _16245_/X sky130_fd_sc_hd__mux4_1
XFILLER_12_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32291_ _32871_/CLK _32291_/D VGND VGND VPWR VPWR _32291_/Q sky130_fd_sc_hd__dfxtp_1
X_34030_ _35630_/CLK _34030_/D VGND VGND VPWR VPWR _34030_/Q sky130_fd_sc_hd__dfxtp_1
X_31242_ _27779_/X _35842_/Q _31252_/S VGND VGND VPWR VPWR _31243_/A sky130_fd_sc_hd__mux2_1
X_16176_ _16176_/A _16176_/B _16176_/C _16176_/D VGND VGND VPWR VPWR _16177_/A sky130_fd_sc_hd__or4_1
XFILLER_217_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput106 _31982_/Q VGND VGND VPWR VPWR D1[24] sky130_fd_sc_hd__buf_2
XFILLER_103_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput117 _31992_/Q VGND VGND VPWR VPWR D1[34] sky130_fd_sc_hd__buf_2
Xoutput128 _32002_/Q VGND VGND VPWR VPWR D1[44] sky130_fd_sc_hd__buf_2
X_31173_ _27677_/X _35809_/Q _31189_/S VGND VGND VPWR VPWR _31174_/A sky130_fd_sc_hd__mux2_1
Xoutput139 _32012_/Q VGND VGND VPWR VPWR D1[54] sky130_fd_sc_hd__buf_2
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19935_ _32898_/Q _32834_/Q _32770_/Q _32706_/Q _19646_/X _19647_/X VGND VGND VPWR
+ VPWR _19935_/X sky130_fd_sc_hd__mux4_1
X_30124_ _30124_/A VGND VGND VPWR VPWR _35312_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35981_ _35983_/CLK _35981_/D VGND VGND VPWR VPWR _35981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30055_ _35280_/Q _29509_/X _30057_/S VGND VGND VPWR VPWR _30056_/A sky130_fd_sc_hd__mux2_1
X_34932_ _35828_/CLK _34932_/D VGND VGND VPWR VPWR _34932_/Q sky130_fd_sc_hd__dfxtp_1
X_19866_ _33152_/Q _36032_/Q _33024_/Q _32960_/Q _19715_/X _19716_/X VGND VGND VPWR
+ VPWR _19866_/X sky130_fd_sc_hd__mux4_1
XFILLER_214_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18817_ _33058_/Q _32034_/Q _35810_/Q _35746_/Q _18672_/X _18673_/X VGND VGND VPWR
+ VPWR _18817_/X sky130_fd_sc_hd__mux4_1
XFILLER_233_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34863_ _35438_/CLK _34863_/D VGND VGND VPWR VPWR _34863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19797_ _20150_/A VGND VGND VPWR VPWR _19797_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_110_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33814_ _36054_/CLK _33814_/D VGND VGND VPWR VPWR _33814_/Q sky130_fd_sc_hd__dfxtp_1
X_18748_ _34656_/Q _34592_/Q _34528_/Q _34464_/Q _18533_/X _18534_/X VGND VGND VPWR
+ VPWR _18748_/X sky130_fd_sc_hd__mux4_1
XFILLER_23_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34794_ _35692_/CLK _34794_/D VGND VGND VPWR VPWR _34794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33745_ _35728_/CLK _33745_/D VGND VGND VPWR VPWR _33745_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18679_ _18378_/X _18677_/X _18678_/X _18388_/X VGND VGND VPWR VPWR _18679_/X sky130_fd_sc_hd__a22o_1
X_30957_ _30957_/A VGND VGND VPWR VPWR _35707_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_1106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20710_ _20581_/X _20708_/X _20709_/X _20591_/X VGND VGND VPWR VPWR _20710_/X sky130_fd_sc_hd__a22o_1
XFILLER_24_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33676_ _33934_/CLK _33676_/D VGND VGND VPWR VPWR _33676_/Q sky130_fd_sc_hd__dfxtp_1
X_21690_ _21690_/A _21690_/B _21690_/C _21690_/D VGND VGND VPWR VPWR _21691_/A sky130_fd_sc_hd__or4_1
XFILLER_212_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30888_ _30888_/A VGND VGND VPWR VPWR _35674_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35415_ _36118_/CLK _35415_/D VGND VGND VPWR VPWR _35415_/Q sky130_fd_sc_hd__dfxtp_1
X_20641_ _22515_/A VGND VGND VPWR VPWR _20641_/X sky130_fd_sc_hd__clkbuf_4
X_32627_ _36019_/CLK _32627_/D VGND VGND VPWR VPWR _32627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35346_ _35858_/CLK _35346_/D VGND VGND VPWR VPWR _35346_/Q sky130_fd_sc_hd__dfxtp_1
X_23360_ _23360_/A VGND VGND VPWR VPWR _32196_/D sky130_fd_sc_hd__clkbuf_1
X_20572_ _18348_/X _20570_/X _20571_/X _18358_/X VGND VGND VPWR VPWR _20572_/X sky130_fd_sc_hd__a22o_1
X_32558_ _35951_/CLK _32558_/D VGND VGND VPWR VPWR _32558_/Q sky130_fd_sc_hd__dfxtp_1
X_22311_ _33092_/Q _32068_/Q _35844_/Q _35780_/Q _22031_/X _22032_/X VGND VGND VPWR
+ VPWR _22311_/X sky130_fd_sc_hd__mux4_1
X_31509_ _31509_/A VGND VGND VPWR VPWR _35968_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35277_ _35471_/CLK _35277_/D VGND VGND VPWR VPWR _35277_/Q sky130_fd_sc_hd__dfxtp_1
X_23291_ _23291_/A VGND VGND VPWR VPWR _32169_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_1016 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32489_ _35944_/CLK _32489_/D VGND VGND VPWR VPWR _32489_/Q sky130_fd_sc_hd__dfxtp_1
X_25030_ _24846_/X _32997_/Q _25038_/S VGND VGND VPWR VPWR _25031_/A sky130_fd_sc_hd__mux2_1
X_22242_ _33090_/Q _32066_/Q _35842_/Q _35778_/Q _22031_/X _22032_/X VGND VGND VPWR
+ VPWR _22242_/X sky130_fd_sc_hd__mux4_1
X_34228_ _35187_/CLK _34228_/D VGND VGND VPWR VPWR _34228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22173_ _35648_/Q _35008_/Q _34368_/Q _33728_/Q _22097_/X _22098_/X VGND VGND VPWR
+ VPWR _22173_/X sky130_fd_sc_hd__mux4_1
X_34159_ _34991_/CLK _34159_/D VGND VGND VPWR VPWR _34159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21124_ _21477_/A VGND VGND VPWR VPWR _21124_/X sky130_fd_sc_hd__buf_4
XFILLER_121_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26981_ _33917_/Q _23417_/X _26981_/S VGND VGND VPWR VPWR _26982_/A sky130_fd_sc_hd__mux2_1
XFILLER_236_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28720_ _34678_/Q _27134_/X _28734_/S VGND VGND VPWR VPWR _28721_/A sky130_fd_sc_hd__mux2_1
X_25932_ _25932_/A VGND VGND VPWR VPWR _33422_/D sky130_fd_sc_hd__clkbuf_1
X_21055_ _21761_/A VGND VGND VPWR VPWR _21055_/X sky130_fd_sc_hd__clkbuf_4
X_20006_ _35652_/Q _35012_/Q _34372_/Q _33732_/Q _19797_/X _19798_/X VGND VGND VPWR
+ VPWR _20006_/X sky130_fd_sc_hd__mux4_1
XFILLER_219_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28651_ _28651_/A VGND VGND VPWR VPWR _28784_/S sky130_fd_sc_hd__buf_12
XFILLER_143_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25863_ _25863_/A VGND VGND VPWR VPWR _33389_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27602_ _34180_/Q _27177_/X _27608_/S VGND VGND VPWR VPWR _27603_/A sky130_fd_sc_hd__mux2_1
XFILLER_228_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24814_ _24814_/A VGND VGND VPWR VPWR _32922_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_246_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28582_ _27739_/X _34613_/Q _28598_/S VGND VGND VPWR VPWR _28583_/A sky130_fd_sc_hd__mux2_1
X_25794_ _24970_/X _33357_/Q _25802_/S VGND VGND VPWR VPWR _25795_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27533_ _34147_/Q _27075_/X _27545_/S VGND VGND VPWR VPWR _27534_/A sky130_fd_sc_hd__mux2_1
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24745_ _24745_/A VGND VGND VPWR VPWR _32893_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21957_ _35450_/Q _35386_/Q _35322_/Q _35258_/Q _21854_/X _21855_/X VGND VGND VPWR
+ VPWR _21957_/X sky130_fd_sc_hd__mux4_1
XFILLER_215_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_270_CLK clkbuf_6_60__f_CLK/X VGND VGND VPWR VPWR _35717_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20908_ _34396_/Q _36124_/Q _34268_/Q _34204_/Q _20770_/X _20771_/X VGND VGND VPWR
+ VPWR _20908_/X sky130_fd_sc_hd__mux4_1
XFILLER_27_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27464_ _27464_/A VGND VGND VPWR VPWR _34114_/D sky130_fd_sc_hd__clkbuf_1
X_24676_ _24676_/A VGND VGND VPWR VPWR _32860_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_587 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21888_ _35448_/Q _35384_/Q _35320_/Q _35256_/Q _21854_/X _21855_/X VGND VGND VPWR
+ VPWR _21888_/X sky130_fd_sc_hd__mux4_1
XFILLER_230_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29203_ _34906_/Q _27047_/X _29213_/S VGND VGND VPWR VPWR _29204_/A sky130_fd_sc_hd__mux2_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26415_ _33651_/Q _23384_/X _26415_/S VGND VGND VPWR VPWR _26416_/A sky130_fd_sc_hd__mux2_1
X_23627_ _22971_/X _32305_/Q _23631_/S VGND VGND VPWR VPWR _23628_/A sky130_fd_sc_hd__mux2_1
X_20839_ _34906_/Q _34842_/Q _34778_/Q _34714_/Q _20696_/X _20698_/X VGND VGND VPWR
+ VPWR _20839_/X sky130_fd_sc_hd__mux4_1
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27395_ _27395_/A VGND VGND VPWR VPWR _34081_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_10 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29134_ _29134_/A VGND VGND VPWR VPWR _34873_/D sky130_fd_sc_hd__clkbuf_1
X_26346_ _24988_/X _33619_/Q _26350_/S VGND VGND VPWR VPWR _26347_/A sky130_fd_sc_hd__mux2_1
X_23558_ _23558_/A VGND VGND VPWR VPWR _32273_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22509_ _34186_/Q _34122_/Q _34058_/Q _33994_/Q _22399_/X _22400_/X VGND VGND VPWR
+ VPWR _22509_/X sky130_fd_sc_hd__mux4_1
XFILLER_156_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput19 DW[26] VGND VGND VPWR VPWR input19/X sky130_fd_sc_hd__clkbuf_8
X_29065_ _29065_/A VGND VGND VPWR VPWR _34840_/D sky130_fd_sc_hd__clkbuf_1
X_26277_ _24886_/X _33586_/Q _26279_/S VGND VGND VPWR VPWR _26278_/A sky130_fd_sc_hd__mux2_1
X_23489_ _23489_/A VGND VGND VPWR VPWR _32241_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16030_ _17912_/A VGND VGND VPWR VPWR _16030_/X sky130_fd_sc_hd__buf_4
X_28016_ _34345_/Q _27093_/X _28016_/S VGND VGND VPWR VPWR _28017_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25228_ _33090_/Q _23435_/X _25238_/S VGND VGND VPWR VPWR _25229_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25159_ _33057_/Q _23265_/X _25175_/S VGND VGND VPWR VPWR _25160_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17981_ _17977_/X _17980_/X _17838_/X VGND VGND VPWR VPWR _18007_/A sky130_fd_sc_hd__o21ba_2
X_29967_ _35238_/Q _29379_/X _29973_/S VGND VGND VPWR VPWR _29968_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19720_ _20212_/A VGND VGND VPWR VPWR _19720_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_111_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28918_ _28918_/A VGND VGND VPWR VPWR _34771_/D sky130_fd_sc_hd__clkbuf_1
X_16932_ _35694_/Q _32202_/Q _35566_/Q _35502_/Q _16611_/X _16612_/X VGND VGND VPWR
+ VPWR _16932_/X sky130_fd_sc_hd__mux4_1
XFILLER_2_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29898_ _29898_/A VGND VGND VPWR VPWR _35205_/D sky130_fd_sc_hd__clkbuf_1
X_19651_ _20159_/A VGND VGND VPWR VPWR _19651_/X sky130_fd_sc_hd__buf_6
X_16863_ _32876_/Q _32812_/Q _32748_/Q _32684_/Q _16640_/X _16641_/X VGND VGND VPWR
+ VPWR _16863_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_718 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28849_ _28849_/A VGND VGND VPWR VPWR _34738_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18602_ _18596_/X _18601_/X _18375_/X VGND VGND VPWR VPWR _18612_/C sky130_fd_sc_hd__o21ba_1
XFILLER_111_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31860_ _23283_/X _36135_/Q _31864_/S VGND VGND VPWR VPWR _31861_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19582_ _32888_/Q _32824_/Q _32760_/Q _32696_/Q _19293_/X _19294_/X VGND VGND VPWR
+ VPWR _19582_/X sky130_fd_sc_hd__mux4_1
XFILLER_219_882 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16794_ _16645_/X _16790_/X _16793_/X _16648_/X VGND VGND VPWR VPWR _16794_/X sky130_fd_sc_hd__a22o_1
XFILLER_206_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18533_ _20298_/A VGND VGND VPWR VPWR _18533_/X sky130_fd_sc_hd__buf_6
X_30811_ _35638_/Q input26/X _30825_/S VGND VGND VPWR VPWR _30812_/A sky130_fd_sc_hd__mux2_1
XFILLER_218_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31791_ _31791_/A VGND VGND VPWR VPWR _36102_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_261_CLK clkbuf_6_62__f_CLK/X VGND VGND VPWR VPWR _36102_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33530_ _33913_/CLK _33530_/D VGND VGND VPWR VPWR _33530_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18464_ _33048_/Q _32024_/Q _35800_/Q _35736_/Q _18367_/X _18369_/X VGND VGND VPWR
+ VPWR _18464_/X sky130_fd_sc_hd__mux4_1
X_30742_ _31147_/A _30877_/B VGND VGND VPWR VPWR _30875_/S sky130_fd_sc_hd__nor2_8
XFILLER_248_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17415_ _17986_/A VGND VGND VPWR VPWR _17415_/X sky130_fd_sc_hd__buf_6
XFILLER_60_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33461_ _36085_/CLK _33461_/D VGND VGND VPWR VPWR _33461_/Q sky130_fd_sc_hd__dfxtp_1
X_18395_ _34390_/Q _36118_/Q _34262_/Q _34198_/Q _18392_/X _18394_/X VGND VGND VPWR
+ VPWR _18395_/X sky130_fd_sc_hd__mux4_1
XFILLER_21_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30673_ _30673_/A VGND VGND VPWR VPWR _35572_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35200_ _35715_/CLK _35200_/D VGND VGND VPWR VPWR _35200_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32412_ _34151_/CLK _32412_/D VGND VGND VPWR VPWR _32412_/Q sky130_fd_sc_hd__dfxtp_1
X_36180_ _36180_/CLK _36180_/D VGND VGND VPWR VPWR _36180_/Q sky130_fd_sc_hd__dfxtp_1
X_17346_ _17833_/A VGND VGND VPWR VPWR _17346_/X sky130_fd_sc_hd__buf_4
XFILLER_92_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33392_ _33904_/CLK _33392_/D VGND VGND VPWR VPWR _33392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35131_ _35197_/CLK _35131_/D VGND VGND VPWR VPWR _35131_/Q sky130_fd_sc_hd__dfxtp_1
X_32343_ _35863_/CLK _32343_/D VGND VGND VPWR VPWR _32343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17277_ _32632_/Q _32568_/Q _32504_/Q _35960_/Q _17276_/X _17060_/X VGND VGND VPWR
+ VPWR _17277_/X sky130_fd_sc_hd__mux4_1
X_19016_ _32104_/Q _32296_/Q _32360_/Q _35880_/Q _18874_/X _19015_/X VGND VGND VPWR
+ VPWR _19016_/X sky130_fd_sc_hd__mux4_1
X_16228_ _16048_/X _16226_/X _16227_/X _16058_/X VGND VGND VPWR VPWR _16228_/X sky130_fd_sc_hd__a22o_1
X_35062_ _35829_/CLK _35062_/D VGND VGND VPWR VPWR _35062_/Q sky130_fd_sc_hd__dfxtp_1
X_32274_ _36114_/CLK _32274_/D VGND VGND VPWR VPWR _32274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34013_ _36188_/CLK _34013_/D VGND VGND VPWR VPWR _34013_/Q sky130_fd_sc_hd__dfxtp_1
X_31225_ _27754_/X _35834_/Q _31231_/S VGND VGND VPWR VPWR _31226_/A sky130_fd_sc_hd__mux2_1
X_16159_ _16155_/X _16158_/X _16044_/X _16046_/X VGND VGND VPWR VPWR _16176_/B sky130_fd_sc_hd__o211a_1
XFILLER_114_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31156_ _27652_/X _35801_/Q _31168_/S VGND VGND VPWR VPWR _31157_/A sky130_fd_sc_hd__mux2_1
X_30107_ _30107_/A VGND VGND VPWR VPWR _35304_/D sky130_fd_sc_hd__clkbuf_1
X_19918_ _19811_/X _19916_/X _19917_/X _19816_/X VGND VGND VPWR VPWR _19918_/X sky130_fd_sc_hd__a22o_1
XFILLER_87_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31087_ _35769_/Q input29/X _31095_/S VGND VGND VPWR VPWR _31088_/A sky130_fd_sc_hd__mux2_1
X_35964_ _35964_/CLK _35964_/D VGND VGND VPWR VPWR _35964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19849_ _19845_/X _19848_/X _19818_/X VGND VGND VPWR VPWR _19850_/D sky130_fd_sc_hd__o21ba_1
X_30038_ _30065_/S VGND VGND VPWR VPWR _30057_/S sky130_fd_sc_hd__buf_4
XFILLER_111_973 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34915_ _34915_/CLK _34915_/D VGND VGND VPWR VPWR _34915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35895_ _35895_/CLK _35895_/D VGND VGND VPWR VPWR _35895_/Q sky130_fd_sc_hd__dfxtp_1
X_22860_ _32917_/Q _32853_/Q _32789_/Q _32725_/Q _20584_/X _20587_/X VGND VGND VPWR
+ VPWR _22860_/X sky130_fd_sc_hd__mux4_1
X_34846_ _36245_/CLK _34846_/D VGND VGND VPWR VPWR _34846_/Q sky130_fd_sc_hd__dfxtp_1
X_21811_ _21805_/X _21810_/X _21732_/X VGND VGND VPWR VPWR _21835_/A sky130_fd_sc_hd__o21ba_1
XFILLER_3_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34777_ _34911_/CLK _34777_/D VGND VGND VPWR VPWR _34777_/Q sky130_fd_sc_hd__dfxtp_1
X_22791_ _22505_/X _22789_/X _22790_/X _22510_/X VGND VGND VPWR VPWR _22791_/X sky130_fd_sc_hd__a22o_1
XFILLER_25_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31989_ _34914_/CLK _31989_/D VGND VGND VPWR VPWR _31989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_252_CLK clkbuf_6_63__f_CLK/X VGND VGND VPWR VPWR _34185_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_3_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24530_ _22891_/X _32791_/Q _24546_/S VGND VGND VPWR VPWR _24531_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33728_ _35646_/CLK _33728_/D VGND VGND VPWR VPWR _33728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21742_ _21736_/X _21739_/X _21740_/X _21741_/X VGND VGND VPWR VPWR _21767_/B sky130_fd_sc_hd__o211a_1
XPHY_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24461_ _24461_/A VGND VGND VPWR VPWR _32758_/D sky130_fd_sc_hd__clkbuf_1
X_33659_ _33661_/CLK _33659_/D VGND VGND VPWR VPWR _33659_/Q sky130_fd_sc_hd__dfxtp_1
X_21673_ _21666_/X _21672_/X _21387_/X _21388_/X VGND VGND VPWR VPWR _21690_/B sky130_fd_sc_hd__o211a_1
XFILLER_24_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26200_ _26200_/A VGND VGND VPWR VPWR _33549_/D sky130_fd_sc_hd__clkbuf_1
X_23412_ _32216_/Q _23411_/X _23418_/S VGND VGND VPWR VPWR _23413_/A sky130_fd_sc_hd__mux2_1
X_20624_ _22506_/A VGND VGND VPWR VPWR _20624_/X sky130_fd_sc_hd__clkbuf_8
X_27180_ input42/X VGND VGND VPWR VPWR _27180_/X sky130_fd_sc_hd__buf_4
X_24392_ _24524_/S VGND VGND VPWR VPWR _24411_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_162_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26131_ _26131_/A VGND VGND VPWR VPWR _33516_/D sky130_fd_sc_hd__clkbuf_1
X_35329_ _35841_/CLK _35329_/D VGND VGND VPWR VPWR _35329_/Q sky130_fd_sc_hd__dfxtp_1
X_23343_ _32188_/Q _23265_/X _23359_/S VGND VGND VPWR VPWR _23344_/A sky130_fd_sc_hd__mux2_1
X_20555_ _20551_/X _20554_/X _20138_/A VGND VGND VPWR VPWR _20577_/A sky130_fd_sc_hd__o21ba_1
XFILLER_20_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26062_ _24967_/X _33484_/Q _26072_/S VGND VGND VPWR VPWR _26063_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23274_ input6/X VGND VGND VPWR VPWR _23274_/X sky130_fd_sc_hd__buf_6
X_20486_ _20482_/X _20485_/X _20171_/A VGND VGND VPWR VPWR _20487_/D sky130_fd_sc_hd__o21ba_1
X_25013_ _24821_/X _32989_/Q _25017_/S VGND VGND VPWR VPWR _25014_/A sky130_fd_sc_hd__mux2_1
X_22225_ _33410_/Q _33346_/Q _33282_/Q _33218_/Q _22080_/X _22081_/X VGND VGND VPWR
+ VPWR _22225_/X sky130_fd_sc_hd__mux4_1
XFILLER_69_1152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29821_ _29821_/A VGND VGND VPWR VPWR _35168_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22156_ _34176_/Q _34112_/Q _34048_/Q _33984_/Q _22046_/X _22047_/X VGND VGND VPWR
+ VPWR _22156_/X sky130_fd_sc_hd__mux4_1
XFILLER_65_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_900 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21107_ _33122_/Q _36002_/Q _32994_/Q _32930_/Q _20956_/X _20957_/X VGND VGND VPWR
+ VPWR _21107_/X sky130_fd_sc_hd__mux4_1
X_29752_ _35136_/Q _29460_/X _29766_/S VGND VGND VPWR VPWR _29753_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_1472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22087_ _32638_/Q _32574_/Q _32510_/Q _35966_/Q _21876_/X _22013_/X VGND VGND VPWR
+ VPWR _22087_/X sky130_fd_sc_hd__mux4_1
X_26964_ _26964_/A VGND VGND VPWR VPWR _33908_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28703_ _34670_/Q _27109_/X _28713_/S VGND VGND VPWR VPWR _28704_/A sky130_fd_sc_hd__mux2_1
X_25915_ _25915_/A VGND VGND VPWR VPWR _33414_/D sky130_fd_sc_hd__clkbuf_1
X_21038_ _22598_/A VGND VGND VPWR VPWR _21038_/X sky130_fd_sc_hd__buf_6
X_29683_ _29683_/A VGND VGND VPWR VPWR _35103_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26895_ _26895_/A VGND VGND VPWR VPWR _33876_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_491_CLK clkbuf_6_9__f_CLK/X VGND VGND VPWR VPWR _35685_/CLK sky130_fd_sc_hd__clkbuf_16
X_28634_ _27816_/X _34638_/Q _28640_/S VGND VGND VPWR VPWR _28635_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25846_ _25846_/A VGND VGND VPWR VPWR _33381_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28565_ _27714_/X _34605_/Q _28577_/S VGND VGND VPWR VPWR _28566_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25777_ _24945_/X _33349_/Q _25781_/S VGND VGND VPWR VPWR _25778_/A sky130_fd_sc_hd__mux2_1
X_22989_ _22989_/A VGND VGND VPWR VPWR _32054_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_243_CLK clkbuf_6_61__f_CLK/X VGND VGND VPWR VPWR _36105_/CLK sky130_fd_sc_hd__clkbuf_16
X_27516_ _34139_/Q _27050_/X _27524_/S VGND VGND VPWR VPWR _27517_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24728_ _22984_/X _32885_/Q _24744_/S VGND VGND VPWR VPWR _24729_/A sky130_fd_sc_hd__mux2_1
X_28496_ _28496_/A VGND VGND VPWR VPWR _34572_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_242_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27447_ _27447_/A VGND VGND VPWR VPWR _34106_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_230_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24659_ _23082_/X _32853_/Q _24659_/S VGND VGND VPWR VPWR _24660_/A sky130_fd_sc_hd__mux2_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17200_ _17906_/A VGND VGND VPWR VPWR _17200_/X sky130_fd_sc_hd__buf_6
XFILLER_204_1112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18180_ _34706_/Q _34642_/Q _34578_/Q _34514_/Q _17998_/X _17999_/X VGND VGND VPWR
+ VPWR _18180_/X sky130_fd_sc_hd__mux4_1
X_27378_ _27378_/A VGND VGND VPWR VPWR _34073_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17131_ _16853_/X _17129_/X _17130_/X _16856_/X VGND VGND VPWR VPWR _17131_/X sky130_fd_sc_hd__a22o_1
X_29117_ _29117_/A VGND VGND VPWR VPWR _34865_/D sky130_fd_sc_hd__clkbuf_1
X_26329_ _26329_/A VGND VGND VPWR VPWR _33610_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29048_ _34833_/Q _27217_/X _29048_/S VGND VGND VPWR VPWR _29049_/A sky130_fd_sc_hd__mux2_1
X_17062_ _17986_/A VGND VGND VPWR VPWR _17062_/X sky130_fd_sc_hd__buf_4
XFILLER_144_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_870 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16013_ _16001_/X _16004_/X _16007_/X _16012_/X VGND VGND VPWR VPWR _16013_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31010_ _35733_/Q input60/X _31010_/S VGND VGND VPWR VPWR _31011_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17964_ _17709_/X _17962_/X _17963_/X _17712_/X VGND VGND VPWR VPWR _17964_/X sky130_fd_sc_hd__a22o_1
XFILLER_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19703_ _19703_/A _19703_/B _19703_/C _19703_/D VGND VGND VPWR VPWR _19704_/A sky130_fd_sc_hd__or4_2
XFILLER_111_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16915_ _16915_/A VGND VGND VPWR VPWR _31981_/D sky130_fd_sc_hd__clkbuf_1
X_32961_ _36033_/CLK _32961_/D VGND VGND VPWR VPWR _32961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17895_ _17891_/X _17894_/X _17857_/X VGND VGND VPWR VPWR _17903_/C sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_482_CLK _35560_/CLK VGND VGND VPWR VPWR _36075_/CLK sky130_fd_sc_hd__clkbuf_16
X_34700_ _35147_/CLK _34700_/D VGND VGND VPWR VPWR _34700_/Q sky130_fd_sc_hd__dfxtp_1
X_31912_ _31912_/A VGND VGND VPWR VPWR _36159_/D sky130_fd_sc_hd__clkbuf_1
X_19634_ _19634_/A VGND VGND VPWR VPWR _32441_/D sky130_fd_sc_hd__buf_2
X_16846_ _17905_/A VGND VGND VPWR VPWR _16846_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_38_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35680_ _35747_/CLK _35680_/D VGND VGND VPWR VPWR _35680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32892_ _35964_/CLK _32892_/D VGND VGND VPWR VPWR _32892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34631_ _34633_/CLK _34631_/D VGND VGND VPWR VPWR _34631_/Q sky130_fd_sc_hd__dfxtp_1
X_31843_ _23258_/X _36127_/Q _31843_/S VGND VGND VPWR VPWR _31844_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19565_ _19458_/X _19563_/X _19564_/X _19463_/X VGND VGND VPWR VPWR _19565_/X sky130_fd_sc_hd__a22o_1
XFILLER_59_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16777_ _33898_/Q _33834_/Q _33770_/Q _36074_/Q _16671_/X _16672_/X VGND VGND VPWR
+ VPWR _16777_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_234_CLK clkbuf_6_55__f_CLK/X VGND VGND VPWR VPWR _36113_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_207_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18516_ _18512_/X _18515_/X _18315_/X VGND VGND VPWR VPWR _18542_/A sky130_fd_sc_hd__o21ba_1
XFILLER_222_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34562_ _34691_/CLK _34562_/D VGND VGND VPWR VPWR _34562_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31774_ _36094_/Q input35/X _31792_/S VGND VGND VPWR VPWR _31775_/A sky130_fd_sc_hd__mux2_1
X_19496_ _19492_/X _19495_/X _19465_/X VGND VGND VPWR VPWR _19497_/D sky130_fd_sc_hd__o21ba_1
XFILLER_146_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33513_ _33897_/CLK _33513_/D VGND VGND VPWR VPWR _33513_/Q sky130_fd_sc_hd__dfxtp_1
X_30725_ _30725_/A VGND VGND VPWR VPWR _35597_/D sky130_fd_sc_hd__clkbuf_1
X_18447_ _20164_/A VGND VGND VPWR VPWR _18447_/X sky130_fd_sc_hd__buf_6
X_34493_ _35194_/CLK _34493_/D VGND VGND VPWR VPWR _34493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36232_ _36235_/CLK _36232_/D VGND VGND VPWR VPWR _36232_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33444_ _34151_/CLK _33444_/D VGND VGND VPWR VPWR _33444_/Q sky130_fd_sc_hd__dfxtp_1
X_18378_ _19453_/A VGND VGND VPWR VPWR _18378_/X sky130_fd_sc_hd__buf_4
X_30656_ _30656_/A VGND VGND VPWR VPWR _35564_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36163_ _36163_/CLK _36163_/D VGND VGND VPWR VPWR _36163_/Q sky130_fd_sc_hd__dfxtp_1
X_17329_ _34425_/Q _36153_/Q _34297_/Q _34233_/Q _17229_/X _17230_/X VGND VGND VPWR
+ VPWR _17329_/X sky130_fd_sc_hd__mux4_1
X_33375_ _35615_/CLK _33375_/D VGND VGND VPWR VPWR _33375_/Q sky130_fd_sc_hd__dfxtp_1
X_30587_ _35532_/Q _29497_/X _30597_/S VGND VGND VPWR VPWR _30588_/A sky130_fd_sc_hd__mux2_1
XFILLER_222_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35114_ _35564_/CLK _35114_/D VGND VGND VPWR VPWR _35114_/Q sky130_fd_sc_hd__dfxtp_1
X_20340_ _34190_/Q _34126_/Q _34062_/Q _33998_/Q _20099_/X _20100_/X VGND VGND VPWR
+ VPWR _20340_/X sky130_fd_sc_hd__mux4_1
X_32326_ _32905_/CLK _32326_/D VGND VGND VPWR VPWR _32326_/Q sky130_fd_sc_hd__dfxtp_1
X_36094_ _36095_/CLK _36094_/D VGND VGND VPWR VPWR _36094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_49__f_CLK clkbuf_5_24_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_49__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_35045_ _35168_/CLK _35045_/D VGND VGND VPWR VPWR _35045_/Q sky130_fd_sc_hd__dfxtp_1
X_20271_ _20164_/X _20269_/X _20270_/X _20169_/X VGND VGND VPWR VPWR _20271_/X sky130_fd_sc_hd__a22o_1
X_32257_ _34626_/CLK _32257_/D VGND VGND VPWR VPWR _32257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22010_ _21806_/X _22008_/X _22009_/X _21809_/X VGND VGND VPWR VPWR _22010_/X sky130_fd_sc_hd__a22o_1
X_31208_ _27729_/X _35826_/Q _31210_/S VGND VGND VPWR VPWR _31209_/A sky130_fd_sc_hd__mux2_1
XFILLER_216_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_1016 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32188_ _36135_/CLK _32188_/D VGND VGND VPWR VPWR _32188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31139_ _35794_/Q input57/X _31145_/S VGND VGND VPWR VPWR _31140_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23961_ _23058_/X _32525_/Q _23969_/S VGND VGND VPWR VPWR _23962_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35947_ _35947_/CLK _35947_/D VGND VGND VPWR VPWR _35947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_233_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_473_CLK clkbuf_6_10__f_CLK/X VGND VGND VPWR VPWR _35630_/CLK sky130_fd_sc_hd__clkbuf_16
X_25700_ _24830_/X _33312_/Q _25718_/S VGND VGND VPWR VPWR _25701_/A sky130_fd_sc_hd__mux2_1
X_22912_ input63/X VGND VGND VPWR VPWR _22912_/X sky130_fd_sc_hd__buf_2
XFILLER_96_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26680_ _33774_/Q _23305_/X _26690_/S VGND VGND VPWR VPWR _26681_/A sky130_fd_sc_hd__mux2_1
X_23892_ _22956_/X _32492_/Q _23906_/S VGND VGND VPWR VPWR _23893_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35878_ _35945_/CLK _35878_/D VGND VGND VPWR VPWR _35878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22843_ _34452_/Q _36180_/Q _34324_/Q _34260_/Q _20667_/X _20669_/X VGND VGND VPWR
+ VPWR _22843_/X sky130_fd_sc_hd__mux4_1
X_25631_ _25631_/A VGND VGND VPWR VPWR _33279_/D sky130_fd_sc_hd__clkbuf_1
X_34829_ _34956_/CLK _34829_/D VGND VGND VPWR VPWR _34829_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_225_CLK clkbuf_6_53__f_CLK/X VGND VGND VPWR VPWR _34441_/CLK sky130_fd_sc_hd__clkbuf_16
X_28350_ _28350_/A VGND VGND VPWR VPWR _34503_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22774_ _35666_/Q _35026_/Q _34386_/Q _33746_/Q _20712_/X _20713_/X VGND VGND VPWR
+ VPWR _22774_/X sky130_fd_sc_hd__mux4_1
X_25562_ _24827_/X _33247_/Q _25562_/S VGND VGND VPWR VPWR _25563_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27301_ _34037_/Q _27131_/X _27317_/S VGND VGND VPWR VPWR _27302_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24513_ _24513_/A VGND VGND VPWR VPWR _32783_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21725_ _34164_/Q _34100_/Q _34036_/Q _33972_/Q _21693_/X _21694_/X VGND VGND VPWR
+ VPWR _21725_/X sky130_fd_sc_hd__mux4_1
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25493_ _24923_/X _33214_/Q _25511_/S VGND VGND VPWR VPWR _25494_/A sky130_fd_sc_hd__mux2_1
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28281_ _28281_/A VGND VGND VPWR VPWR _34470_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_223_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27232_ _27232_/A _27232_/B _25132_/A VGND VGND VPWR VPWR _27233_/A sky130_fd_sc_hd__or3b_1
XFILLER_157_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_578 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21656_ _33906_/Q _33842_/Q _33778_/Q _36082_/Q _21624_/X _21625_/X VGND VGND VPWR
+ VPWR _21656_/X sky130_fd_sc_hd__mux4_1
XFILLER_40_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24444_ _24444_/A VGND VGND VPWR VPWR _32750_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_185_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20607_ _22515_/A VGND VGND VPWR VPWR _20607_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_137_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27163_ _33983_/Q _27162_/X _27187_/S VGND VGND VPWR VPWR _27164_/A sky130_fd_sc_hd__mux2_1
X_24375_ _23061_/X _32718_/Q _24381_/S VGND VGND VPWR VPWR _24376_/A sky130_fd_sc_hd__mux2_1
X_21587_ _21453_/X _21585_/X _21586_/X _21456_/X VGND VGND VPWR VPWR _21587_/X sky130_fd_sc_hd__a22o_1
XFILLER_32_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23326_ _23326_/A VGND VGND VPWR VPWR _32180_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26114_ _26114_/A VGND VGND VPWR VPWR _33508_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20538_ _18301_/X _20536_/X _20537_/X _18307_/X VGND VGND VPWR VPWR _20538_/X sky130_fd_sc_hd__a22o_1
XFILLER_197_1255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27094_ _33961_/Q _27093_/X _27094_/S VGND VGND VPWR VPWR _27095_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26045_ _24942_/X _33476_/Q _26051_/S VGND VGND VPWR VPWR _26046_/A sky130_fd_sc_hd__mux2_1
X_23257_ _23257_/A VGND VGND VPWR VPWR _32158_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20469_ _32146_/Q _32338_/Q _32402_/Q _35922_/Q _20286_/X _19311_/A VGND VGND VPWR
+ VPWR _20469_/X sky130_fd_sc_hd__mux4_1
XFILLER_84_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22208_ _22561_/A VGND VGND VPWR VPWR _22208_/X sky130_fd_sc_hd__buf_4
XFILLER_165_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23188_ _23030_/X _32132_/Q _23194_/S VGND VGND VPWR VPWR _23189_/A sky130_fd_sc_hd__mux2_1
XTAP_6611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29804_ _29804_/A VGND VGND VPWR VPWR _35160_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22139_ _35455_/Q _35391_/Q _35327_/Q _35263_/Q _21854_/X _21855_/X VGND VGND VPWR
+ VPWR _22139_/X sky130_fd_sc_hd__mux4_1
XTAP_6644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27996_ _27996_/A VGND VGND VPWR VPWR _34335_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29735_ _35128_/Q _29435_/X _29745_/S VGND VGND VPWR VPWR _29736_/A sky130_fd_sc_hd__mux2_1
XTAP_6688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26947_ _26947_/A VGND VGND VPWR VPWR _33900_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16700_ _34152_/Q _34088_/Q _34024_/Q _33960_/Q _16387_/X _16388_/X VGND VGND VPWR
+ VPWR _16700_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_464_CLK clkbuf_6_11__f_CLK/X VGND VGND VPWR VPWR _35692_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_248_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29666_ _35095_/Q _29333_/X _29682_/S VGND VGND VPWR VPWR _29667_/A sky130_fd_sc_hd__mux2_1
XTAP_5987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17680_ _35203_/Q _35139_/Q _35075_/Q _32259_/Q _17363_/X _17364_/X VGND VGND VPWR
+ VPWR _17680_/X sky130_fd_sc_hd__mux4_1
XFILLER_43_1188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26878_ _33868_/Q _23469_/X _26888_/S VGND VGND VPWR VPWR _26879_/A sky130_fd_sc_hd__mux2_1
XTAP_5998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28617_ _27791_/X _34630_/Q _28619_/S VGND VGND VPWR VPWR _28618_/A sky130_fd_sc_hd__mux2_1
X_16631_ _16493_/X _16629_/X _16630_/X _16498_/X VGND VGND VPWR VPWR _16631_/X sky130_fd_sc_hd__a22o_1
X_25829_ _25829_/A VGND VGND VPWR VPWR _33373_/D sky130_fd_sc_hd__clkbuf_1
X_29597_ _29597_/A VGND VGND VPWR VPWR _35062_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_216_CLK clkbuf_6_52__f_CLK/X VGND VGND VPWR VPWR _35147_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_204_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_732 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19350_ _19350_/A _19350_/B _19350_/C _19350_/D VGND VGND VPWR VPWR _19351_/A sky130_fd_sc_hd__or4_4
XFILLER_62_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16562_ _16562_/A VGND VGND VPWR VPWR _31971_/D sky130_fd_sc_hd__clkbuf_1
X_28548_ _27689_/X _34597_/Q _28556_/S VGND VGND VPWR VPWR _28549_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18301_ _20164_/A VGND VGND VPWR VPWR _18301_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_243_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19281_ _19281_/A VGND VGND VPWR VPWR _32431_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28479_ _28479_/A VGND VGND VPWR VPWR _34564_/D sky130_fd_sc_hd__clkbuf_1
X_16493_ _17905_/A VGND VGND VPWR VPWR _16493_/X sky130_fd_sc_hd__buf_4
XFILLER_231_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18232_ _18228_/X _18231_/X _17846_/A _17847_/A VGND VGND VPWR VPWR _18247_/B sky130_fd_sc_hd__o211a_1
X_30510_ _30510_/A VGND VGND VPWR VPWR _35495_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31490_ _31490_/A VGND VGND VPWR VPWR _35959_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18163_ _33938_/Q _33874_/Q _33810_/Q _36114_/Q _16062_/X _16064_/X VGND VGND VPWR
+ VPWR _18163_/X sky130_fd_sc_hd__mux4_1
X_30441_ _35463_/Q _29481_/X _30441_/S VGND VGND VPWR VPWR _30442_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_1352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17114_ _17110_/X _17113_/X _16798_/X VGND VGND VPWR VPWR _17122_/C sky130_fd_sc_hd__o21ba_1
XFILLER_184_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33160_ _33160_/CLK _33160_/D VGND VGND VPWR VPWR _33160_/Q sky130_fd_sc_hd__dfxtp_1
X_18094_ _34959_/Q _34895_/Q _34831_/Q _34767_/Q _17866_/X _17867_/X VGND VGND VPWR
+ VPWR _18094_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30372_ _35430_/Q _29379_/X _30378_/S VGND VGND VPWR VPWR _30373_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_1238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32111_ _35952_/CLK _32111_/D VGND VGND VPWR VPWR _32111_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17045_ _16800_/X _17043_/X _17044_/X _16803_/X VGND VGND VPWR VPWR _17045_/X sky130_fd_sc_hd__a22o_1
X_33091_ _35779_/CLK _33091_/D VGND VGND VPWR VPWR _33091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_873 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32042_ _35820_/CLK _32042_/D VGND VGND VPWR VPWR _32042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18996_ _18992_/X _18995_/X _18759_/X VGND VGND VPWR VPWR _18997_/D sky130_fd_sc_hd__o21ba_1
XFILLER_225_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35801_ _35801_/CLK _35801_/D VGND VGND VPWR VPWR _35801_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17947_ _33931_/Q _33867_/Q _33803_/Q _36107_/Q _17730_/X _17731_/X VGND VGND VPWR
+ VPWR _17947_/X sky130_fd_sc_hd__mux4_1
XFILLER_113_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33993_ _34121_/CLK _33993_/D VGND VGND VPWR VPWR _33993_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_455_CLK clkbuf_6_14__f_CLK/X VGND VGND VPWR VPWR _36141_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_239_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35732_ _35733_/CLK _35732_/D VGND VGND VPWR VPWR _35732_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32944_ _36144_/CLK _32944_/D VGND VGND VPWR VPWR _32944_/Q sky130_fd_sc_hd__dfxtp_1
X_17878_ _33417_/Q _33353_/Q _33289_/Q _33225_/Q _17833_/X _17834_/X VGND VGND VPWR
+ VPWR _17878_/X sky130_fd_sc_hd__mux4_1
XFILLER_241_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19617_ _20099_/A VGND VGND VPWR VPWR _19617_/X sky130_fd_sc_hd__buf_6
XFILLER_66_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16829_ _16825_/X _16828_/X _16787_/X _16788_/X VGND VGND VPWR VPWR _16844_/B sky130_fd_sc_hd__o211a_1
XFILLER_96_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35663_ _35663_/CLK _35663_/D VGND VGND VPWR VPWR _35663_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32875_ _32875_/CLK _32875_/D VGND VGND VPWR VPWR _32875_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_207_CLK clkbuf_6_54__f_CLK/X VGND VGND VPWR VPWR _35658_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_207_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31826_ _31826_/A VGND VGND VPWR VPWR _36118_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34614_ _36024_/CLK _34614_/D VGND VGND VPWR VPWR _34614_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19548_ _32887_/Q _32823_/Q _32759_/Q _32695_/Q _19293_/X _19294_/X VGND VGND VPWR
+ VPWR _19548_/X sky130_fd_sc_hd__mux4_1
X_35594_ _35723_/CLK _35594_/D VGND VGND VPWR VPWR _35594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34545_ _35056_/CLK _34545_/D VGND VGND VPWR VPWR _34545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31757_ _36086_/Q input26/X _31771_/S VGND VGND VPWR VPWR _31758_/A sky130_fd_sc_hd__mux2_1
X_19479_ _32117_/Q _32309_/Q _32373_/Q _35893_/Q _19227_/X _19368_/X VGND VGND VPWR
+ VPWR _19479_/X sky130_fd_sc_hd__mux4_1
XFILLER_55_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21510_ _34413_/Q _36141_/Q _34285_/Q _34221_/Q _21476_/X _21477_/X VGND VGND VPWR
+ VPWR _21510_/X sky130_fd_sc_hd__mux4_1
X_30708_ _30708_/A VGND VGND VPWR VPWR _35589_/D sky130_fd_sc_hd__clkbuf_1
X_22490_ _35657_/Q _35017_/Q _34377_/Q _33737_/Q _22450_/X _22451_/X VGND VGND VPWR
+ VPWR _22490_/X sky130_fd_sc_hd__mux4_1
XFILLER_167_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34476_ _35754_/CLK _34476_/D VGND VGND VPWR VPWR _34476_/Q sky130_fd_sc_hd__dfxtp_1
X_31688_ _31688_/A _31688_/B VGND VGND VPWR VPWR _31821_/S sky130_fd_sc_hd__nor2_8
X_33427_ _36179_/CLK _33427_/D VGND VGND VPWR VPWR _33427_/Q sky130_fd_sc_hd__dfxtp_1
X_36215_ _36219_/CLK _36215_/D VGND VGND VPWR VPWR _36215_/Q sky130_fd_sc_hd__dfxtp_1
X_21441_ _34923_/Q _34859_/Q _34795_/Q _34731_/Q _21407_/X _21408_/X VGND VGND VPWR
+ VPWR _21441_/X sky130_fd_sc_hd__mux4_1
XFILLER_222_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30639_ _30639_/A VGND VGND VPWR VPWR _35556_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36146_ _36146_/CLK _36146_/D VGND VGND VPWR VPWR _36146_/Q sky130_fd_sc_hd__dfxtp_1
X_24160_ _24160_/A VGND VGND VPWR VPWR _32617_/D sky130_fd_sc_hd__clkbuf_1
X_33358_ _33425_/CLK _33358_/D VGND VGND VPWR VPWR _33358_/Q sky130_fd_sc_hd__dfxtp_1
X_21372_ _34154_/Q _34090_/Q _34026_/Q _33962_/Q _21340_/X _21341_/X VGND VGND VPWR
+ VPWR _21372_/X sky130_fd_sc_hd__mux4_1
XFILLER_174_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23111_ _23111_/A VGND VGND VPWR VPWR _32095_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_1351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20323_ _35725_/Q _32236_/Q _35597_/Q _35533_/Q _18293_/X _18295_/X VGND VGND VPWR
+ VPWR _20323_/X sky130_fd_sc_hd__mux4_1
XFILLER_135_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32309_ _32885_/CLK _32309_/D VGND VGND VPWR VPWR _32309_/Q sky130_fd_sc_hd__dfxtp_1
X_24091_ _23049_/X _32586_/Q _24105_/S VGND VGND VPWR VPWR _24092_/A sky130_fd_sc_hd__mux2_1
X_36077_ _36077_/CLK _36077_/D VGND VGND VPWR VPWR _36077_/Q sky130_fd_sc_hd__dfxtp_1
X_33289_ _33420_/CLK _33289_/D VGND VGND VPWR VPWR _33289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35028_ _35668_/CLK _35028_/D VGND VGND VPWR VPWR _35028_/Q sky130_fd_sc_hd__dfxtp_1
X_23042_ input46/X VGND VGND VPWR VPWR _23042_/X sky130_fd_sc_hd__buf_2
XFILLER_118_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20254_ _32907_/Q _32843_/Q _32779_/Q _32715_/Q _19999_/X _20000_/X VGND VGND VPWR
+ VPWR _20254_/X sky130_fd_sc_hd__mux4_1
XFILLER_143_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27850_ _27655_/X _34266_/Q _27860_/S VGND VGND VPWR VPWR _27851_/A sky130_fd_sc_hd__mux2_1
XFILLER_135_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20185_ _32137_/Q _32329_/Q _32393_/Q _35913_/Q _19933_/X _20074_/X VGND VGND VPWR
+ VPWR _20185_/X sky130_fd_sc_hd__mux4_1
XFILLER_27_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26801_ _26801_/A VGND VGND VPWR VPWR _33831_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27781_ _27781_/A VGND VGND VPWR VPWR _34242_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24993_ _24993_/A VGND VGND VPWR VPWR _32980_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_229_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29520_ _29520_/A VGND VGND VPWR VPWR _35027_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_446_CLK clkbuf_leaf_61_CLK/A VGND VGND VPWR VPWR _35951_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_218_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26732_ _33799_/Q _23450_/X _26732_/S VGND VGND VPWR VPWR _26733_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23944_ _23033_/X _32517_/Q _23948_/S VGND VGND VPWR VPWR _23945_/A sky130_fd_sc_hd__mux2_1
XTAP_3804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29451_ _35005_/Q _29450_/X _29451_/S VGND VGND VPWR VPWR _29452_/A sky130_fd_sc_hd__mux2_1
XTAP_3848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26663_ _33766_/Q _23280_/X _26669_/S VGND VGND VPWR VPWR _26664_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_245_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23875_ _22931_/X _32484_/Q _23885_/S VGND VGND VPWR VPWR _23876_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28402_ _28513_/S VGND VGND VPWR VPWR _28421_/S sky130_fd_sc_hd__buf_6
X_25614_ _25614_/A VGND VGND VPWR VPWR _33271_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_226_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22826_ _32660_/Q _32596_/Q _32532_/Q _35988_/Q _22582_/X _21477_/A VGND VGND VPWR
+ VPWR _22826_/X sky130_fd_sc_hd__mux4_1
X_29382_ input9/X VGND VGND VPWR VPWR _29382_/X sky130_fd_sc_hd__buf_2
XFILLER_77_1240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26594_ _26594_/A VGND VGND VPWR VPWR _33735_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_832 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28333_ _27770_/X _34495_/Q _28349_/S VGND VGND VPWR VPWR _28334_/A sky130_fd_sc_hd__mux2_1
X_25545_ _25545_/A VGND VGND VPWR VPWR _33238_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22757_ _22757_/A _22757_/B _22757_/C _22757_/D VGND VGND VPWR VPWR _22758_/A sky130_fd_sc_hd__or4_4
XFILLER_12_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28264_ _28264_/A VGND VGND VPWR VPWR _34462_/D sky130_fd_sc_hd__clkbuf_1
X_21708_ _35699_/Q _32207_/Q _35571_/Q _35507_/Q _21564_/X _21565_/X VGND VGND VPWR
+ VPWR _21708_/X sky130_fd_sc_hd__mux4_1
XFILLER_201_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22688_ _20601_/X _22686_/X _22687_/X _20607_/X VGND VGND VPWR VPWR _22688_/X sky130_fd_sc_hd__a22o_1
XFILLER_13_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25476_ _24899_/X _33206_/Q _25490_/S VGND VGND VPWR VPWR _25477_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_1298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27215_ _34000_/Q _27214_/X _27218_/S VGND VGND VPWR VPWR _27216_/A sky130_fd_sc_hd__mux2_1
X_21639_ _35441_/Q _35377_/Q _35313_/Q _35249_/Q _21501_/X _21502_/X VGND VGND VPWR
+ VPWR _21639_/X sky130_fd_sc_hd__mux4_1
X_24427_ _24427_/A VGND VGND VPWR VPWR _32742_/D sky130_fd_sc_hd__clkbuf_1
X_28195_ _28243_/S VGND VGND VPWR VPWR _28214_/S sky130_fd_sc_hd__buf_4
XFILLER_166_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_1030 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27146_ input30/X VGND VGND VPWR VPWR _27146_/X sky130_fd_sc_hd__buf_2
X_24358_ _23036_/X _32710_/Q _24360_/S VGND VGND VPWR VPWR _24359_/A sky130_fd_sc_hd__mux2_1
XFILLER_176_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23309_ _23309_/A VGND VGND VPWR VPWR _30877_/A sky130_fd_sc_hd__buf_12
XFILLER_153_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24289_ _22934_/X _32677_/Q _24297_/S VGND VGND VPWR VPWR _24290_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27077_ _27077_/A VGND VGND VPWR VPWR _33955_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_862 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_6_32__f_CLK clkbuf_5_16_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_32__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_26028_ _24917_/X _33468_/Q _26030_/S VGND VGND VPWR VPWR _26029_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18850_ _35427_/Q _35363_/Q _35299_/Q _35235_/Q _18848_/X _18849_/X VGND VGND VPWR
+ VPWR _18850_/X sky130_fd_sc_hd__mux4_1
XTAP_6430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17801_ _34183_/Q _34119_/Q _34055_/Q _33991_/Q _17799_/X _17800_/X VGND VGND VPWR
+ VPWR _17801_/X sky130_fd_sc_hd__mux4_1
XTAP_6452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18781_ _33057_/Q _32033_/Q _35809_/Q _35745_/Q _18672_/X _18673_/X VGND VGND VPWR
+ VPWR _18781_/X sky130_fd_sc_hd__mux4_1
XTAP_6485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27979_ _34327_/Q _27038_/X _27995_/S VGND VGND VPWR VPWR _27980_/A sky130_fd_sc_hd__mux2_1
XTAP_5740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15993_ _17799_/A VGND VGND VPWR VPWR _15993_/X sky130_fd_sc_hd__buf_4
XTAP_5751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_437_CLK clkbuf_6_36__f_CLK/X VGND VGND VPWR VPWR _36144_/CLK sky130_fd_sc_hd__clkbuf_16
X_17732_ _33925_/Q _33861_/Q _33797_/Q _36101_/Q _17730_/X _17731_/X VGND VGND VPWR
+ VPWR _17732_/X sky130_fd_sc_hd__mux4_1
XTAP_5762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29718_ _35120_/Q _29410_/X _29724_/S VGND VGND VPWR VPWR _29719_/A sky130_fd_sc_hd__mux2_1
XTAP_5773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30990_ _35723_/Q input49/X _31002_/S VGND VGND VPWR VPWR _30991_/A sky130_fd_sc_hd__mux2_1
XTAP_5795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_1299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29649_ _29649_/A VGND VGND VPWR VPWR _35087_/D sky130_fd_sc_hd__clkbuf_1
X_17663_ _32643_/Q _32579_/Q _32515_/Q _35971_/Q _17629_/X _17413_/X VGND VGND VPWR
+ VPWR _17663_/X sky130_fd_sc_hd__mux4_1
XFILLER_63_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_996 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_635 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19402_ _33139_/Q _36019_/Q _33011_/Q _32947_/Q _19362_/X _19363_/X VGND VGND VPWR
+ VPWR _19402_/X sky130_fd_sc_hd__mux4_1
X_16614_ _35621_/Q _34981_/Q _34341_/Q _33701_/Q _16438_/X _16439_/X VGND VGND VPWR
+ VPWR _16614_/X sky130_fd_sc_hd__mux4_1
X_32660_ _35988_/CLK _32660_/D VGND VGND VPWR VPWR _32660_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17594_ _33921_/Q _33857_/Q _33793_/Q _36097_/Q _17377_/X _17378_/X VGND VGND VPWR
+ VPWR _17594_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31611_ _27726_/X _36017_/Q _31615_/S VGND VGND VPWR VPWR _31612_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19333_ _32881_/Q _32817_/Q _32753_/Q _32689_/Q _19293_/X _19294_/X VGND VGND VPWR
+ VPWR _19333_/X sky130_fd_sc_hd__mux4_1
XFILLER_245_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16545_ _35683_/Q _32190_/Q _35555_/Q _35491_/Q _16258_/X _16259_/X VGND VGND VPWR
+ VPWR _16545_/X sky130_fd_sc_hd__mux4_1
X_32591_ _35983_/CLK _32591_/D VGND VGND VPWR VPWR _32591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34330_ _35610_/CLK _34330_/D VGND VGND VPWR VPWR _34330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31542_ _31542_/A VGND VGND VPWR VPWR _35984_/D sky130_fd_sc_hd__clkbuf_1
X_19264_ _20099_/A VGND VGND VPWR VPWR _19264_/X sky130_fd_sc_hd__buf_4
XFILLER_149_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16476_ _16472_/X _16475_/X _16434_/X _16435_/X VGND VGND VPWR VPWR _16491_/B sky130_fd_sc_hd__o211a_1
X_18215_ _16060_/X _18213_/X _18214_/X _16072_/X VGND VGND VPWR VPWR _18215_/X sky130_fd_sc_hd__a22o_1
XFILLER_31_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34261_ _36181_/CLK _34261_/D VGND VGND VPWR VPWR _34261_/Q sky130_fd_sc_hd__dfxtp_1
X_31473_ _31473_/A VGND VGND VPWR VPWR _35951_/D sky130_fd_sc_hd__clkbuf_1
X_19195_ _32877_/Q _32813_/Q _32749_/Q _32685_/Q _18940_/X _18941_/X VGND VGND VPWR
+ VPWR _19195_/X sky130_fd_sc_hd__mux4_1
X_36000_ _36003_/CLK _36000_/D VGND VGND VPWR VPWR _36000_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_762 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33212_ _33913_/CLK _33212_/D VGND VGND VPWR VPWR _33212_/Q sky130_fd_sc_hd__dfxtp_1
X_18146_ _35473_/Q _35409_/Q _35345_/Q _35281_/Q _17960_/X _17961_/X VGND VGND VPWR
+ VPWR _18146_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30424_ _30424_/A VGND VGND VPWR VPWR _35454_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34192_ _34192_/CLK _34192_/D VGND VGND VPWR VPWR _34192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33143_ _36024_/CLK _33143_/D VGND VGND VPWR VPWR _33143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18077_ _33167_/Q _36047_/Q _33039_/Q _32975_/Q _17768_/X _17769_/X VGND VGND VPWR
+ VPWR _18077_/X sky130_fd_sc_hd__mux4_1
X_30355_ _35422_/Q _29354_/X _30357_/S VGND VGND VPWR VPWR _30356_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1079 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17028_ _17022_/X _17027_/X _16779_/X VGND VGND VPWR VPWR _17050_/A sky130_fd_sc_hd__o21ba_1
XFILLER_176_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33074_ _35187_/CLK _33074_/D VGND VGND VPWR VPWR _33074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30286_ _30286_/A VGND VGND VPWR VPWR _35389_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32025_ _34135_/CLK _32025_/D VGND VGND VPWR VPWR _32025_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18979_ _32103_/Q _32295_/Q _32359_/Q _35879_/Q _18874_/X _18662_/X VGND VGND VPWR
+ VPWR _18979_/X sky130_fd_sc_hd__mux4_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_428_CLK clkbuf_6_38__f_CLK/X VGND VGND VPWR VPWR _36149_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21990_ _35643_/Q _35003_/Q _34363_/Q _33723_/Q _21744_/X _21745_/X VGND VGND VPWR
+ VPWR _21990_/X sky130_fd_sc_hd__mux4_1
X_33976_ _35320_/CLK _33976_/D VGND VGND VPWR VPWR _33976_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20941_ _34909_/Q _34845_/Q _34781_/Q _34717_/Q _20696_/X _20698_/X VGND VGND VPWR
+ VPWR _20941_/X sky130_fd_sc_hd__mux4_1
X_35715_ _35715_/CLK _35715_/D VGND VGND VPWR VPWR _35715_/Q sky130_fd_sc_hd__dfxtp_1
X_32927_ _35807_/CLK _32927_/D VGND VGND VPWR VPWR _32927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20872_ _20691_/X _20870_/X _20871_/X _20701_/X VGND VGND VPWR VPWR _20872_/X sky130_fd_sc_hd__a22o_1
X_35646_ _35646_/CLK _35646_/D VGND VGND VPWR VPWR _35646_/Q sky130_fd_sc_hd__dfxtp_1
X_23660_ _23660_/A VGND VGND VPWR VPWR _32320_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32858_ _34070_/CLK _32858_/D VGND VGND VPWR VPWR _32858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22611_ _22505_/X _22609_/X _22610_/X _22510_/X VGND VGND VPWR VPWR _22611_/X sky130_fd_sc_hd__a22o_1
XFILLER_35_882 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31809_ _36111_/Q input53/X _31813_/S VGND VGND VPWR VPWR _31810_/A sky130_fd_sc_hd__mux2_1
X_23591_ _23702_/S VGND VGND VPWR VPWR _23610_/S sky130_fd_sc_hd__buf_4
XFILLER_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32789_ _32802_/CLK _32789_/D VGND VGND VPWR VPWR _32789_/Q sky130_fd_sc_hd__dfxtp_1
X_35577_ _35577_/CLK _35577_/D VGND VGND VPWR VPWR _35577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22542_ _22542_/A VGND VGND VPWR VPWR _36234_/D sky130_fd_sc_hd__clkbuf_1
X_25330_ _33138_/Q _23381_/X _25332_/S VGND VGND VPWR VPWR _25331_/A sky130_fd_sc_hd__mux2_1
X_34528_ _34594_/CLK _34528_/D VGND VGND VPWR VPWR _34528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22473_ _22473_/A _22473_/B _22473_/C _22473_/D VGND VGND VPWR VPWR _22474_/A sky130_fd_sc_hd__or4_4
X_25261_ _33106_/Q _23487_/X _25267_/S VGND VGND VPWR VPWR _25262_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34459_ _36127_/CLK _34459_/D VGND VGND VPWR VPWR _34459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27000_ _33926_/Q _23447_/X _27002_/S VGND VGND VPWR VPWR _27001_/A sky130_fd_sc_hd__mux2_1
X_24212_ _32642_/Q _23435_/X _24222_/S VGND VGND VPWR VPWR _24213_/A sky130_fd_sc_hd__mux2_1
X_21424_ _33131_/Q _36011_/Q _33003_/Q _32939_/Q _21309_/X _21310_/X VGND VGND VPWR
+ VPWR _21424_/X sky130_fd_sc_hd__mux4_1
XFILLER_147_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25192_ _33073_/Q _23364_/X _25196_/S VGND VGND VPWR VPWR _25193_/A sky130_fd_sc_hd__mux2_1
X_24143_ _32609_/Q _23265_/X _24159_/S VGND VGND VPWR VPWR _24144_/A sky130_fd_sc_hd__mux2_1
X_36129_ _36129_/CLK _36129_/D VGND VGND VPWR VPWR _36129_/Q sky130_fd_sc_hd__dfxtp_1
X_21355_ _35689_/Q _32196_/Q _35561_/Q _35497_/Q _21211_/X _21212_/X VGND VGND VPWR
+ VPWR _21355_/X sky130_fd_sc_hd__mux4_1
XFILLER_135_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20306_ _20302_/X _20305_/X _20171_/X VGND VGND VPWR VPWR _20307_/D sky130_fd_sc_hd__o21ba_1
X_24074_ _23024_/X _32578_/Q _24084_/S VGND VGND VPWR VPWR _24075_/A sky130_fd_sc_hd__mux2_1
X_28951_ _28951_/A VGND VGND VPWR VPWR _34786_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21286_ _35431_/Q _35367_/Q _35303_/Q _35239_/Q _21148_/X _21149_/X VGND VGND VPWR
+ VPWR _21286_/X sky130_fd_sc_hd__mux4_1
XFILLER_122_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23025_ _23024_/X _32066_/Q _23040_/S VGND VGND VPWR VPWR _23026_/A sky130_fd_sc_hd__mux2_1
X_27902_ _27732_/X _34291_/Q _27902_/S VGND VGND VPWR VPWR _27903_/A sky130_fd_sc_hd__mux2_1
X_20237_ _34442_/Q _36170_/Q _34314_/Q _34250_/Q _20235_/X _20236_/X VGND VGND VPWR
+ VPWR _20237_/X sky130_fd_sc_hd__mux4_1
XFILLER_104_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28882_ _34754_/Q _27171_/X _28892_/S VGND VGND VPWR VPWR _28883_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27833_ _27833_/A VGND VGND VPWR VPWR _34259_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20168_ _34952_/Q _34888_/Q _34824_/Q _34760_/Q _20166_/X _20167_/X VGND VGND VPWR
+ VPWR _20168_/X sky130_fd_sc_hd__mux4_1
XFILLER_77_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_419_CLK clkbuf_6_33__f_CLK/X VGND VGND VPWR VPWR _35439_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_44_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27764_ _27763_/X _34237_/Q _27764_/S VGND VGND VPWR VPWR _27765_/A sky130_fd_sc_hd__mux2_1
X_20099_ _20099_/A VGND VGND VPWR VPWR _20099_/X sky130_fd_sc_hd__clkbuf_8
X_24976_ input53/X VGND VGND VPWR VPWR _24976_/X sky130_fd_sc_hd__buf_6
XTAP_3601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29503_ input52/X VGND VGND VPWR VPWR _29503_/X sky130_fd_sc_hd__buf_2
XTAP_4357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26715_ _26715_/A VGND VGND VPWR VPWR _33790_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23927_ _23008_/X _32509_/Q _23927_/S VGND VGND VPWR VPWR _23928_/A sky130_fd_sc_hd__mux2_1
XTAP_3645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27695_ input9/X VGND VGND VPWR VPWR _27695_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29434_ _29434_/A VGND VGND VPWR VPWR _34999_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_229_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26646_ _33758_/Q _23255_/X _26648_/S VGND VGND VPWR VPWR _26647_/A sky130_fd_sc_hd__mux2_1
XTAP_3678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23858_ _22906_/X _32476_/Q _23864_/S VGND VGND VPWR VPWR _23859_/A sky130_fd_sc_hd__mux2_1
XTAP_3689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22809_ _22805_/X _22808_/X _22457_/A VGND VGND VPWR VPWR _22817_/C sky130_fd_sc_hd__o21ba_1
X_29365_ _34977_/Q _29364_/X _29389_/S VGND VGND VPWR VPWR _29366_/A sky130_fd_sc_hd__mux2_1
X_26577_ _24927_/X _33727_/Q _26593_/S VGND VGND VPWR VPWR _26578_/A sky130_fd_sc_hd__mux2_1
XTAP_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23789_ _23789_/A VGND VGND VPWR VPWR _32380_/D sky130_fd_sc_hd__clkbuf_1
X_16330_ _35677_/Q _32183_/Q _35549_/Q _35485_/Q _16258_/X _16259_/X VGND VGND VPWR
+ VPWR _16330_/X sky130_fd_sc_hd__mux4_1
XFILLER_125_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28316_ _27745_/X _34487_/Q _28328_/S VGND VGND VPWR VPWR _28317_/A sky130_fd_sc_hd__mux2_1
X_25528_ _24976_/X _33231_/Q _25532_/S VGND VGND VPWR VPWR _25529_/A sky130_fd_sc_hd__mux2_1
X_29296_ _29296_/A VGND VGND VPWR VPWR _34950_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28247_ _27639_/X _34454_/Q _28265_/S VGND VGND VPWR VPWR _28248_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16261_ _35611_/Q _34971_/Q _34331_/Q _33691_/Q _16053_/X _16055_/X VGND VGND VPWR
+ VPWR _16261_/X sky130_fd_sc_hd__mux4_1
X_25459_ _24874_/X _33198_/Q _25469_/S VGND VGND VPWR VPWR _25460_/A sky130_fd_sc_hd__mux2_1
X_18000_ _34700_/Q _34636_/Q _34572_/Q _34508_/Q _17998_/X _17999_/X VGND VGND VPWR
+ VPWR _18000_/X sky130_fd_sc_hd__mux4_1
XFILLER_127_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16192_ _35673_/Q _32179_/Q _35545_/Q _35481_/Q _16049_/X _16050_/X VGND VGND VPWR
+ VPWR _16192_/X sky130_fd_sc_hd__mux4_1
X_28178_ _28178_/A VGND VGND VPWR VPWR _34421_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27129_ _33972_/Q _27127_/X _27156_/S VGND VGND VPWR VPWR _27130_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30140_ _35320_/Q _29435_/X _30150_/S VGND VGND VPWR VPWR _30141_/A sky130_fd_sc_hd__mux2_1
X_19951_ _34946_/Q _34882_/Q _34818_/Q _34754_/Q _19813_/X _19814_/X VGND VGND VPWR
+ VPWR _19951_/X sky130_fd_sc_hd__mux4_1
XFILLER_218_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18902_ _18800_/X _18900_/X _18901_/X _18803_/X VGND VGND VPWR VPWR _18902_/X sky130_fd_sc_hd__a22o_1
X_30071_ _35287_/Q _29333_/X _30087_/S VGND VGND VPWR VPWR _30072_/A sky130_fd_sc_hd__mux2_1
X_19882_ _20235_/A VGND VGND VPWR VPWR _19882_/X sky130_fd_sc_hd__buf_6
XFILLER_49_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_727 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18833_ _18793_/X _18831_/X _18832_/X _18798_/X VGND VGND VPWR VPWR _18833_/X sky130_fd_sc_hd__a22o_1
XTAP_6260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33830_ _36066_/CLK _33830_/D VGND VGND VPWR VPWR _33830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18764_ _34145_/Q _34081_/Q _34017_/Q _33953_/Q _18687_/X _18688_/X VGND VGND VPWR
+ VPWR _18764_/X sky130_fd_sc_hd__mux4_1
XTAP_5570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17715_ _34692_/Q _34628_/Q _34564_/Q _34500_/Q _17645_/X _17646_/X VGND VGND VPWR
+ VPWR _17715_/X sky130_fd_sc_hd__mux4_1
XTAP_5592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33761_ _36065_/CLK _33761_/D VGND VGND VPWR VPWR _33761_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30973_ _35715_/Q input40/X _30981_/S VGND VGND VPWR VPWR _30974_/A sky130_fd_sc_hd__mux2_1
X_18695_ _32607_/Q _32543_/Q _32479_/Q _35935_/Q _18517_/X _18654_/X VGND VGND VPWR
+ VPWR _18695_/X sky130_fd_sc_hd__mux4_1
XTAP_4880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35500_ _35564_/CLK _35500_/D VGND VGND VPWR VPWR _35500_/Q sky130_fd_sc_hd__dfxtp_1
X_17646_ _17999_/A VGND VGND VPWR VPWR _17646_/X sky130_fd_sc_hd__clkbuf_4
X_32712_ _32906_/CLK _32712_/D VGND VGND VPWR VPWR _32712_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_1359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33692_ _36060_/CLK _33692_/D VGND VGND VPWR VPWR _33692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32643_ _35779_/CLK _32643_/D VGND VGND VPWR VPWR _32643_/Q sky130_fd_sc_hd__dfxtp_1
X_35431_ _35433_/CLK _35431_/D VGND VGND VPWR VPWR _35431_/Q sky130_fd_sc_hd__dfxtp_1
X_17577_ _17356_/X _17575_/X _17576_/X _17359_/X VGND VGND VPWR VPWR _17577_/X sky130_fd_sc_hd__a22o_1
XFILLER_56_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19316_ _19105_/X _19314_/X _19315_/X _19110_/X VGND VGND VPWR VPWR _19316_/X sky130_fd_sc_hd__a22o_1
X_16528_ _16522_/X _16527_/X _16459_/X VGND VGND VPWR VPWR _16529_/D sky130_fd_sc_hd__o21ba_1
X_35362_ _35553_/CLK _35362_/D VGND VGND VPWR VPWR _35362_/Q sky130_fd_sc_hd__dfxtp_1
X_32574_ _36031_/CLK _32574_/D VGND VGND VPWR VPWR _32574_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34313_ _36171_/CLK _34313_/D VGND VGND VPWR VPWR _34313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31525_ _27797_/X _35976_/Q _31543_/S VGND VGND VPWR VPWR _31526_/A sky130_fd_sc_hd__mux2_1
X_19247_ _19243_/X _19246_/X _19112_/X VGND VGND VPWR VPWR _19248_/D sky130_fd_sc_hd__o21ba_1
XFILLER_91_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35293_ _35677_/CLK _35293_/D VGND VGND VPWR VPWR _35293_/Q sky130_fd_sc_hd__dfxtp_1
X_16459_ _17871_/A VGND VGND VPWR VPWR _16459_/X sky130_fd_sc_hd__buf_2
XFILLER_34_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_1181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34244_ _36164_/CLK _34244_/D VGND VGND VPWR VPWR _34244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19178_ _34412_/Q _36140_/Q _34284_/Q _34220_/Q _19176_/X _19177_/X VGND VGND VPWR
+ VPWR _19178_/X sky130_fd_sc_hd__mux4_1
X_31456_ _31456_/A VGND VGND VPWR VPWR _35943_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18129_ _33681_/Q _33617_/Q _33553_/Q _33489_/Q _17906_/X _17907_/X VGND VGND VPWR
+ VPWR _18129_/X sky130_fd_sc_hd__mux4_1
X_30407_ _30407_/A VGND VGND VPWR VPWR _35446_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_754 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34175_ _35456_/CLK _34175_/D VGND VGND VPWR VPWR _34175_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31387_ _27794_/X _35911_/Q _31387_/S VGND VGND VPWR VPWR _31388_/A sky130_fd_sc_hd__mux2_1
X_33126_ _36007_/CLK _33126_/D VGND VGND VPWR VPWR _33126_/Q sky130_fd_sc_hd__dfxtp_1
X_21140_ _20953_/X _21138_/X _21139_/X _20959_/X VGND VGND VPWR VPWR _21140_/X sky130_fd_sc_hd__a22o_1
X_30338_ _30470_/S VGND VGND VPWR VPWR _30357_/S sky130_fd_sc_hd__buf_6
XFILLER_172_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21071_ _33121_/Q _36001_/Q _32993_/Q _32929_/Q _20956_/X _20957_/X VGND VGND VPWR
+ VPWR _21071_/X sky130_fd_sc_hd__mux4_1
X_33057_ _35812_/CLK _33057_/D VGND VGND VPWR VPWR _33057_/Q sky130_fd_sc_hd__dfxtp_1
X_30269_ _35381_/Q _29426_/X _30285_/S VGND VGND VPWR VPWR _30270_/A sky130_fd_sc_hd__mux2_1
X_20022_ _19811_/X _20020_/X _20021_/X _19816_/X VGND VGND VPWR VPWR _20022_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_1204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32008_ _36209_/CLK _32008_/D VGND VGND VPWR VPWR _32008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24830_ input2/X VGND VGND VPWR VPWR _24830_/X sky130_fd_sc_hd__buf_4
XFILLER_41_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24761_ _23033_/X _32901_/Q _24765_/S VGND VGND VPWR VPWR _24762_/A sky130_fd_sc_hd__mux2_1
X_21973_ _33659_/Q _33595_/Q _33531_/Q _33467_/Q _21800_/X _21801_/X VGND VGND VPWR
+ VPWR _21973_/X sky130_fd_sc_hd__mux4_1
X_33959_ _34149_/CLK _33959_/D VGND VGND VPWR VPWR _33959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26500_ _26500_/A VGND VGND VPWR VPWR _33690_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23712_ _23712_/A VGND VGND VPWR VPWR _32343_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27480_ _34122_/Q _27196_/X _27494_/S VGND VGND VPWR VPWR _27481_/A sky130_fd_sc_hd__mux2_1
XFILLER_187_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20924_ _33117_/Q _35997_/Q _32989_/Q _32925_/Q _20624_/X _20625_/X VGND VGND VPWR
+ VPWR _20924_/X sky130_fd_sc_hd__mux4_1
XFILLER_55_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_242_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24692_ _22931_/X _32868_/Q _24702_/S VGND VGND VPWR VPWR _24693_/A sky130_fd_sc_hd__mux2_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26431_ _26431_/A VGND VGND VPWR VPWR _33658_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20855_ _32859_/Q _32795_/Q _32731_/Q _32667_/Q _20637_/X _20639_/X VGND VGND VPWR
+ VPWR _20855_/X sky130_fd_sc_hd__mux4_1
X_35629_ _35630_/CLK _35629_/D VGND VGND VPWR VPWR _35629_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23643_ _23643_/A VGND VGND VPWR VPWR _32312_/D sky130_fd_sc_hd__clkbuf_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29150_ _34881_/Q _27168_/X _29162_/S VGND VGND VPWR VPWR _29151_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26362_ _26362_/A VGND VGND VPWR VPWR _33625_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23574_ _23574_/A VGND VGND VPWR VPWR _32279_/D sky130_fd_sc_hd__clkbuf_1
X_20786_ _33113_/Q _35993_/Q _32985_/Q _32921_/Q _20624_/X _20625_/X VGND VGND VPWR
+ VPWR _20786_/X sky130_fd_sc_hd__mux4_1
X_28101_ _28101_/A VGND VGND VPWR VPWR _34385_/D sky130_fd_sc_hd__clkbuf_1
X_25313_ _25403_/S VGND VGND VPWR VPWR _25332_/S sky130_fd_sc_hd__buf_4
X_22525_ _35722_/Q _32233_/Q _35594_/Q _35530_/Q _22270_/X _22271_/X VGND VGND VPWR
+ VPWR _22525_/X sky130_fd_sc_hd__mux4_1
XFILLER_161_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29081_ _34848_/Q _27065_/X _29099_/S VGND VGND VPWR VPWR _29082_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26293_ _26293_/A VGND VGND VPWR VPWR _33593_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28032_ _28032_/A VGND VGND VPWR VPWR _34352_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25244_ _25244_/A VGND VGND VPWR VPWR _33097_/D sky130_fd_sc_hd__clkbuf_1
X_22456_ _22309_/X _22454_/X _22455_/X _22312_/X VGND VGND VPWR VPWR _22456_/X sky130_fd_sc_hd__a22o_1
XFILLER_157_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21407_ _22466_/A VGND VGND VPWR VPWR _21407_/X sky130_fd_sc_hd__buf_4
X_22387_ _22309_/X _22383_/X _22386_/X _22312_/X VGND VGND VPWR VPWR _22387_/X sky130_fd_sc_hd__a22o_1
X_25175_ _33065_/Q _23289_/X _25175_/S VGND VGND VPWR VPWR _25176_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24126_ _32601_/Q _23240_/X _24138_/S VGND VGND VPWR VPWR _24127_/A sky130_fd_sc_hd__mux2_1
X_21338_ _21338_/A VGND VGND VPWR VPWR _36200_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29983_ _29983_/A VGND VGND VPWR VPWR _35245_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28934_ _28934_/A VGND VGND VPWR VPWR _34778_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21269_ _21093_/X _21267_/X _21268_/X _21098_/X VGND VGND VPWR VPWR _21269_/X sky130_fd_sc_hd__a22o_1
X_24057_ _22999_/X _32570_/Q _24063_/S VGND VGND VPWR VPWR _24058_/A sky130_fd_sc_hd__mux2_1
XFILLER_235_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23008_ input33/X VGND VGND VPWR VPWR _23008_/X sky130_fd_sc_hd__buf_2
XFILLER_104_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28865_ _34746_/Q _27146_/X _28871_/S VGND VGND VPWR VPWR _28866_/A sky130_fd_sc_hd__mux2_1
XFILLER_238_817 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27816_ input52/X VGND VGND VPWR VPWR _27816_/X sky130_fd_sc_hd__clkbuf_4
XTAP_4110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28796_ _34713_/Q _27044_/X _28808_/S VGND VGND VPWR VPWR _28797_/A sky130_fd_sc_hd__mux2_1
XTAP_4121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27747_ _27747_/A VGND VGND VPWR VPWR _34231_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24959_ _24958_/X _32969_/Q _24983_/S VGND VGND VPWR VPWR _24960_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17500_ _17351_/X _17496_/X _17499_/X _17354_/X VGND VGND VPWR VPWR _17500_/X sky130_fd_sc_hd__a22o_1
XTAP_4187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18480_ _18440_/X _18478_/X _18479_/X _18445_/X VGND VGND VPWR VPWR _18480_/X sky130_fd_sc_hd__a22o_1
XTAP_3464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27678_ _27677_/X _34209_/Q _27702_/S VGND VGND VPWR VPWR _27679_/A sky130_fd_sc_hd__mux2_1
XTAP_3475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17431_ _17935_/A VGND VGND VPWR VPWR _17431_/X sky130_fd_sc_hd__buf_6
XTAP_3497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29417_ _34994_/Q _29416_/X _29420_/S VGND VGND VPWR VPWR _29418_/A sky130_fd_sc_hd__mux2_1
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26629_ _26761_/S VGND VGND VPWR VPWR _26648_/S sky130_fd_sc_hd__buf_6
XFILLER_17_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29348_ input61/X VGND VGND VPWR VPWR _29348_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_144_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17362_ _34682_/Q _34618_/Q _34554_/Q _34490_/Q _17292_/X _17293_/X VGND VGND VPWR
+ VPWR _17362_/X sky130_fd_sc_hd__mux4_1
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19101_ _34666_/Q _34602_/Q _34538_/Q _34474_/Q _18886_/X _18887_/X VGND VGND VPWR
+ VPWR _19101_/X sky130_fd_sc_hd__mux4_1
XFILLER_198_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16313_ _16313_/A VGND VGND VPWR VPWR _31964_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29279_ _34942_/Q _27158_/X _29297_/S VGND VGND VPWR VPWR _29280_/A sky130_fd_sc_hd__mux2_1
XFILLER_203_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17293_ _17999_/A VGND VGND VPWR VPWR _17293_/X sky130_fd_sc_hd__buf_6
XFILLER_207_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31310_ _27680_/X _35874_/Q _31324_/S VGND VGND VPWR VPWR _31311_/A sky130_fd_sc_hd__mux2_1
X_19032_ _18747_/X _19030_/X _19031_/X _18750_/X VGND VGND VPWR VPWR _19032_/X sky130_fd_sc_hd__a22o_1
X_16244_ _33627_/Q _33563_/Q _33499_/Q _33435_/Q _16141_/X _16142_/X VGND VGND VPWR
+ VPWR _16244_/X sky130_fd_sc_hd__mux4_1
X_32290_ _32871_/CLK _32290_/D VGND VGND VPWR VPWR _32290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31241_ _31241_/A VGND VGND VPWR VPWR _35841_/D sky130_fd_sc_hd__clkbuf_1
X_16175_ _16169_/X _16174_/X _16104_/X VGND VGND VPWR VPWR _16176_/D sky130_fd_sc_hd__o21ba_1
XFILLER_154_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_916 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput107 _31983_/Q VGND VGND VPWR VPWR D1[25] sky130_fd_sc_hd__buf_2
XFILLER_217_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput118 _31993_/Q VGND VGND VPWR VPWR D1[35] sky130_fd_sc_hd__buf_2
XFILLER_114_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput129 _32003_/Q VGND VGND VPWR VPWR D1[45] sky130_fd_sc_hd__buf_2
X_31172_ _31172_/A VGND VGND VPWR VPWR _35808_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30123_ _35312_/Q _29410_/X _30129_/S VGND VGND VPWR VPWR _30124_/A sky130_fd_sc_hd__mux2_1
X_19934_ _32130_/Q _32322_/Q _32386_/Q _35906_/Q _19933_/X _19721_/X VGND VGND VPWR
+ VPWR _19934_/X sky130_fd_sc_hd__mux4_1
XFILLER_190_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35980_ _35980_/CLK _35980_/D VGND VGND VPWR VPWR _35980_/Q sky130_fd_sc_hd__dfxtp_1
X_30054_ _30054_/A VGND VGND VPWR VPWR _35279_/D sky130_fd_sc_hd__clkbuf_1
X_34931_ _35056_/CLK _34931_/D VGND VGND VPWR VPWR _34931_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19865_ _32640_/Q _32576_/Q _32512_/Q _35968_/Q _19576_/X _19713_/X VGND VGND VPWR
+ VPWR _19865_/X sky130_fd_sc_hd__mux4_1
XFILLER_96_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18816_ _35426_/Q _35362_/Q _35298_/Q _35234_/Q _18495_/X _18496_/X VGND VGND VPWR
+ VPWR _18816_/X sky130_fd_sc_hd__mux4_1
XFILLER_228_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34862_ _34926_/CLK _34862_/D VGND VGND VPWR VPWR _34862_/Q sky130_fd_sc_hd__dfxtp_1
X_19796_ _35710_/Q _32219_/Q _35582_/Q _35518_/Q _19617_/X _19618_/X VGND VGND VPWR
+ VPWR _19796_/X sky130_fd_sc_hd__mux4_1
XFILLER_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_888 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33813_ _36119_/CLK _33813_/D VGND VGND VPWR VPWR _33813_/Q sky130_fd_sc_hd__dfxtp_1
X_18747_ _19453_/A VGND VGND VPWR VPWR _18747_/X sky130_fd_sc_hd__buf_4
X_34793_ _34921_/CLK _34793_/D VGND VGND VPWR VPWR _34793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18678_ _35166_/Q _35102_/Q _35038_/Q _32158_/Q _18604_/X _18605_/X VGND VGND VPWR
+ VPWR _18678_/X sky130_fd_sc_hd__mux4_1
X_33744_ _35728_/CLK _33744_/D VGND VGND VPWR VPWR _33744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30956_ _35707_/Q input31/X _30960_/S VGND VGND VPWR VPWR _30957_/A sky130_fd_sc_hd__mux2_1
XFILLER_224_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17629_ _17982_/A VGND VGND VPWR VPWR _17629_/X sky130_fd_sc_hd__buf_6
X_33675_ _33869_/CLK _33675_/D VGND VGND VPWR VPWR _33675_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30887_ _35674_/Q input45/X _30897_/S VGND VGND VPWR VPWR _30888_/A sky130_fd_sc_hd__mux2_1
XFILLER_225_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35414_ _36119_/CLK _35414_/D VGND VGND VPWR VPWR _35414_/Q sky130_fd_sc_hd__dfxtp_1
X_20640_ _32854_/Q _32790_/Q _32726_/Q _32662_/Q _20637_/X _20639_/X VGND VGND VPWR
+ VPWR _20640_/X sky130_fd_sc_hd__mux4_1
X_32626_ _35955_/CLK _32626_/D VGND VGND VPWR VPWR _32626_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20571_ _35221_/Q _35157_/Q _35093_/Q _32277_/Q _18392_/X _18394_/X VGND VGND VPWR
+ VPWR _20571_/X sky130_fd_sc_hd__mux4_1
X_35345_ _35729_/CLK _35345_/D VGND VGND VPWR VPWR _35345_/Q sky130_fd_sc_hd__dfxtp_1
X_32557_ _35951_/CLK _32557_/D VGND VGND VPWR VPWR _32557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22310_ _35460_/Q _35396_/Q _35332_/Q _35268_/Q _22207_/X _22208_/X VGND VGND VPWR
+ VPWR _22310_/X sky130_fd_sc_hd__mux4_1
X_31508_ _27773_/X _35968_/Q _31522_/S VGND VGND VPWR VPWR _31509_/A sky130_fd_sc_hd__mux2_1
X_23290_ _32169_/Q _23289_/X _23290_/S VGND VGND VPWR VPWR _23291_/A sky130_fd_sc_hd__mux2_1
X_35276_ _35727_/CLK _35276_/D VGND VGND VPWR VPWR _35276_/Q sky130_fd_sc_hd__dfxtp_1
X_32488_ _35944_/CLK _32488_/D VGND VGND VPWR VPWR _32488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22241_ _35458_/Q _35394_/Q _35330_/Q _35266_/Q _22207_/X _22208_/X VGND VGND VPWR
+ VPWR _22241_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_1135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31439_ _31439_/A VGND VGND VPWR VPWR _35935_/D sky130_fd_sc_hd__clkbuf_1
X_34227_ _36017_/CLK _34227_/D VGND VGND VPWR VPWR _34227_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22172_ _35712_/Q _32222_/Q _35584_/Q _35520_/Q _21917_/X _21918_/X VGND VGND VPWR
+ VPWR _22172_/X sky130_fd_sc_hd__mux4_1
XFILLER_127_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34158_ _35630_/CLK _34158_/D VGND VGND VPWR VPWR _34158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21123_ _22316_/A VGND VGND VPWR VPWR _21123_/X sky130_fd_sc_hd__buf_6
X_33109_ _36052_/CLK _33109_/D VGND VGND VPWR VPWR _33109_/Q sky130_fd_sc_hd__dfxtp_1
X_34089_ _34153_/CLK _34089_/D VGND VGND VPWR VPWR _34089_/Q sky130_fd_sc_hd__dfxtp_1
X_26980_ _26980_/A VGND VGND VPWR VPWR _33916_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25931_ _24973_/X _33422_/Q _25937_/S VGND VGND VPWR VPWR _25932_/A sky130_fd_sc_hd__mux2_1
X_21054_ _22466_/A VGND VGND VPWR VPWR _21054_/X sky130_fd_sc_hd__buf_4
XFILLER_236_1394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20005_ _35716_/Q _32226_/Q _35588_/Q _35524_/Q _19970_/X _19971_/X VGND VGND VPWR
+ VPWR _20005_/X sky130_fd_sc_hd__mux4_1
XFILLER_28_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28650_ _30877_/B _31823_/B VGND VGND VPWR VPWR _28651_/A sky130_fd_sc_hd__and2b_1
XFILLER_86_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25862_ _24871_/X _33389_/Q _25874_/S VGND VGND VPWR VPWR _25863_/A sky130_fd_sc_hd__mux2_1
XFILLER_246_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27601_ _27601_/A VGND VGND VPWR VPWR _34179_/D sky130_fd_sc_hd__clkbuf_1
X_24813_ _24812_/X _32922_/Q _24828_/S VGND VGND VPWR VPWR _24814_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28581_ _28581_/A VGND VGND VPWR VPWR _34612_/D sky130_fd_sc_hd__clkbuf_1
X_25793_ _25793_/A VGND VGND VPWR VPWR _33356_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_966 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27532_ _27532_/A VGND VGND VPWR VPWR _34146_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24744_ _23008_/X _32893_/Q _24744_/S VGND VGND VPWR VPWR _24745_/A sky130_fd_sc_hd__mux2_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21956_ _22464_/A VGND VGND VPWR VPWR _21956_/X sky130_fd_sc_hd__buf_4
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27463_ _34114_/Q _27171_/X _27473_/S VGND VGND VPWR VPWR _27464_/A sky130_fd_sc_hd__mux2_1
X_20907_ _20678_/X _20903_/X _20906_/X _20688_/X VGND VGND VPWR VPWR _20907_/X sky130_fd_sc_hd__a22o_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24675_ _22906_/X _32860_/Q _24681_/S VGND VGND VPWR VPWR _24676_/A sky130_fd_sc_hd__mux2_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21887_ _21598_/X _21885_/X _21886_/X _21601_/X VGND VGND VPWR VPWR _21887_/X sky130_fd_sc_hd__a22o_1
X_29202_ _29202_/A VGND VGND VPWR VPWR _34905_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_215_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26414_ _26414_/A VGND VGND VPWR VPWR _33650_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23626_ _23626_/A VGND VGND VPWR VPWR _32304_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_1332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20838_ _34394_/Q _36122_/Q _34266_/Q _34202_/Q _20770_/X _20771_/X VGND VGND VPWR
+ VPWR _20838_/X sky130_fd_sc_hd__mux4_1
X_27394_ _34081_/Q _27069_/X _27410_/S VGND VGND VPWR VPWR _27395_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_243_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29133_ _34873_/Q _27143_/X _29141_/S VGND VGND VPWR VPWR _29134_/A sky130_fd_sc_hd__mux2_1
X_26345_ _26345_/A VGND VGND VPWR VPWR _33618_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23557_ _32273_/Q _23484_/X _23557_/S VGND VGND VPWR VPWR _23558_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20769_ _20678_/X _20767_/X _20768_/X _20688_/X VGND VGND VPWR VPWR _20769_/X sky130_fd_sc_hd__a22o_1
XFILLER_204_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29064_ _34840_/Q _27041_/X _29078_/S VGND VGND VPWR VPWR _29065_/A sky130_fd_sc_hd__mux2_1
X_22508_ _33674_/Q _33610_/Q _33546_/Q _33482_/Q _22506_/X _22507_/X VGND VGND VPWR
+ VPWR _22508_/X sky130_fd_sc_hd__mux4_1
XFILLER_195_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26276_ _26276_/A VGND VGND VPWR VPWR _33585_/D sky130_fd_sc_hd__clkbuf_1
X_23488_ _32241_/Q _23487_/X _23499_/S VGND VGND VPWR VPWR _23489_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28015_ _28015_/A VGND VGND VPWR VPWR _34344_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25227_ _25227_/A VGND VGND VPWR VPWR _33089_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22439_ _22432_/X _22437_/X _22438_/X VGND VGND VPWR VPWR _22473_/A sky130_fd_sc_hd__o21ba_1
XFILLER_182_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25158_ _25158_/A VGND VGND VPWR VPWR _33056_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_1478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24109_ _23076_/X _32595_/Q _24113_/S VGND VGND VPWR VPWR _24110_/A sky130_fd_sc_hd__mux2_1
X_17980_ _17912_/X _17978_/X _17979_/X _17915_/X VGND VGND VPWR VPWR _17980_/X sky130_fd_sc_hd__a22o_1
XFILLER_123_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25089_ _24933_/X _33025_/Q _25101_/S VGND VGND VPWR VPWR _25090_/A sky130_fd_sc_hd__mux2_1
X_29966_ _29966_/A VGND VGND VPWR VPWR _35237_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_215_1423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16931_ _16926_/X _16930_/X _16787_/X _16788_/X VGND VGND VPWR VPWR _16948_/B sky130_fd_sc_hd__o211a_1
X_28917_ _34771_/Q _27223_/X _28921_/S VGND VGND VPWR VPWR _28918_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29897_ _35205_/Q _29475_/X _29901_/S VGND VGND VPWR VPWR _29898_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_1478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19650_ _19644_/X _19649_/X _19440_/X _19441_/X VGND VGND VPWR VPWR _19671_/B sky130_fd_sc_hd__o211a_1
X_16862_ _32108_/Q _32300_/Q _32364_/Q _35884_/Q _16574_/X _16715_/X VGND VGND VPWR
+ VPWR _16862_/X sky130_fd_sc_hd__mux4_1
X_28848_ _34738_/Q _27121_/X _28850_/S VGND VGND VPWR VPWR _28849_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18601_ _18597_/X _18598_/X _18599_/X _18600_/X VGND VGND VPWR VPWR _18601_/X sky130_fd_sc_hd__a22o_1
X_19581_ _32120_/Q _32312_/Q _32376_/Q _35896_/Q _19580_/X _19368_/X VGND VGND VPWR
+ VPWR _19581_/X sky130_fd_sc_hd__mux4_1
X_28779_ _28779_/A VGND VGND VPWR VPWR _34706_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16793_ _35626_/Q _34986_/Q _34346_/Q _33706_/Q _16791_/X _16792_/X VGND VGND VPWR
+ VPWR _16793_/X sky130_fd_sc_hd__mux4_1
XFILLER_18_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18532_ _18528_/X _18531_/X _18375_/X VGND VGND VPWR VPWR _18542_/C sky130_fd_sc_hd__o21ba_1
X_30810_ _30810_/A VGND VGND VPWR VPWR _35637_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31790_ _36102_/Q input43/X _31792_/S VGND VGND VPWR VPWR _31791_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18463_ _35416_/Q _35352_/Q _35288_/Q _35224_/Q _18362_/X _18364_/X VGND VGND VPWR
+ VPWR _18463_/X sky130_fd_sc_hd__mux4_1
X_30741_ _30741_/A VGND VGND VPWR VPWR _35605_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_5_4_0_CLK clkbuf_5_7_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_4_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XTAP_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17414_ _32636_/Q _32572_/Q _32508_/Q _35964_/Q _17276_/X _17413_/X VGND VGND VPWR
+ VPWR _17414_/X sky130_fd_sc_hd__mux4_1
X_33460_ _36085_/CLK _33460_/D VGND VGND VPWR VPWR _33460_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18394_ _19177_/A VGND VGND VPWR VPWR _18394_/X sky130_fd_sc_hd__buf_4
X_30672_ _35572_/Q _29422_/X _30690_/S VGND VGND VPWR VPWR _30673_/A sky130_fd_sc_hd__mux2_1
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32411_ _34151_/CLK _32411_/D VGND VGND VPWR VPWR _32411_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17345_ _32122_/Q _32314_/Q _32378_/Q _35898_/Q _17280_/X _17068_/X VGND VGND VPWR
+ VPWR _17345_/X sky130_fd_sc_hd__mux4_1
X_33391_ _36080_/CLK _33391_/D VGND VGND VPWR VPWR _33391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32342_ _32856_/CLK _32342_/D VGND VGND VPWR VPWR _32342_/Q sky130_fd_sc_hd__dfxtp_1
X_35130_ _35577_/CLK _35130_/D VGND VGND VPWR VPWR _35130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17276_ _17982_/A VGND VGND VPWR VPWR _17276_/X sky130_fd_sc_hd__buf_6
XFILLER_174_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19015_ _20074_/A VGND VGND VPWR VPWR _19015_/X sky130_fd_sc_hd__clkbuf_4
X_16227_ _35610_/Q _34970_/Q _34330_/Q _33690_/Q _16053_/X _16055_/X VGND VGND VPWR
+ VPWR _16227_/X sky130_fd_sc_hd__mux4_1
XFILLER_173_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35061_ _36149_/CLK _35061_/D VGND VGND VPWR VPWR _35061_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32273_ _36115_/CLK _32273_/D VGND VGND VPWR VPWR _32273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34012_ _36211_/CLK _34012_/D VGND VGND VPWR VPWR _34012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31224_ _31224_/A VGND VGND VPWR VPWR _35833_/D sky130_fd_sc_hd__clkbuf_1
X_16158_ _16030_/X _16156_/X _16157_/X _16041_/X VGND VGND VPWR VPWR _16158_/X sky130_fd_sc_hd__a22o_1
XFILLER_177_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31155_ _31155_/A VGND VGND VPWR VPWR _35800_/D sky130_fd_sc_hd__clkbuf_1
X_16089_ _16078_/X _16081_/X _16086_/X _16088_/X VGND VGND VPWR VPWR _16089_/X sky130_fd_sc_hd__a22o_1
XFILLER_9_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30106_ _35304_/Q _29385_/X _30108_/S VGND VGND VPWR VPWR _30107_/A sky130_fd_sc_hd__mux2_1
X_19917_ _34945_/Q _34881_/Q _34817_/Q _34753_/Q _19813_/X _19814_/X VGND VGND VPWR
+ VPWR _19917_/X sky130_fd_sc_hd__mux4_1
X_31086_ _31086_/A VGND VGND VPWR VPWR _35768_/D sky130_fd_sc_hd__clkbuf_1
X_35963_ _36027_/CLK _35963_/D VGND VGND VPWR VPWR _35963_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_218_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30037_ _30037_/A VGND VGND VPWR VPWR _35271_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34914_ _34914_/CLK _34914_/D VGND VGND VPWR VPWR _34914_/Q sky130_fd_sc_hd__dfxtp_1
X_19848_ _19811_/X _19846_/X _19847_/X _19816_/X VGND VGND VPWR VPWR _19848_/X sky130_fd_sc_hd__a22o_1
XFILLER_69_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35894_ _35895_/CLK _35894_/D VGND VGND VPWR VPWR _35894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34845_ _36242_/CLK _34845_/D VGND VGND VPWR VPWR _34845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19779_ _19499_/X _19777_/X _19778_/X _19504_/X VGND VGND VPWR VPWR _19779_/X sky130_fd_sc_hd__a22o_1
XFILLER_84_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21810_ _21806_/X _21807_/X _21808_/X _21809_/X VGND VGND VPWR VPWR _21810_/X sky130_fd_sc_hd__a22o_1
X_34776_ _34907_/CLK _34776_/D VGND VGND VPWR VPWR _34776_/Q sky130_fd_sc_hd__dfxtp_1
X_22790_ _34195_/Q _34131_/Q _34067_/Q _34003_/Q _20649_/X _20650_/X VGND VGND VPWR
+ VPWR _22790_/X sky130_fd_sc_hd__mux4_1
XFILLER_58_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31988_ _34914_/CLK _31988_/D VGND VGND VPWR VPWR _31988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33727_ _36096_/CLK _33727_/D VGND VGND VPWR VPWR _33727_/Q sky130_fd_sc_hd__dfxtp_1
X_21741_ _22447_/A VGND VGND VPWR VPWR _21741_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_224_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30939_ _35699_/Q input22/X _30939_/S VGND VGND VPWR VPWR _30940_/A sky130_fd_sc_hd__mux2_1
XFILLER_212_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24460_ _22987_/X _32758_/Q _24474_/S VGND VGND VPWR VPWR _24461_/A sky130_fd_sc_hd__mux2_1
X_33658_ _34172_/CLK _33658_/D VGND VGND VPWR VPWR _33658_/Q sky130_fd_sc_hd__dfxtp_1
X_21672_ _21667_/X _21669_/X _21670_/X _21671_/X VGND VGND VPWR VPWR _21672_/X sky130_fd_sc_hd__a22o_1
X_23411_ input31/X VGND VGND VPWR VPWR _23411_/X sky130_fd_sc_hd__buf_4
X_20623_ _32598_/Q _32534_/Q _32470_/Q _35926_/Q _22466_/A _22317_/A VGND VGND VPWR
+ VPWR _20623_/X sky130_fd_sc_hd__mux4_1
X_32609_ _36002_/CLK _32609_/D VGND VGND VPWR VPWR _32609_/Q sky130_fd_sc_hd__dfxtp_1
X_24391_ _27840_/A _31553_/B VGND VGND VPWR VPWR _24524_/S sky130_fd_sc_hd__nand2_8
X_33589_ _34100_/CLK _33589_/D VGND VGND VPWR VPWR _33589_/Q sky130_fd_sc_hd__dfxtp_1
X_26130_ _24868_/X _33516_/Q _26144_/S VGND VGND VPWR VPWR _26131_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20554_ _18330_/X _20552_/X _20553_/X _18341_/X VGND VGND VPWR VPWR _20554_/X sky130_fd_sc_hd__a22o_1
X_35328_ _35839_/CLK _35328_/D VGND VGND VPWR VPWR _35328_/Q sky130_fd_sc_hd__dfxtp_1
X_23342_ _23342_/A VGND VGND VPWR VPWR _32187_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26061_ _26061_/A VGND VGND VPWR VPWR _33483_/D sky130_fd_sc_hd__clkbuf_1
X_20485_ _18360_/X _20483_/X _20484_/X _18372_/X VGND VGND VPWR VPWR _20485_/X sky130_fd_sc_hd__a22o_1
XFILLER_180_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23273_ _23273_/A VGND VGND VPWR VPWR _32163_/D sky130_fd_sc_hd__clkbuf_1
X_35259_ _35451_/CLK _35259_/D VGND VGND VPWR VPWR _35259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25012_ _25012_/A VGND VGND VPWR VPWR _32988_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22224_ _22152_/X _22222_/X _22223_/X _22157_/X VGND VGND VPWR VPWR _22224_/X sky130_fd_sc_hd__a22o_1
XFILLER_69_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22155_ _33664_/Q _33600_/Q _33536_/Q _33472_/Q _22153_/X _22154_/X VGND VGND VPWR
+ VPWR _22155_/X sky130_fd_sc_hd__mux4_1
X_29820_ _35168_/Q _29360_/X _29838_/S VGND VGND VPWR VPWR _29821_/A sky130_fd_sc_hd__mux2_1
XTAP_6804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21106_ _32610_/Q _32546_/Q _32482_/Q _35938_/Q _20817_/X _20954_/X VGND VGND VPWR
+ VPWR _21106_/X sky130_fd_sc_hd__mux4_1
XFILLER_47_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29751_ _29751_/A VGND VGND VPWR VPWR _35135_/D sky130_fd_sc_hd__clkbuf_1
X_22086_ _22079_/X _22084_/X _22085_/X VGND VGND VPWR VPWR _22120_/A sky130_fd_sc_hd__o21ba_1
X_26963_ _33908_/Q _23387_/X _26981_/S VGND VGND VPWR VPWR _26964_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_912 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25914_ _24948_/X _33414_/Q _25916_/S VGND VGND VPWR VPWR _25915_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28702_ _28702_/A VGND VGND VPWR VPWR _34669_/D sky130_fd_sc_hd__clkbuf_1
X_21037_ _35680_/Q _32186_/Q _35552_/Q _35488_/Q _20858_/X _20859_/X VGND VGND VPWR
+ VPWR _21037_/X sky130_fd_sc_hd__mux4_1
XFILLER_87_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29682_ _35103_/Q _29357_/X _29682_/S VGND VGND VPWR VPWR _29683_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26894_ _33876_/Q _23495_/X _26896_/S VGND VGND VPWR VPWR _26895_/A sky130_fd_sc_hd__mux2_1
XFILLER_219_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_248_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28633_ _28633_/A VGND VGND VPWR VPWR _34637_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_247_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25845_ _24846_/X _33381_/Q _25853_/S VGND VGND VPWR VPWR _25846_/A sky130_fd_sc_hd__mux2_1
XFILLER_235_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28564_ _28564_/A VGND VGND VPWR VPWR _34604_/D sky130_fd_sc_hd__clkbuf_1
X_25776_ _25776_/A VGND VGND VPWR VPWR _33348_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22988_ _22987_/X _32054_/Q _23009_/S VGND VGND VPWR VPWR _22989_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27515_ _27515_/A VGND VGND VPWR VPWR _34138_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24727_ _24727_/A VGND VGND VPWR VPWR _32884_/D sky130_fd_sc_hd__clkbuf_1
X_28495_ _27810_/X _34572_/Q _28505_/S VGND VGND VPWR VPWR _28496_/A sky130_fd_sc_hd__mux2_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21939_ _33914_/Q _33850_/Q _33786_/Q _36090_/Q _21624_/X _21625_/X VGND VGND VPWR
+ VPWR _21939_/X sky130_fd_sc_hd__mux4_1
XFILLER_76_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27446_ _34106_/Q _27146_/X _27452_/S VGND VGND VPWR VPWR _27447_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24658_ _24658_/A VGND VGND VPWR VPWR _32852_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_203_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_939 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23609_ _23609_/A VGND VGND VPWR VPWR _32296_/D sky130_fd_sc_hd__clkbuf_1
X_27377_ _34073_/Q _27044_/X _27389_/S VGND VGND VPWR VPWR _27378_/A sky130_fd_sc_hd__mux2_1
XFILLER_208_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24589_ _24589_/A VGND VGND VPWR VPWR _32819_/D sky130_fd_sc_hd__clkbuf_1
X_17130_ _33908_/Q _33844_/Q _33780_/Q _36084_/Q _17024_/X _17025_/X VGND VGND VPWR
+ VPWR _17130_/X sky130_fd_sc_hd__mux4_1
X_29116_ _34865_/Q _27118_/X _29120_/S VGND VGND VPWR VPWR _29117_/A sky130_fd_sc_hd__mux2_1
X_26328_ _24961_/X _33610_/Q _26342_/S VGND VGND VPWR VPWR _26329_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29047_ _29047_/A VGND VGND VPWR VPWR _34832_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_221_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17061_ _32626_/Q _32562_/Q _32498_/Q _35954_/Q _16923_/X _17060_/X VGND VGND VPWR
+ VPWR _17061_/X sky130_fd_sc_hd__mux4_1
X_26259_ _26259_/A VGND VGND VPWR VPWR _33577_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16012_ _33878_/Q _33814_/Q _33750_/Q _36054_/Q _16009_/X _16011_/X VGND VGND VPWR
+ VPWR _16012_/X sky130_fd_sc_hd__mux4_1
XFILLER_137_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_1253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17963_ _33099_/Q _32075_/Q _35851_/Q _35787_/Q _17784_/X _17785_/X VGND VGND VPWR
+ VPWR _17963_/X sky130_fd_sc_hd__mux4_1
X_29949_ _29949_/A VGND VGND VPWR VPWR _35229_/D sky130_fd_sc_hd__clkbuf_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19702_ _19698_/X _19701_/X _19465_/X VGND VGND VPWR VPWR _19703_/D sky130_fd_sc_hd__o21ba_1
XFILLER_239_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16914_ _16914_/A _16914_/B _16914_/C _16914_/D VGND VGND VPWR VPWR _16915_/A sky130_fd_sc_hd__or4_4
X_32960_ _35646_/CLK _32960_/D VGND VGND VPWR VPWR _32960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_215_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17894_ _17709_/X _17892_/X _17893_/X _17712_/X VGND VGND VPWR VPWR _17894_/X sky130_fd_sc_hd__a22o_1
XFILLER_38_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31911_ _23426_/X _36159_/Q _31927_/S VGND VGND VPWR VPWR _31912_/A sky130_fd_sc_hd__mux2_1
X_19633_ _19633_/A _19633_/B _19633_/C _19633_/D VGND VGND VPWR VPWR _19634_/A sky130_fd_sc_hd__or4_2
X_16845_ _16845_/A VGND VGND VPWR VPWR _31979_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32891_ _32891_/CLK _32891_/D VGND VGND VPWR VPWR _32891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34630_ _34694_/CLK _34630_/D VGND VGND VPWR VPWR _34630_/Q sky130_fd_sc_hd__dfxtp_1
X_31842_ _31842_/A VGND VGND VPWR VPWR _36126_/D sky130_fd_sc_hd__clkbuf_1
X_16776_ _33386_/Q _33322_/Q _33258_/Q _33194_/Q _16774_/X _16775_/X VGND VGND VPWR
+ VPWR _16776_/X sky130_fd_sc_hd__mux4_1
X_19564_ _34935_/Q _34871_/Q _34807_/Q _34743_/Q _19460_/X _19461_/X VGND VGND VPWR
+ VPWR _19564_/X sky130_fd_sc_hd__mux4_1
XFILLER_19_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18515_ _18447_/X _18513_/X _18514_/X _18450_/X VGND VGND VPWR VPWR _18515_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_722 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34561_ _34690_/CLK _34561_/D VGND VGND VPWR VPWR _34561_/Q sky130_fd_sc_hd__dfxtp_1
X_31773_ _31821_/S VGND VGND VPWR VPWR _31792_/S sky130_fd_sc_hd__clkbuf_8
XTAP_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19495_ _19458_/X _19493_/X _19494_/X _19463_/X VGND VGND VPWR VPWR _19495_/X sky130_fd_sc_hd__a22o_1
XTAP_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33512_ _35622_/CLK _33512_/D VGND VGND VPWR VPWR _33512_/Q sky130_fd_sc_hd__dfxtp_1
X_30724_ _35597_/Q _29500_/X _30732_/S VGND VGND VPWR VPWR _30725_/A sky130_fd_sc_hd__mux2_1
X_18446_ _18440_/X _18443_/X _18444_/X _18445_/X VGND VGND VPWR VPWR _18446_/X sky130_fd_sc_hd__a22o_1
X_34492_ _35197_/CLK _34492_/D VGND VGND VPWR VPWR _34492_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_36231_ _36235_/CLK _36231_/D VGND VGND VPWR VPWR _36231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18377_ _20065_/A VGND VGND VPWR VPWR _19453_/A sky130_fd_sc_hd__clkbuf_16
X_33443_ _34151_/CLK _33443_/D VGND VGND VPWR VPWR _33443_/Q sky130_fd_sc_hd__dfxtp_1
X_30655_ _35564_/Q _29398_/X _30669_/S VGND VGND VPWR VPWR _30656_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17328_ _17153_/X _17326_/X _17327_/X _17156_/X VGND VGND VPWR VPWR _17328_/X sky130_fd_sc_hd__a22o_1
XFILLER_239_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36162_ _36163_/CLK _36162_/D VGND VGND VPWR VPWR _36162_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33374_ _36205_/CLK _33374_/D VGND VGND VPWR VPWR _33374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30586_ _30586_/A VGND VGND VPWR VPWR _35531_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_1096 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35113_ _35177_/CLK _35113_/D VGND VGND VPWR VPWR _35113_/Q sky130_fd_sc_hd__dfxtp_1
X_32325_ _32901_/CLK _32325_/D VGND VGND VPWR VPWR _32325_/Q sky130_fd_sc_hd__dfxtp_1
X_17259_ _17253_/X _17258_/X _17151_/X VGND VGND VPWR VPWR _17267_/C sky130_fd_sc_hd__o21ba_1
X_36093_ _36093_/CLK _36093_/D VGND VGND VPWR VPWR _36093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20270_ _34955_/Q _34891_/Q _34827_/Q _34763_/Q _20166_/X _20167_/X VGND VGND VPWR
+ VPWR _20270_/X sky130_fd_sc_hd__mux4_1
X_32256_ _35715_/CLK _32256_/D VGND VGND VPWR VPWR _32256_/Q sky130_fd_sc_hd__dfxtp_1
X_35044_ _35490_/CLK _35044_/D VGND VGND VPWR VPWR _35044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31207_ _31207_/A VGND VGND VPWR VPWR _35825_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_170_CLK clkbuf_6_28__f_CLK/X VGND VGND VPWR VPWR _35221_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_157_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32187_ _35056_/CLK _32187_/D VGND VGND VPWR VPWR _32187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31138_ _31138_/A VGND VGND VPWR VPWR _35793_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23960_ _23960_/A VGND VGND VPWR VPWR _32524_/D sky130_fd_sc_hd__clkbuf_1
X_31069_ _31069_/A VGND VGND VPWR VPWR _35760_/D sky130_fd_sc_hd__clkbuf_1
X_35946_ _35946_/CLK _35946_/D VGND VGND VPWR VPWR _35946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22911_ _22911_/A VGND VGND VPWR VPWR _32029_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_229_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23891_ _23891_/A VGND VGND VPWR VPWR _32491_/D sky130_fd_sc_hd__clkbuf_1
X_35877_ _35945_/CLK _35877_/D VGND VGND VPWR VPWR _35877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_216_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25630_ _24927_/X _33279_/Q _25646_/S VGND VGND VPWR VPWR _25631_/A sky130_fd_sc_hd__mux2_1
X_34828_ _34956_/CLK _34828_/D VGND VGND VPWR VPWR _34828_/Q sky130_fd_sc_hd__dfxtp_1
X_22842_ _20648_/X _22840_/X _22841_/X _20658_/X VGND VGND VPWR VPWR _22842_/X sky130_fd_sc_hd__a22o_1
XFILLER_204_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25561_ _25561_/A VGND VGND VPWR VPWR _33246_/D sky130_fd_sc_hd__clkbuf_1
X_34759_ _36113_/CLK _34759_/D VGND VGND VPWR VPWR _34759_/Q sky130_fd_sc_hd__dfxtp_1
X_22773_ _35730_/Q _32241_/Q _35602_/Q _35538_/Q _20593_/X _20595_/X VGND VGND VPWR
+ VPWR _22773_/X sky130_fd_sc_hd__mux4_1
X_27300_ _27300_/A VGND VGND VPWR VPWR _34036_/D sky130_fd_sc_hd__clkbuf_1
X_24512_ _23064_/X _32783_/Q _24516_/S VGND VGND VPWR VPWR _24513_/A sky130_fd_sc_hd__mux2_1
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21724_ _33652_/Q _33588_/Q _33524_/Q _33460_/Q _21447_/X _21448_/X VGND VGND VPWR
+ VPWR _21724_/X sky130_fd_sc_hd__mux4_1
X_28280_ _27692_/X _34470_/Q _28286_/S VGND VGND VPWR VPWR _28281_/A sky130_fd_sc_hd__mux2_1
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25492_ _25540_/S VGND VGND VPWR VPWR _25511_/S sky130_fd_sc_hd__clkbuf_8
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27231_ _27231_/A VGND VGND VPWR VPWR _34005_/D sky130_fd_sc_hd__clkbuf_1
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24443_ _22962_/X _32750_/Q _24453_/S VGND VGND VPWR VPWR _24444_/A sky130_fd_sc_hd__mux2_1
X_21655_ _33394_/Q _33330_/Q _33266_/Q _33202_/Q _21374_/X _21375_/X VGND VGND VPWR
+ VPWR _21655_/X sky130_fd_sc_hd__mux4_1
XFILLER_200_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20606_ _22377_/A VGND VGND VPWR VPWR _22515_/A sky130_fd_sc_hd__buf_12
X_27162_ input36/X VGND VGND VPWR VPWR _27162_/X sky130_fd_sc_hd__buf_4
XFILLER_71_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24374_ _24374_/A VGND VGND VPWR VPWR _32717_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21586_ _33904_/Q _33840_/Q _33776_/Q _36080_/Q _21271_/X _21272_/X VGND VGND VPWR
+ VPWR _21586_/X sky130_fd_sc_hd__mux4_1
X_26113_ _24843_/X _33508_/Q _26123_/S VGND VGND VPWR VPWR _26114_/A sky130_fd_sc_hd__mux2_1
X_23325_ _32180_/Q _23243_/X _23335_/S VGND VGND VPWR VPWR _23326_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20537_ _33108_/Q _32084_/Q _35860_/Q _35796_/Q _18379_/X _18380_/X VGND VGND VPWR
+ VPWR _20537_/X sky130_fd_sc_hd__mux4_1
X_27093_ input11/X VGND VGND VPWR VPWR _27093_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_166_999 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26044_ _26044_/A VGND VGND VPWR VPWR _33475_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23256_ _32158_/Q _23255_/X _23259_/S VGND VGND VPWR VPWR _23257_/A sky130_fd_sc_hd__mux2_1
X_20468_ _19453_/A _20466_/X _20467_/X _19456_/A VGND VGND VPWR VPWR _20468_/X sky130_fd_sc_hd__a22o_1
XFILLER_101_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22207_ _22560_/A VGND VGND VPWR VPWR _22207_/X sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_161_CLK clkbuf_6_31__f_CLK/X VGND VGND VPWR VPWR _36115_/CLK sky130_fd_sc_hd__clkbuf_16
X_20399_ _33680_/Q _33616_/Q _33552_/Q _33488_/Q _20206_/X _20207_/X VGND VGND VPWR
+ VPWR _20399_/X sky130_fd_sc_hd__mux4_1
XFILLER_165_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23187_ _23187_/A VGND VGND VPWR VPWR _32131_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_885 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29803_ _35160_/Q _29336_/X _29817_/S VGND VGND VPWR VPWR _29804_/A sky130_fd_sc_hd__mux2_1
XTAP_6634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22138_ _21951_/X _22136_/X _22137_/X _21954_/X VGND VGND VPWR VPWR _22138_/X sky130_fd_sc_hd__a22o_1
XTAP_5900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27995_ _34335_/Q _27062_/X _27995_/S VGND VGND VPWR VPWR _27996_/A sky130_fd_sc_hd__mux2_1
XTAP_6645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26946_ _33900_/Q _23299_/X _26960_/S VGND VGND VPWR VPWR _26947_/A sky130_fd_sc_hd__mux2_1
X_29734_ _29734_/A VGND VGND VPWR VPWR _35127_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22069_ _35197_/Q _35133_/Q _35069_/Q _32253_/Q _21963_/X _21964_/X VGND VGND VPWR
+ VPWR _22069_/X sky130_fd_sc_hd__mux4_1
XFILLER_212_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29665_ _29665_/A VGND VGND VPWR VPWR _35094_/D sky130_fd_sc_hd__clkbuf_1
X_26877_ _26877_/A VGND VGND VPWR VPWR _33867_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_948 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16630_ _34150_/Q _34086_/Q _34022_/Q _33958_/Q _16387_/X _16388_/X VGND VGND VPWR
+ VPWR _16630_/X sky130_fd_sc_hd__mux4_1
X_28616_ _28616_/A VGND VGND VPWR VPWR _34629_/D sky130_fd_sc_hd__clkbuf_1
X_25828_ _24821_/X _33373_/Q _25832_/S VGND VGND VPWR VPWR _25829_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29596_ _35062_/Q _29429_/X _29610_/S VGND VGND VPWR VPWR _29597_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16561_ _16561_/A _16561_/B _16561_/C _16561_/D VGND VGND VPWR VPWR _16562_/A sky130_fd_sc_hd__or4_2
XFILLER_244_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25759_ _25759_/A VGND VGND VPWR VPWR _33340_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28547_ _28547_/A VGND VGND VPWR VPWR _34596_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18300_ _20073_/A VGND VGND VPWR VPWR _20164_/A sky130_fd_sc_hd__buf_12
XFILLER_71_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19280_ _19280_/A _19280_/B _19280_/C _19280_/D VGND VGND VPWR VPWR _19281_/A sky130_fd_sc_hd__or4_4
Xclkbuf_6_55__f_CLK clkbuf_5_27_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_55__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_28478_ _27785_/X _34564_/Q _28484_/S VGND VGND VPWR VPWR _28479_/A sky130_fd_sc_hd__mux2_1
X_16492_ _16492_/A VGND VGND VPWR VPWR _31969_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18231_ _17158_/A _18229_/X _18230_/X _17163_/A VGND VGND VPWR VPWR _18231_/X sky130_fd_sc_hd__a22o_1
X_27429_ _34098_/Q _27121_/X _27431_/S VGND VGND VPWR VPWR _27430_/A sky130_fd_sc_hd__mux2_1
X_18162_ _33426_/Q _33362_/Q _33298_/Q _33234_/Q _16037_/X _16039_/X VGND VGND VPWR
+ VPWR _18162_/X sky130_fd_sc_hd__mux4_1
X_30440_ _30440_/A VGND VGND VPWR VPWR _35462_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17113_ _17003_/X _17111_/X _17112_/X _17006_/X VGND VGND VPWR VPWR _17113_/X sky130_fd_sc_hd__a22o_1
XFILLER_128_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18093_ _34447_/Q _36175_/Q _34319_/Q _34255_/Q _17935_/X _17936_/X VGND VGND VPWR
+ VPWR _18093_/X sky130_fd_sc_hd__mux4_1
XFILLER_184_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30371_ _30371_/A VGND VGND VPWR VPWR _35429_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32110_ _32877_/CLK _32110_/D VGND VGND VPWR VPWR _32110_/Q sky130_fd_sc_hd__dfxtp_1
X_17044_ _35185_/Q _35121_/Q _35057_/Q _32198_/Q _17010_/X _17011_/X VGND VGND VPWR
+ VPWR _17044_/X sky130_fd_sc_hd__mux4_1
X_33090_ _36034_/CLK _33090_/D VGND VGND VPWR VPWR _33090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32041_ _35753_/CLK _32041_/D VGND VGND VPWR VPWR _32041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_152_CLK clkbuf_6_29__f_CLK/X VGND VGND VPWR VPWR _36180_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_217_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18995_ _18752_/X _18993_/X _18994_/X _18757_/X VGND VGND VPWR VPWR _18995_/X sky130_fd_sc_hd__a22o_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35800_ _35800_/CLK _35800_/D VGND VGND VPWR VPWR _35800_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17946_ _33419_/Q _33355_/Q _33291_/Q _33227_/Q _17833_/X _17834_/X VGND VGND VPWR
+ VPWR _17946_/X sky130_fd_sc_hd__mux4_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33992_ _34121_/CLK _33992_/D VGND VGND VPWR VPWR _33992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35731_ _35731_/CLK _35731_/D VGND VGND VPWR VPWR _35731_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32943_ _36015_/CLK _32943_/D VGND VGND VPWR VPWR _32943_/Q sky130_fd_sc_hd__dfxtp_1
X_17877_ _17552_/X _17875_/X _17876_/X _17557_/X VGND VGND VPWR VPWR _17877_/X sky130_fd_sc_hd__a22o_1
XFILLER_38_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19616_ _19612_/X _19615_/X _19440_/X _19441_/X VGND VGND VPWR VPWR _19633_/B sky130_fd_sc_hd__o211a_1
X_35662_ _35663_/CLK _35662_/D VGND VGND VPWR VPWR _35662_/Q sky130_fd_sc_hd__dfxtp_1
X_16828_ _16714_/X _16826_/X _16827_/X _16718_/X VGND VGND VPWR VPWR _16828_/X sky130_fd_sc_hd__a22o_1
X_32874_ _32875_/CLK _32874_/D VGND VGND VPWR VPWR _32874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34613_ _36024_/CLK _34613_/D VGND VGND VPWR VPWR _34613_/Q sky130_fd_sc_hd__dfxtp_1
X_31825_ _23225_/X _36118_/Q _31843_/S VGND VGND VPWR VPWR _31826_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_1081 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19547_ _32119_/Q _32311_/Q _32375_/Q _35895_/Q _19227_/X _19368_/X VGND VGND VPWR
+ VPWR _19547_/X sky130_fd_sc_hd__mux4_1
X_35593_ _35722_/CLK _35593_/D VGND VGND VPWR VPWR _35593_/Q sky130_fd_sc_hd__dfxtp_1
X_16759_ _33065_/Q _32041_/Q _35817_/Q _35753_/Q _16725_/X _16726_/X VGND VGND VPWR
+ VPWR _16759_/X sky130_fd_sc_hd__mux4_1
XFILLER_206_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34544_ _36143_/CLK _34544_/D VGND VGND VPWR VPWR _34544_/Q sky130_fd_sc_hd__dfxtp_1
X_31756_ _31756_/A VGND VGND VPWR VPWR _36085_/D sky130_fd_sc_hd__clkbuf_1
X_19478_ _19359_/X _19476_/X _19477_/X _19365_/X VGND VGND VPWR VPWR _19478_/X sky130_fd_sc_hd__a22o_1
XFILLER_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18429_ _18360_/X _18427_/X _18428_/X _18372_/X VGND VGND VPWR VPWR _18429_/X sky130_fd_sc_hd__a22o_1
X_30707_ _35589_/Q _29475_/X _30711_/S VGND VGND VPWR VPWR _30708_/A sky130_fd_sc_hd__mux2_1
X_34475_ _35820_/CLK _34475_/D VGND VGND VPWR VPWR _34475_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31687_ _31687_/A VGND VGND VPWR VPWR _36053_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_222_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36214_ _36219_/CLK _36214_/D VGND VGND VPWR VPWR _36214_/Q sky130_fd_sc_hd__dfxtp_1
X_33426_ _36115_/CLK _33426_/D VGND VGND VPWR VPWR _33426_/Q sky130_fd_sc_hd__dfxtp_1
X_21440_ _34411_/Q _36139_/Q _34283_/Q _34219_/Q _21123_/X _21124_/X VGND VGND VPWR
+ VPWR _21440_/X sky130_fd_sc_hd__mux4_1
XFILLER_147_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30638_ _35556_/Q _29373_/X _30648_/S VGND VGND VPWR VPWR _30639_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_222_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21371_ _33642_/Q _33578_/Q _33514_/Q _33450_/Q _21094_/X _21095_/X VGND VGND VPWR
+ VPWR _21371_/X sky130_fd_sc_hd__mux4_1
X_36145_ _36147_/CLK _36145_/D VGND VGND VPWR VPWR _36145_/Q sky130_fd_sc_hd__dfxtp_1
X_33357_ _34186_/CLK _33357_/D VGND VGND VPWR VPWR _33357_/Q sky130_fd_sc_hd__dfxtp_1
X_30569_ _30569_/A VGND VGND VPWR VPWR _35523_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_391_CLK clkbuf_6_40__f_CLK/X VGND VGND VPWR VPWR _33910_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_175_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20322_ _20318_/X _20321_/X _20146_/X _20147_/X VGND VGND VPWR VPWR _20337_/B sky130_fd_sc_hd__o211a_1
X_23110_ _22915_/X _32095_/Q _23110_/S VGND VGND VPWR VPWR _23111_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32308_ _32882_/CLK _32308_/D VGND VGND VPWR VPWR _32308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24090_ _24090_/A VGND VGND VPWR VPWR _32585_/D sky130_fd_sc_hd__clkbuf_1
X_36076_ _36076_/CLK _36076_/D VGND VGND VPWR VPWR _36076_/Q sky130_fd_sc_hd__dfxtp_1
X_33288_ _33420_/CLK _33288_/D VGND VGND VPWR VPWR _33288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35027_ _35729_/CLK _35027_/D VGND VGND VPWR VPWR _35027_/Q sky130_fd_sc_hd__dfxtp_1
X_23041_ _23041_/A VGND VGND VPWR VPWR _32071_/D sky130_fd_sc_hd__clkbuf_1
X_20253_ _32139_/Q _32331_/Q _32395_/Q _35915_/Q _19933_/X _20074_/X VGND VGND VPWR
+ VPWR _20253_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_143_CLK clkbuf_6_28__f_CLK/X VGND VGND VPWR VPWR _35990_/CLK sky130_fd_sc_hd__clkbuf_16
X_32239_ _35728_/CLK _32239_/D VGND VGND VPWR VPWR _32239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20184_ _20065_/X _20182_/X _20183_/X _20071_/X VGND VGND VPWR VPWR _20184_/X sky130_fd_sc_hd__a22o_1
XFILLER_192_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26800_ _33831_/Q _23283_/X _26804_/S VGND VGND VPWR VPWR _26801_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27780_ _27779_/X _34242_/Q _27795_/S VGND VGND VPWR VPWR _27781_/A sky130_fd_sc_hd__mux2_1
X_24992_ _24991_/X _32980_/Q _24995_/S VGND VGND VPWR VPWR _24993_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26731_ _26731_/A VGND VGND VPWR VPWR _33798_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35929_ _35929_/CLK _35929_/D VGND VGND VPWR VPWR _35929_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23943_ _23943_/A VGND VGND VPWR VPWR _32516_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29450_ input33/X VGND VGND VPWR VPWR _29450_/X sky130_fd_sc_hd__buf_2
XFILLER_245_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26662_ _26662_/A VGND VGND VPWR VPWR _33765_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_986 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23874_ _23874_/A VGND VGND VPWR VPWR _32483_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_217_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28401_ _28401_/A VGND VGND VPWR VPWR _34527_/D sky130_fd_sc_hd__clkbuf_1
X_25613_ _24902_/X _33271_/Q _25625_/S VGND VGND VPWR VPWR _25614_/A sky130_fd_sc_hd__mux2_1
X_22825_ _22821_/X _22824_/X _22438_/A VGND VGND VPWR VPWR _22847_/A sky130_fd_sc_hd__o21ba_1
X_29381_ _29381_/A VGND VGND VPWR VPWR _34982_/D sky130_fd_sc_hd__clkbuf_1
X_26593_ _24951_/X _33735_/Q _26593_/S VGND VGND VPWR VPWR _26594_/A sky130_fd_sc_hd__mux2_1
XFILLER_198_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28332_ _28332_/A VGND VGND VPWR VPWR _34494_/D sky130_fd_sc_hd__clkbuf_1
X_25544_ _24796_/X _33238_/Q _25562_/S VGND VGND VPWR VPWR _25545_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22756_ _22752_/X _22755_/X _22471_/X VGND VGND VPWR VPWR _22757_/D sky130_fd_sc_hd__o21ba_1
XFILLER_213_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28263_ _27667_/X _34462_/Q _28265_/S VGND VGND VPWR VPWR _28264_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21707_ _21703_/X _21706_/X _21387_/X _21388_/X VGND VGND VPWR VPWR _21722_/B sky130_fd_sc_hd__o211a_1
XFILLER_129_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25475_ _25475_/A VGND VGND VPWR VPWR _33205_/D sky130_fd_sc_hd__clkbuf_1
X_22687_ _33103_/Q _32079_/Q _35855_/Q _35791_/Q _22384_/X _22385_/X VGND VGND VPWR
+ VPWR _22687_/X sky130_fd_sc_hd__mux4_1
X_27214_ input54/X VGND VGND VPWR VPWR _27214_/X sky130_fd_sc_hd__buf_4
XFILLER_157_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24426_ _22937_/X _32742_/Q _24432_/S VGND VGND VPWR VPWR _24427_/A sky130_fd_sc_hd__mux2_1
X_21638_ _21598_/X _21636_/X _21637_/X _21601_/X VGND VGND VPWR VPWR _21638_/X sky130_fd_sc_hd__a22o_1
X_28194_ _28194_/A VGND VGND VPWR VPWR _34429_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27145_ _27145_/A VGND VGND VPWR VPWR _33977_/D sky130_fd_sc_hd__clkbuf_1
X_24357_ _24357_/A VGND VGND VPWR VPWR _32709_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_382_CLK clkbuf_6_42__f_CLK/X VGND VGND VPWR VPWR _36092_/CLK sky130_fd_sc_hd__clkbuf_16
X_21569_ _35439_/Q _35375_/Q _35311_/Q _35247_/Q _21501_/X _21502_/X VGND VGND VPWR
+ VPWR _21569_/X sky130_fd_sc_hd__mux4_1
XFILLER_197_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23308_ input88/X input87/X input86/X VGND VGND VPWR VPWR _23309_/A sky130_fd_sc_hd__or3b_1
XFILLER_126_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27076_ _33955_/Q _27075_/X _27094_/S VGND VGND VPWR VPWR _27077_/A sky130_fd_sc_hd__mux2_1
X_24288_ _24288_/A VGND VGND VPWR VPWR _32676_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26027_ _26027_/A VGND VGND VPWR VPWR _33467_/D sky130_fd_sc_hd__clkbuf_1
XTAP_7110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_134_CLK clkbuf_6_23__f_CLK/X VGND VGND VPWR VPWR _34585_/CLK sky130_fd_sc_hd__clkbuf_16
X_23239_ _23239_/A VGND VGND VPWR VPWR _32152_/D sky130_fd_sc_hd__clkbuf_1
XTAP_7121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17800_ _17800_/A VGND VGND VPWR VPWR _17800_/X sky130_fd_sc_hd__buf_4
XTAP_6453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15992_ _16061_/A VGND VGND VPWR VPWR _17799_/A sky130_fd_sc_hd__buf_12
XTAP_6464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18780_ _35425_/Q _35361_/Q _35297_/Q _35233_/Q _18495_/X _18496_/X VGND VGND VPWR
+ VPWR _18780_/X sky130_fd_sc_hd__mux4_1
XTAP_6475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27978_ _27978_/A VGND VGND VPWR VPWR _34326_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17731_ _17851_/A VGND VGND VPWR VPWR _17731_/X sky130_fd_sc_hd__buf_4
XTAP_5763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29717_ _29717_/A VGND VGND VPWR VPWR _35119_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26929_ _33892_/Q _23274_/X _26939_/S VGND VGND VPWR VPWR _26930_/A sky130_fd_sc_hd__mux2_1
XTAP_5785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29648_ _35087_/Q _29506_/X _29652_/S VGND VGND VPWR VPWR _29649_/A sky130_fd_sc_hd__mux2_1
X_17662_ _17658_/X _17661_/X _17485_/X VGND VGND VPWR VPWR _17686_/A sky130_fd_sc_hd__o21ba_1
XFILLER_48_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_907 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19401_ _32627_/Q _32563_/Q _32499_/Q _35955_/Q _19223_/X _19360_/X VGND VGND VPWR
+ VPWR _19401_/X sky130_fd_sc_hd__mux4_1
X_16613_ _35685_/Q _32192_/Q _35557_/Q _35493_/Q _16611_/X _16612_/X VGND VGND VPWR
+ VPWR _16613_/X sky130_fd_sc_hd__mux4_2
XFILLER_63_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17593_ _33409_/Q _33345_/Q _33281_/Q _33217_/Q _17480_/X _17481_/X VGND VGND VPWR
+ VPWR _17593_/X sky130_fd_sc_hd__mux4_1
XFILLER_169_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29579_ _35054_/Q _29404_/X _29589_/S VGND VGND VPWR VPWR _29580_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31610_ _31610_/A VGND VGND VPWR VPWR _36016_/D sky130_fd_sc_hd__clkbuf_1
X_19332_ _32113_/Q _32305_/Q _32369_/Q _35889_/Q _19227_/X _19015_/X VGND VGND VPWR
+ VPWR _19332_/X sky130_fd_sc_hd__mux4_1
X_16544_ _16540_/X _16543_/X _16434_/X _16435_/X VGND VGND VPWR VPWR _16561_/B sky130_fd_sc_hd__o211a_1
X_32590_ _35982_/CLK _32590_/D VGND VGND VPWR VPWR _32590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31541_ _27822_/X _35984_/Q _31543_/S VGND VGND VPWR VPWR _31542_/A sky130_fd_sc_hd__mux2_1
X_16475_ _16361_/X _16473_/X _16474_/X _16365_/X VGND VGND VPWR VPWR _16475_/X sky130_fd_sc_hd__a22o_1
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19263_ _19259_/X _19262_/X _19087_/X _19088_/X VGND VGND VPWR VPWR _19280_/B sky130_fd_sc_hd__o211a_1
XFILLER_188_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18214_ _34963_/Q _34899_/Q _34835_/Q _34771_/Q _16083_/X _16085_/X VGND VGND VPWR
+ VPWR _18214_/X sky130_fd_sc_hd__mux4_1
X_34260_ _36181_/CLK _34260_/D VGND VGND VPWR VPWR _34260_/Q sky130_fd_sc_hd__dfxtp_1
X_31472_ _27720_/X _35951_/Q _31480_/S VGND VGND VPWR VPWR _31473_/A sky130_fd_sc_hd__mux2_1
X_19194_ _32109_/Q _32301_/Q _32365_/Q _35885_/Q _18874_/X _19015_/X VGND VGND VPWR
+ VPWR _19194_/X sky130_fd_sc_hd__mux4_1
XFILLER_54_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30423_ _35454_/Q _29453_/X _30441_/S VGND VGND VPWR VPWR _30424_/A sky130_fd_sc_hd__mux2_1
X_33211_ _33531_/CLK _33211_/D VGND VGND VPWR VPWR _33211_/Q sky130_fd_sc_hd__dfxtp_1
X_18145_ _15981_/X _18143_/X _18144_/X _15991_/X VGND VGND VPWR VPWR _18145_/X sky130_fd_sc_hd__a22o_1
X_34191_ _34192_/CLK _34191_/D VGND VGND VPWR VPWR _34191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_373_CLK clkbuf_6_43__f_CLK/X VGND VGND VPWR VPWR _36157_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_200_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30354_ _30354_/A VGND VGND VPWR VPWR _35421_/D sky130_fd_sc_hd__clkbuf_1
X_18076_ _32655_/Q _32591_/Q _32527_/Q _35983_/Q _17982_/X _17766_/X VGND VGND VPWR
+ VPWR _18076_/X sky130_fd_sc_hd__mux4_1
X_33142_ _34485_/CLK _33142_/D VGND VGND VPWR VPWR _33142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17027_ _16853_/X _17023_/X _17026_/X _16856_/X VGND VGND VPWR VPWR _17027_/X sky130_fd_sc_hd__a22o_1
X_33073_ _36147_/CLK _33073_/D VGND VGND VPWR VPWR _33073_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_125_CLK clkbuf_6_21__f_CLK/X VGND VGND VPWR VPWR _36245_/CLK sky130_fd_sc_hd__clkbuf_16
X_30285_ _35389_/Q _29450_/X _30285_/S VGND VGND VPWR VPWR _30286_/A sky130_fd_sc_hd__mux2_1
XFILLER_131_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32024_ _35735_/CLK _32024_/D VGND VGND VPWR VPWR _32024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18978_ _18653_/X _18976_/X _18977_/X _18659_/X VGND VGND VPWR VPWR _18978_/X sky130_fd_sc_hd__a22o_1
XFILLER_85_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17929_ _33098_/Q _32074_/Q _35850_/Q _35786_/Q _17784_/X _17785_/X VGND VGND VPWR
+ VPWR _17929_/X sky130_fd_sc_hd__mux4_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33975_ _35703_/CLK _33975_/D VGND VGND VPWR VPWR _33975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35714_ _36033_/CLK _35714_/D VGND VGND VPWR VPWR _35714_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20940_ _34397_/Q _36125_/Q _34269_/Q _34205_/Q _20770_/X _20771_/X VGND VGND VPWR
+ VPWR _20940_/X sky130_fd_sc_hd__mux4_1
X_32926_ _35999_/CLK _32926_/D VGND VGND VPWR VPWR _32926_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_1059 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35645_ _35645_/CLK _35645_/D VGND VGND VPWR VPWR _35645_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20871_ _34907_/Q _34843_/Q _34779_/Q _34715_/Q _20696_/X _20698_/X VGND VGND VPWR
+ VPWR _20871_/X sky130_fd_sc_hd__mux4_1
X_32857_ _35733_/CLK _32857_/D VGND VGND VPWR VPWR _32857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22610_ _34189_/Q _34125_/Q _34061_/Q _33997_/Q _22399_/X _22400_/X VGND VGND VPWR
+ VPWR _22610_/X sky130_fd_sc_hd__mux4_1
XFILLER_228_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31808_ _31808_/A VGND VGND VPWR VPWR _36110_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_223_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23590_ _23590_/A VGND VGND VPWR VPWR _32287_/D sky130_fd_sc_hd__clkbuf_1
X_35576_ _35768_/CLK _35576_/D VGND VGND VPWR VPWR _35576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32788_ _32869_/CLK _32788_/D VGND VGND VPWR VPWR _32788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22541_ _22541_/A _22541_/B _22541_/C _22541_/D VGND VGND VPWR VPWR _22542_/A sky130_fd_sc_hd__or4_4
X_34527_ _35544_/CLK _34527_/D VGND VGND VPWR VPWR _34527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31739_ _31739_/A VGND VGND VPWR VPWR _36077_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25260_ _25260_/A VGND VGND VPWR VPWR _33105_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22472_ _22463_/X _22470_/X _22471_/X VGND VGND VPWR VPWR _22473_/D sky130_fd_sc_hd__o21ba_1
X_34458_ _34654_/CLK _34458_/D VGND VGND VPWR VPWR _34458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24211_ _24211_/A VGND VGND VPWR VPWR _32641_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33409_ _33924_/CLK _33409_/D VGND VGND VPWR VPWR _33409_/Q sky130_fd_sc_hd__dfxtp_1
X_21423_ _32619_/Q _32555_/Q _32491_/Q _35947_/Q _21170_/X _21307_/X VGND VGND VPWR
+ VPWR _21423_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_364_CLK clkbuf_6_44__f_CLK/X VGND VGND VPWR VPWR _35191_/CLK sky130_fd_sc_hd__clkbuf_16
X_25191_ _25191_/A VGND VGND VPWR VPWR _33072_/D sky130_fd_sc_hd__clkbuf_1
X_34389_ _35733_/CLK _34389_/D VGND VGND VPWR VPWR _34389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_1294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24142_ _24142_/A VGND VGND VPWR VPWR _32608_/D sky130_fd_sc_hd__clkbuf_1
X_36128_ _36128_/CLK _36128_/D VGND VGND VPWR VPWR _36128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21354_ _21350_/X _21353_/X _21034_/X _21035_/X VGND VGND VPWR VPWR _21369_/B sky130_fd_sc_hd__o211a_1
X_20305_ _20164_/X _20303_/X _20304_/X _20169_/X VGND VGND VPWR VPWR _20305_/X sky130_fd_sc_hd__a22o_1
XFILLER_123_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_116_CLK clkbuf_6_20__f_CLK/X VGND VGND VPWR VPWR _36219_/CLK sky130_fd_sc_hd__clkbuf_16
X_36059_ _36059_/CLK _36059_/D VGND VGND VPWR VPWR _36059_/Q sky130_fd_sc_hd__dfxtp_1
X_24073_ _24073_/A VGND VGND VPWR VPWR _32577_/D sky130_fd_sc_hd__clkbuf_1
X_28950_ _34786_/Q _27072_/X _28964_/S VGND VGND VPWR VPWR _28951_/A sky130_fd_sc_hd__mux2_1
X_21285_ _21245_/X _21283_/X _21284_/X _21248_/X VGND VGND VPWR VPWR _21285_/X sky130_fd_sc_hd__a22o_1
X_23024_ input39/X VGND VGND VPWR VPWR _23024_/X sky130_fd_sc_hd__buf_2
XFILLER_122_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27901_ _27901_/A VGND VGND VPWR VPWR _34290_/D sky130_fd_sc_hd__clkbuf_1
X_20236_ _20236_/A VGND VGND VPWR VPWR _20236_/X sky130_fd_sc_hd__buf_4
XFILLER_235_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28881_ _28881_/A VGND VGND VPWR VPWR _34753_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27832_ _27831_/X _34259_/Q _27838_/S VGND VGND VPWR VPWR _27833_/A sky130_fd_sc_hd__mux2_1
X_20167_ _20167_/A VGND VGND VPWR VPWR _20167_/X sky130_fd_sc_hd__clkbuf_4
XTAP_5015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20098_ _33671_/Q _33607_/Q _33543_/Q _33479_/Q _19853_/X _19854_/X VGND VGND VPWR
+ VPWR _20098_/X sky130_fd_sc_hd__mux4_1
X_24975_ _24975_/A VGND VGND VPWR VPWR _32974_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27763_ input33/X VGND VGND VPWR VPWR _27763_/X sky130_fd_sc_hd__clkbuf_4
XTAP_4336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_218_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29502_ _29502_/A VGND VGND VPWR VPWR _35021_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26714_ _33790_/Q _23420_/X _26732_/S VGND VGND VPWR VPWR _26715_/A sky130_fd_sc_hd__mux2_1
XTAP_3624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23926_ _23926_/A VGND VGND VPWR VPWR _32508_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27694_ _27694_/A VGND VGND VPWR VPWR _34214_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26645_ _26645_/A VGND VGND VPWR VPWR _33757_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29433_ _34999_/Q _29432_/X _29451_/S VGND VGND VPWR VPWR _29434_/A sky130_fd_sc_hd__mux2_1
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23857_ _23857_/A VGND VGND VPWR VPWR _32475_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22808_ _20601_/X _22806_/X _22807_/X _20607_/X VGND VGND VPWR VPWR _22808_/X sky130_fd_sc_hd__a22o_1
XFILLER_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26576_ _26576_/A VGND VGND VPWR VPWR _33726_/D sky130_fd_sc_hd__clkbuf_1
X_29364_ input3/X VGND VGND VPWR VPWR _29364_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23788_ _23005_/X _32380_/Q _23790_/S VGND VGND VPWR VPWR _23789_/A sky130_fd_sc_hd__mux2_1
XFILLER_246_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25527_ _25527_/A VGND VGND VPWR VPWR _33230_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28315_ _28315_/A VGND VGND VPWR VPWR _34486_/D sky130_fd_sc_hd__clkbuf_1
X_29295_ _34950_/Q _27183_/X _29297_/S VGND VGND VPWR VPWR _29296_/A sky130_fd_sc_hd__mux2_1
X_22739_ _32145_/Q _32337_/Q _32401_/Q _35921_/Q _22586_/X _21611_/A VGND VGND VPWR
+ VPWR _22739_/X sky130_fd_sc_hd__mux4_1
XFILLER_41_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28246_ _28378_/S VGND VGND VPWR VPWR _28265_/S sky130_fd_sc_hd__buf_6
XFILLER_186_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16260_ _35675_/Q _32181_/Q _35547_/Q _35483_/Q _16258_/X _16259_/X VGND VGND VPWR
+ VPWR _16260_/X sky130_fd_sc_hd__mux4_1
X_25458_ _25458_/A VGND VGND VPWR VPWR _33197_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24409_ _22912_/X _32734_/Q _24411_/S VGND VGND VPWR VPWR _24410_/A sky130_fd_sc_hd__mux2_1
X_16191_ _16187_/X _16190_/X _16044_/X _16046_/X VGND VGND VPWR VPWR _16208_/B sky130_fd_sc_hd__o211a_1
XFILLER_187_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28177_ _27739_/X _34421_/Q _28193_/S VGND VGND VPWR VPWR _28178_/A sky130_fd_sc_hd__mux2_1
X_25389_ _33166_/Q _23475_/X _25395_/S VGND VGND VPWR VPWR _25390_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_355_CLK clkbuf_6_46__f_CLK/X VGND VGND VPWR VPWR _35709_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_51_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27128_ _27230_/S VGND VGND VPWR VPWR _27156_/S sky130_fd_sc_hd__buf_4
XFILLER_86_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_1378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19950_ _34434_/Q _36162_/Q _34306_/Q _34242_/Q _19882_/X _19883_/X VGND VGND VPWR
+ VPWR _19950_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_107_CLK clkbuf_leaf_81_CLK/A VGND VGND VPWR VPWR _35802_/CLK sky130_fd_sc_hd__clkbuf_16
X_27059_ input63/X VGND VGND VPWR VPWR _27059_/X sky130_fd_sc_hd__buf_4
XFILLER_218_1410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18901_ _33893_/Q _33829_/Q _33765_/Q _36069_/Q _18618_/X _18619_/X VGND VGND VPWR
+ VPWR _18901_/X sky130_fd_sc_hd__mux4_1
X_30070_ _30070_/A VGND VGND VPWR VPWR _35286_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_206_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19881_ _19806_/X _19879_/X _19880_/X _19809_/X VGND VGND VPWR VPWR _19881_/X sky130_fd_sc_hd__a22o_1
XFILLER_175_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18832_ _34147_/Q _34083_/Q _34019_/Q _33955_/Q _18687_/X _18688_/X VGND VGND VPWR
+ VPWR _18832_/X sky130_fd_sc_hd__mux4_1
XFILLER_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18763_ _33633_/Q _33569_/Q _33505_/Q _33441_/Q _18441_/X _18442_/X VGND VGND VPWR
+ VPWR _18763_/X sky130_fd_sc_hd__mux4_1
XTAP_5560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17714_ _17708_/X _17713_/X _17504_/X VGND VGND VPWR VPWR _17724_/C sky130_fd_sc_hd__o21ba_1
XFILLER_236_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33760_ _36065_/CLK _33760_/D VGND VGND VPWR VPWR _33760_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30972_ _30972_/A VGND VGND VPWR VPWR _35714_/D sky130_fd_sc_hd__clkbuf_1
X_18694_ _18690_/X _18693_/X _18315_/X VGND VGND VPWR VPWR _18716_/A sky130_fd_sc_hd__o21ba_1
XFILLER_209_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32711_ _32905_/CLK _32711_/D VGND VGND VPWR VPWR _32711_/Q sky130_fd_sc_hd__dfxtp_1
X_17645_ _17998_/A VGND VGND VPWR VPWR _17645_/X sky130_fd_sc_hd__buf_6
X_33691_ _36057_/CLK _33691_/D VGND VGND VPWR VPWR _33691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_940 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35430_ _35685_/CLK _35430_/D VGND VGND VPWR VPWR _35430_/Q sky130_fd_sc_hd__dfxtp_1
X_32642_ _36034_/CLK _32642_/D VGND VGND VPWR VPWR _32642_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17576_ _33088_/Q _32064_/Q _35840_/Q _35776_/Q _17431_/X _17432_/X VGND VGND VPWR
+ VPWR _17576_/X sky130_fd_sc_hd__mux4_1
X_19315_ _34928_/Q _34864_/Q _34800_/Q _34736_/Q _19107_/X _19108_/X VGND VGND VPWR
+ VPWR _19315_/X sky130_fd_sc_hd__mux4_1
XFILLER_17_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16527_ _16452_/X _16525_/X _16526_/X _16457_/X VGND VGND VPWR VPWR _16527_/X sky130_fd_sc_hd__a22o_1
X_35361_ _36005_/CLK _35361_/D VGND VGND VPWR VPWR _35361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_1046 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32573_ _35965_/CLK _32573_/D VGND VGND VPWR VPWR _32573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34312_ _36171_/CLK _34312_/D VGND VGND VPWR VPWR _34312_/Q sky130_fd_sc_hd__dfxtp_1
X_31524_ _31551_/S VGND VGND VPWR VPWR _31543_/S sky130_fd_sc_hd__buf_4
X_19246_ _19105_/X _19244_/X _19245_/X _19110_/X VGND VGND VPWR VPWR _19246_/X sky130_fd_sc_hd__a22o_1
X_35292_ _35804_/CLK _35292_/D VGND VGND VPWR VPWR _35292_/Q sky130_fd_sc_hd__dfxtp_1
X_16458_ _16452_/X _16453_/X _16456_/X _16457_/X VGND VGND VPWR VPWR _16458_/X sky130_fd_sc_hd__a22o_1
XFILLER_121_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34243_ _36164_/CLK _34243_/D VGND VGND VPWR VPWR _34243_/Q sky130_fd_sc_hd__dfxtp_1
X_16389_ _34143_/Q _34079_/Q _34015_/Q _33951_/Q _16387_/X _16388_/X VGND VGND VPWR
+ VPWR _16389_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_346_CLK clkbuf_6_47__f_CLK/X VGND VGND VPWR VPWR _32575_/CLK sky130_fd_sc_hd__clkbuf_16
X_19177_ _19177_/A VGND VGND VPWR VPWR _19177_/X sky130_fd_sc_hd__buf_4
X_31455_ _27695_/X _35943_/Q _31459_/S VGND VGND VPWR VPWR _31456_/A sky130_fd_sc_hd__mux2_1
XFILLER_223_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18128_ _18128_/A VGND VGND VPWR VPWR _32016_/D sky130_fd_sc_hd__buf_2
XFILLER_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30406_ _35446_/Q _29429_/X _30420_/S VGND VGND VPWR VPWR _30407_/A sky130_fd_sc_hd__mux2_1
XFILLER_247_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31386_ _31386_/A VGND VGND VPWR VPWR _35910_/D sky130_fd_sc_hd__clkbuf_1
X_34174_ _34174_/CLK _34174_/D VGND VGND VPWR VPWR _34174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33125_ _36007_/CLK _33125_/D VGND VGND VPWR VPWR _33125_/Q sky130_fd_sc_hd__dfxtp_1
X_18059_ _18055_/X _18058_/X _17857_/X VGND VGND VPWR VPWR _18067_/C sky130_fd_sc_hd__o21ba_1
X_30337_ _30337_/A _30877_/A VGND VGND VPWR VPWR _30470_/S sky130_fd_sc_hd__nor2_8
XFILLER_144_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21070_ _32609_/Q _32545_/Q _32481_/Q _35937_/Q _20817_/X _20954_/X VGND VGND VPWR
+ VPWR _21070_/X sky130_fd_sc_hd__mux4_1
XFILLER_67_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30268_ _30268_/A VGND VGND VPWR VPWR _35380_/D sky130_fd_sc_hd__clkbuf_1
X_33056_ _35810_/CLK _33056_/D VGND VGND VPWR VPWR _33056_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_1270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20021_ _34948_/Q _34884_/Q _34820_/Q _34756_/Q _19813_/X _19814_/X VGND VGND VPWR
+ VPWR _20021_/X sky130_fd_sc_hd__mux4_1
XFILLER_86_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32007_ _36209_/CLK _32007_/D VGND VGND VPWR VPWR _32007_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_232_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30199_ _30199_/A VGND VGND VPWR VPWR _35348_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_1279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24760_ _24760_/A VGND VGND VPWR VPWR _32900_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33958_ _34085_/CLK _33958_/D VGND VGND VPWR VPWR _33958_/Q sky130_fd_sc_hd__dfxtp_1
X_21972_ _21972_/A VGND VGND VPWR VPWR _36218_/D sky130_fd_sc_hd__buf_2
XFILLER_27_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23711_ _22891_/X _32343_/Q _23727_/S VGND VGND VPWR VPWR _23712_/A sky130_fd_sc_hd__mux2_1
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20923_ _32605_/Q _32541_/Q _32477_/Q _35933_/Q _20817_/X _22317_/A VGND VGND VPWR
+ VPWR _20923_/X sky130_fd_sc_hd__mux4_1
X_32909_ _32909_/CLK _32909_/D VGND VGND VPWR VPWR _32909_/Q sky130_fd_sc_hd__dfxtp_1
X_24691_ _24691_/A VGND VGND VPWR VPWR _32867_/D sky130_fd_sc_hd__clkbuf_1
X_33889_ _35618_/CLK _33889_/D VGND VGND VPWR VPWR _33889_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26430_ _33658_/Q _23408_/X _26436_/S VGND VGND VPWR VPWR _26431_/A sky130_fd_sc_hd__mux2_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35628_ _35693_/CLK _35628_/D VGND VGND VPWR VPWR _35628_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23642_ _22993_/X _32312_/Q _23652_/S VGND VGND VPWR VPWR _23643_/A sky130_fd_sc_hd__mux2_1
X_20854_ _32091_/Q _32283_/Q _32347_/Q _35867_/Q _20821_/X _22467_/A VGND VGND VPWR
+ VPWR _20854_/X sky130_fd_sc_hd__mux4_1
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26361_ _33625_/Q _23240_/X _26373_/S VGND VGND VPWR VPWR _26362_/A sky130_fd_sc_hd__mux2_1
XFILLER_223_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23573_ _22891_/X _32279_/Q _23589_/S VGND VGND VPWR VPWR _23574_/A sky130_fd_sc_hd__mux2_1
X_35559_ _35559_/CLK _35559_/D VGND VGND VPWR VPWR _35559_/Q sky130_fd_sc_hd__dfxtp_1
X_20785_ _32601_/Q _32537_/Q _32473_/Q _35929_/Q _22466_/A _22317_/A VGND VGND VPWR
+ VPWR _20785_/X sky130_fd_sc_hd__mux4_1
X_28100_ _34385_/Q _27217_/X _28100_/S VGND VGND VPWR VPWR _28101_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25312_ _25312_/A VGND VGND VPWR VPWR _33129_/D sky130_fd_sc_hd__clkbuf_1
X_22524_ _22520_/X _22523_/X _22446_/X _22447_/X VGND VGND VPWR VPWR _22541_/B sky130_fd_sc_hd__o211a_2
X_29080_ _29191_/S VGND VGND VPWR VPWR _29099_/S sky130_fd_sc_hd__buf_4
XFILLER_194_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26292_ _24908_/X _33593_/Q _26300_/S VGND VGND VPWR VPWR _26293_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28031_ _34352_/Q _27115_/X _28037_/S VGND VGND VPWR VPWR _28032_/A sky130_fd_sc_hd__mux2_1
X_25243_ _33097_/Q _23460_/X _25259_/S VGND VGND VPWR VPWR _25244_/A sky130_fd_sc_hd__mux2_1
X_22455_ _33096_/Q _32072_/Q _35848_/Q _35784_/Q _22384_/X _22385_/X VGND VGND VPWR
+ VPWR _22455_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_337_CLK clkbuf_6_45__f_CLK/X VGND VGND VPWR VPWR _35962_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_183_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21406_ _34410_/Q _36138_/Q _34282_/Q _34218_/Q _21123_/X _21124_/X VGND VGND VPWR
+ VPWR _21406_/X sky130_fd_sc_hd__mux4_1
XFILLER_202_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25174_ _25174_/A VGND VGND VPWR VPWR _33064_/D sky130_fd_sc_hd__clkbuf_1
X_22386_ _33094_/Q _32070_/Q _35846_/Q _35782_/Q _22384_/X _22385_/X VGND VGND VPWR
+ VPWR _22386_/X sky130_fd_sc_hd__mux4_1
XFILLER_159_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24125_ _24125_/A VGND VGND VPWR VPWR _32600_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21337_ _21337_/A _21337_/B _21337_/C _21337_/D VGND VGND VPWR VPWR _21338_/A sky130_fd_sc_hd__or4_4
X_29982_ _35245_/Q _29401_/X _29994_/S VGND VGND VPWR VPWR _29983_/A sky130_fd_sc_hd__mux2_1
X_28933_ _34778_/Q _27047_/X _28943_/S VGND VGND VPWR VPWR _28934_/A sky130_fd_sc_hd__mux2_1
X_24056_ _24056_/A VGND VGND VPWR VPWR _32569_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21268_ _34151_/Q _34087_/Q _34023_/Q _33959_/Q _20987_/X _20988_/X VGND VGND VPWR
+ VPWR _21268_/X sky130_fd_sc_hd__mux4_2
XFILLER_137_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23007_ _23007_/A VGND VGND VPWR VPWR _32060_/D sky130_fd_sc_hd__clkbuf_1
X_20219_ _33162_/Q _36042_/Q _33034_/Q _32970_/Q _20068_/X _20069_/X VGND VGND VPWR
+ VPWR _20219_/X sky130_fd_sc_hd__mux4_1
X_28864_ _28864_/A VGND VGND VPWR VPWR _34745_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21199_ _21093_/X _21197_/X _21198_/X _21098_/X VGND VGND VPWR VPWR _21199_/X sky130_fd_sc_hd__a22o_1
XFILLER_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_829 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27815_ _27815_/A VGND VGND VPWR VPWR _34253_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28795_ _28795_/A VGND VGND VPWR VPWR _34712_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24958_ input47/X VGND VGND VPWR VPWR _24958_/X sky130_fd_sc_hd__buf_4
XFILLER_218_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27746_ _27745_/X _34231_/Q _27764_/S VGND VGND VPWR VPWR _27747_/A sky130_fd_sc_hd__mux2_1
XTAP_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23909_ _22980_/X _32500_/Q _23927_/S VGND VGND VPWR VPWR _23910_/A sky130_fd_sc_hd__mux2_1
XTAP_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24889_ input22/X VGND VGND VPWR VPWR _24889_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_45_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27677_ input3/X VGND VGND VPWR VPWR _27677_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_205_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29416_ input21/X VGND VGND VPWR VPWR _29416_/X sky130_fd_sc_hd__buf_2
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17430_ _35452_/Q _35388_/Q _35324_/Q _35260_/Q _17254_/X _17255_/X VGND VGND VPWR
+ VPWR _17430_/X sky130_fd_sc_hd__mux4_1
X_26628_ _31147_/B _31688_/B VGND VGND VPWR VPWR _26761_/S sky130_fd_sc_hd__nor2_8
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29347_ _29347_/A VGND VGND VPWR VPWR _34971_/D sky130_fd_sc_hd__clkbuf_1
X_17361_ _17355_/X _17360_/X _17151_/X VGND VGND VPWR VPWR _17371_/C sky130_fd_sc_hd__o21ba_1
X_26559_ _26559_/A VGND VGND VPWR VPWR _33718_/D sky130_fd_sc_hd__clkbuf_1
X_19100_ _19453_/A VGND VGND VPWR VPWR _19100_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_201_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16312_ _16312_/A _16312_/B _16312_/C _16312_/D VGND VGND VPWR VPWR _16313_/A sky130_fd_sc_hd__or4_4
X_17292_ _17998_/A VGND VGND VPWR VPWR _17292_/X sky130_fd_sc_hd__buf_6
X_29278_ _29326_/S VGND VGND VPWR VPWR _29297_/S sky130_fd_sc_hd__buf_4
XFILLER_198_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16243_ _16243_/A VGND VGND VPWR VPWR _31962_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_51_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19031_ _35176_/Q _35112_/Q _35048_/Q _32168_/Q _18957_/X _18958_/X VGND VGND VPWR
+ VPWR _19031_/X sky130_fd_sc_hd__mux4_1
X_28229_ _27816_/X _34446_/Q _28235_/S VGND VGND VPWR VPWR _28230_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_328_CLK clkbuf_6_39__f_CLK/X VGND VGND VPWR VPWR _32885_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_173_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31240_ _27776_/X _35841_/Q _31252_/S VGND VGND VPWR VPWR _31241_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16174_ _16091_/X _16172_/X _16173_/X _16101_/X VGND VGND VPWR VPWR _16174_/X sky130_fd_sc_hd__a22o_1
XFILLER_126_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput108 _31984_/Q VGND VGND VPWR VPWR D1[26] sky130_fd_sc_hd__buf_2
X_31171_ _27673_/X _35808_/Q _31189_/S VGND VGND VPWR VPWR _31172_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput119 _31994_/Q VGND VGND VPWR VPWR D1[36] sky130_fd_sc_hd__buf_2
XFILLER_217_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30122_ _30122_/A VGND VGND VPWR VPWR _35311_/D sky130_fd_sc_hd__clkbuf_1
X_19933_ _20286_/A VGND VGND VPWR VPWR _19933_/X sky130_fd_sc_hd__buf_4
XFILLER_99_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30053_ _35279_/Q _29506_/X _30057_/S VGND VGND VPWR VPWR _30054_/A sky130_fd_sc_hd__mux2_1
X_34930_ _35634_/CLK _34930_/D VGND VGND VPWR VPWR _34930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19864_ _19858_/X _19863_/X _19785_/X VGND VGND VPWR VPWR _19888_/A sky130_fd_sc_hd__o21ba_1
XFILLER_141_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_500_CLK clkbuf_6_2__f_CLK/X VGND VGND VPWR VPWR _36072_/CLK sky130_fd_sc_hd__clkbuf_16
Xclkbuf_6_2__f_CLK clkbuf_5_1_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_2__f_CLK/X sky130_fd_sc_hd__clkbuf_16
Xoutput90 _31958_/Q VGND VGND VPWR VPWR D1[0] sky130_fd_sc_hd__buf_2
XFILLER_228_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18815_ _18592_/X _18813_/X _18814_/X _18595_/X VGND VGND VPWR VPWR _18815_/X sky130_fd_sc_hd__a22o_1
XTAP_6080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34861_ _35566_/CLK _34861_/D VGND VGND VPWR VPWR _34861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19795_ _19789_/X _19792_/X _19793_/X _19794_/X VGND VGND VPWR VPWR _19820_/B sky130_fd_sc_hd__o211a_1
X_33812_ _33941_/CLK _33812_/D VGND VGND VPWR VPWR _33812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18746_ _18741_/X _18744_/X _18745_/X VGND VGND VPWR VPWR _18761_/C sky130_fd_sc_hd__o21ba_1
XFILLER_209_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34792_ _34920_/CLK _34792_/D VGND VGND VPWR VPWR _34792_/Q sky130_fd_sc_hd__dfxtp_1
X_33743_ _35661_/CLK _33743_/D VGND VGND VPWR VPWR _33743_/Q sky130_fd_sc_hd__dfxtp_1
X_18677_ _34654_/Q _34590_/Q _34526_/Q _34462_/Q _18533_/X _18534_/X VGND VGND VPWR
+ VPWR _18677_/X sky130_fd_sc_hd__mux4_1
X_30955_ _30955_/A VGND VGND VPWR VPWR _35706_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_1214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17628_ _17624_/X _17627_/X _17485_/X VGND VGND VPWR VPWR _17654_/A sky130_fd_sc_hd__o21ba_1
X_33674_ _33869_/CLK _33674_/D VGND VGND VPWR VPWR _33674_/Q sky130_fd_sc_hd__dfxtp_1
X_30886_ _30886_/A VGND VGND VPWR VPWR _35673_/D sky130_fd_sc_hd__clkbuf_1
X_35413_ _36055_/CLK _35413_/D VGND VGND VPWR VPWR _35413_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32625_ _36017_/CLK _32625_/D VGND VGND VPWR VPWR _32625_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17559_ _17912_/A VGND VGND VPWR VPWR _17559_/X sky130_fd_sc_hd__buf_4
XFILLER_177_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35344_ _35729_/CLK _35344_/D VGND VGND VPWR VPWR _35344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20570_ _34709_/Q _34645_/Q _34581_/Q _34517_/Q _20298_/X _20299_/X VGND VGND VPWR
+ VPWR _20570_/X sky130_fd_sc_hd__mux4_1
X_32556_ _35949_/CLK _32556_/D VGND VGND VPWR VPWR _32556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31507_ _31507_/A VGND VGND VPWR VPWR _35967_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19229_ _32878_/Q _32814_/Q _32750_/Q _32686_/Q _18940_/X _18941_/X VGND VGND VPWR
+ VPWR _19229_/X sky130_fd_sc_hd__mux4_1
X_35275_ _35596_/CLK _35275_/D VGND VGND VPWR VPWR _35275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_319_CLK clkbuf_6_37__f_CLK/X VGND VGND VPWR VPWR _32906_/CLK sky130_fd_sc_hd__clkbuf_16
X_32487_ _35944_/CLK _32487_/D VGND VGND VPWR VPWR _32487_/Q sky130_fd_sc_hd__dfxtp_1
X_22240_ _21951_/X _22238_/X _22239_/X _21954_/X VGND VGND VPWR VPWR _22240_/X sky130_fd_sc_hd__a22o_1
X_34226_ _34611_/CLK _34226_/D VGND VGND VPWR VPWR _34226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31438_ _27670_/X _35935_/Q _31438_/S VGND VGND VPWR VPWR _31439_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_1015 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22171_ _22167_/X _22170_/X _22093_/X _22094_/X VGND VGND VPWR VPWR _22188_/B sky130_fd_sc_hd__o211a_1
XFILLER_117_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34157_ _35630_/CLK _34157_/D VGND VGND VPWR VPWR _34157_/Q sky130_fd_sc_hd__dfxtp_1
X_31369_ _27766_/X _35902_/Q _31387_/S VGND VGND VPWR VPWR _31370_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_1368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33108_ _35858_/CLK _33108_/D VGND VGND VPWR VPWR _33108_/Q sky130_fd_sc_hd__dfxtp_1
X_21122_ _21047_/X _21120_/X _21121_/X _21050_/X VGND VGND VPWR VPWR _21122_/X sky130_fd_sc_hd__a22o_1
XFILLER_105_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34088_ _34920_/CLK _34088_/D VGND VGND VPWR VPWR _34088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25930_ _25930_/A VGND VGND VPWR VPWR _33421_/D sky130_fd_sc_hd__clkbuf_1
X_33039_ _36045_/CLK _33039_/D VGND VGND VPWR VPWR _33039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21053_ _34400_/Q _36128_/Q _34272_/Q _34208_/Q _20770_/X _20771_/X VGND VGND VPWR
+ VPWR _21053_/X sky130_fd_sc_hd__mux4_1
XFILLER_59_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20004_ _20159_/A VGND VGND VPWR VPWR _20004_/X sky130_fd_sc_hd__clkbuf_4
X_25861_ _25861_/A VGND VGND VPWR VPWR _33388_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_247_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27600_ _34179_/Q _27174_/X _27608_/S VGND VGND VPWR VPWR _27601_/A sky130_fd_sc_hd__mux2_1
X_24812_ input45/X VGND VGND VPWR VPWR _24812_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_46_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25792_ _24967_/X _33356_/Q _25802_/S VGND VGND VPWR VPWR _25793_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28580_ _27735_/X _34612_/Q _28598_/S VGND VGND VPWR VPWR _28581_/A sky130_fd_sc_hd__mux2_1
XFILLER_234_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27531_ _34146_/Q _27072_/X _27545_/S VGND VGND VPWR VPWR _27532_/A sky130_fd_sc_hd__mux2_1
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24743_ _24743_/A VGND VGND VPWR VPWR _32892_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21955_ _21951_/X _21952_/X _21953_/X _21954_/X VGND VGND VPWR VPWR _21955_/X sky130_fd_sc_hd__a22o_1
XFILLER_28_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27462_ _27462_/A VGND VGND VPWR VPWR _34113_/D sky130_fd_sc_hd__clkbuf_1
X_20906_ _35164_/Q _35100_/Q _35036_/Q _32156_/Q _20904_/X _20905_/X VGND VGND VPWR
+ VPWR _20906_/X sky130_fd_sc_hd__mux4_1
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24674_ _24674_/A VGND VGND VPWR VPWR _32859_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21886_ _35640_/Q _35000_/Q _34360_/Q _33720_/Q _21744_/X _21745_/X VGND VGND VPWR
+ VPWR _21886_/X sky130_fd_sc_hd__mux4_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29201_ _34905_/Q _27044_/X _29213_/S VGND VGND VPWR VPWR _29202_/A sky130_fd_sc_hd__mux2_1
XFILLER_203_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26413_ _33650_/Q _23381_/X _26415_/S VGND VGND VPWR VPWR _26414_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23625_ _22968_/X _32304_/Q _23631_/S VGND VGND VPWR VPWR _23626_/A sky130_fd_sc_hd__mux2_1
X_20837_ _20678_/X _20835_/X _20836_/X _20688_/X VGND VGND VPWR VPWR _20837_/X sky130_fd_sc_hd__a22o_1
XFILLER_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27393_ _27393_/A VGND VGND VPWR VPWR _34080_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26344_ _24985_/X _33618_/Q _26350_/S VGND VGND VPWR VPWR _26345_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29132_ _29132_/A VGND VGND VPWR VPWR _34872_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23556_ _23556_/A VGND VGND VPWR VPWR _32272_/D sky130_fd_sc_hd__clkbuf_1
X_20768_ _35160_/Q _35096_/Q _35032_/Q _32152_/Q _20683_/X _20685_/X VGND VGND VPWR
+ VPWR _20768_/X sky130_fd_sc_hd__mux4_1
XFILLER_195_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1006 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29063_ _29063_/A VGND VGND VPWR VPWR _34839_/D sky130_fd_sc_hd__clkbuf_1
X_22507_ _22507_/A VGND VGND VPWR VPWR _22507_/X sky130_fd_sc_hd__buf_4
X_26275_ _24883_/X _33585_/Q _26279_/S VGND VGND VPWR VPWR _26276_/A sky130_fd_sc_hd__mux2_1
X_23487_ input57/X VGND VGND VPWR VPWR _23487_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_167_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20699_ _34902_/Q _34838_/Q _34774_/Q _34710_/Q _20696_/X _20698_/X VGND VGND VPWR
+ VPWR _20699_/X sky130_fd_sc_hd__mux4_1
X_25226_ _33089_/Q _23432_/X _25238_/S VGND VGND VPWR VPWR _25227_/A sky130_fd_sc_hd__mux2_1
X_28014_ _34344_/Q _27090_/X _28016_/S VGND VGND VPWR VPWR _28015_/A sky130_fd_sc_hd__mux2_1
X_22438_ _22438_/A VGND VGND VPWR VPWR _22438_/X sky130_fd_sc_hd__buf_2
XFILLER_13_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25157_ _33056_/Q _23261_/X _25175_/S VGND VGND VPWR VPWR _25158_/A sky130_fd_sc_hd__mux2_1
X_22369_ _22374_/A VGND VGND VPWR VPWR _22369_/X sky130_fd_sc_hd__clkbuf_4
X_24108_ _24108_/A VGND VGND VPWR VPWR _32594_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25088_ _25088_/A VGND VGND VPWR VPWR _33024_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29965_ _35237_/Q _29376_/X _29973_/S VGND VGND VPWR VPWR _29966_/A sky130_fd_sc_hd__mux2_1
X_28916_ _28916_/A VGND VGND VPWR VPWR _34770_/D sky130_fd_sc_hd__clkbuf_1
X_24039_ _24039_/A VGND VGND VPWR VPWR _32561_/D sky130_fd_sc_hd__clkbuf_1
X_16930_ _16714_/X _16928_/X _16929_/X _16718_/X VGND VGND VPWR VPWR _16930_/X sky130_fd_sc_hd__a22o_1
XFILLER_215_1435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29896_ _29896_/A VGND VGND VPWR VPWR _35204_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_1271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28847_ _28847_/A VGND VGND VPWR VPWR _34737_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16861_ _16706_/X _16859_/X _16860_/X _16712_/X VGND VGND VPWR VPWR _16861_/X sky130_fd_sc_hd__a22o_1
XFILLER_77_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18600_ _20169_/A VGND VGND VPWR VPWR _18600_/X sky130_fd_sc_hd__buf_4
XFILLER_24_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_912 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19580_ _20286_/A VGND VGND VPWR VPWR _19580_/X sky130_fd_sc_hd__clkbuf_8
X_28778_ _34706_/Q _27220_/X _28784_/S VGND VGND VPWR VPWR _28779_/A sky130_fd_sc_hd__mux2_1
X_16792_ _17999_/A VGND VGND VPWR VPWR _16792_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_237_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18531_ _18360_/X _18529_/X _18530_/X _18372_/X VGND VGND VPWR VPWR _18531_/X sky130_fd_sc_hd__a22o_1
XFILLER_18_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27729_ input21/X VGND VGND VPWR VPWR _27729_/X sky130_fd_sc_hd__buf_2
XTAP_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18462_ _18348_/X _18460_/X _18461_/X _18358_/X VGND VGND VPWR VPWR _18462_/X sky130_fd_sc_hd__a22o_1
X_30740_ _35605_/Q _29524_/X _30740_/S VGND VGND VPWR VPWR _30741_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17413_ _17766_/A VGND VGND VPWR VPWR _17413_/X sky130_fd_sc_hd__buf_4
XFILLER_60_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18393_ _20066_/A VGND VGND VPWR VPWR _19177_/A sky130_fd_sc_hd__buf_8
X_30671_ _30740_/S VGND VGND VPWR VPWR _30690_/S sky130_fd_sc_hd__buf_6
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32410_ _34151_/CLK _32410_/D VGND VGND VPWR VPWR _32410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17344_ _17059_/X _17342_/X _17343_/X _17065_/X VGND VGND VPWR VPWR _17344_/X sky130_fd_sc_hd__a22o_1
XFILLER_144_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33390_ _36079_/CLK _33390_/D VGND VGND VPWR VPWR _33390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32341_ _35922_/CLK _32341_/D VGND VGND VPWR VPWR _32341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17275_ _17271_/X _17274_/X _17132_/X VGND VGND VPWR VPWR _17301_/A sky130_fd_sc_hd__o21ba_1
XFILLER_158_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19014_ _20212_/A VGND VGND VPWR VPWR _19014_/X sky130_fd_sc_hd__clkbuf_4
X_16226_ _35674_/Q _32180_/Q _35546_/Q _35482_/Q _16049_/X _16050_/X VGND VGND VPWR
+ VPWR _16226_/X sky130_fd_sc_hd__mux4_1
X_35060_ _35124_/CLK _35060_/D VGND VGND VPWR VPWR _35060_/Q sky130_fd_sc_hd__dfxtp_1
X_32272_ _36115_/CLK _32272_/D VGND VGND VPWR VPWR _32272_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34011_ _36212_/CLK _34011_/D VGND VGND VPWR VPWR _34011_/Q sky130_fd_sc_hd__dfxtp_1
X_16157_ _32856_/Q _32792_/Q _32728_/Q _32664_/Q _16037_/X _16039_/X VGND VGND VPWR
+ VPWR _16157_/X sky130_fd_sc_hd__mux4_1
X_31223_ _27751_/X _35833_/Q _31231_/S VGND VGND VPWR VPWR _31224_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31154_ _27649_/X _35800_/Q _31168_/S VGND VGND VPWR VPWR _31155_/A sky130_fd_sc_hd__mux2_1
X_16088_ _17156_/A VGND VGND VPWR VPWR _16088_/X sky130_fd_sc_hd__buf_4
XFILLER_103_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19916_ _34433_/Q _36161_/Q _34305_/Q _34241_/Q _19882_/X _19883_/X VGND VGND VPWR
+ VPWR _19916_/X sky130_fd_sc_hd__mux4_1
X_30105_ _30105_/A VGND VGND VPWR VPWR _35303_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31085_ _35768_/Q input28/X _31095_/S VGND VGND VPWR VPWR _31086_/A sky130_fd_sc_hd__mux2_1
X_35962_ _35962_/CLK _35962_/D VGND VGND VPWR VPWR _35962_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30036_ _35271_/Q _29481_/X _30036_/S VGND VGND VPWR VPWR _30037_/A sky130_fd_sc_hd__mux2_1
X_34913_ _34913_/CLK _34913_/D VGND VGND VPWR VPWR _34913_/Q sky130_fd_sc_hd__dfxtp_1
X_19847_ _34943_/Q _34879_/Q _34815_/Q _34751_/Q _19813_/X _19814_/X VGND VGND VPWR
+ VPWR _19847_/X sky130_fd_sc_hd__mux4_1
X_35893_ _35956_/CLK _35893_/D VGND VGND VPWR VPWR _35893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34844_ _36242_/CLK _34844_/D VGND VGND VPWR VPWR _34844_/Q sky130_fd_sc_hd__dfxtp_1
X_19778_ _34174_/Q _34110_/Q _34046_/Q _33982_/Q _19746_/X _19747_/X VGND VGND VPWR
+ VPWR _19778_/X sky130_fd_sc_hd__mux4_1
XFILLER_216_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18729_ _33120_/Q _36000_/Q _32992_/Q _32928_/Q _18656_/X _18657_/X VGND VGND VPWR
+ VPWR _18729_/X sky130_fd_sc_hd__mux4_1
X_34775_ _34904_/CLK _34775_/D VGND VGND VPWR VPWR _34775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31987_ _34914_/CLK _31987_/D VGND VGND VPWR VPWR _31987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33726_ _35646_/CLK _33726_/D VGND VGND VPWR VPWR _33726_/Q sky130_fd_sc_hd__dfxtp_1
X_21740_ _22446_/A VGND VGND VPWR VPWR _21740_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_97_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30938_ _30938_/A VGND VGND VPWR VPWR _35698_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_240_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33657_ _33913_/CLK _33657_/D VGND VGND VPWR VPWR _33657_/Q sky130_fd_sc_hd__dfxtp_1
X_21671_ _22515_/A VGND VGND VPWR VPWR _21671_/X sky130_fd_sc_hd__clkbuf_4
X_30869_ _35666_/Q input57/X _30875_/S VGND VGND VPWR VPWR _30870_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_96_CLK clkbuf_leaf_96_CLK/A VGND VGND VPWR VPWR _36060_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_184_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23410_ _23410_/A VGND VGND VPWR VPWR _32215_/D sky130_fd_sc_hd__clkbuf_1
X_20622_ _22366_/A VGND VGND VPWR VPWR _22317_/A sky130_fd_sc_hd__buf_8
XFILLER_127_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32608_ _36002_/CLK _32608_/D VGND VGND VPWR VPWR _32608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24390_ _24390_/A VGND VGND VPWR VPWR _32725_/D sky130_fd_sc_hd__clkbuf_1
X_33588_ _35699_/CLK _33588_/D VGND VGND VPWR VPWR _33588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35327_ _35839_/CLK _35327_/D VGND VGND VPWR VPWR _35327_/Q sky130_fd_sc_hd__dfxtp_1
X_23341_ _32187_/Q _23340_/X _23424_/S VGND VGND VPWR VPWR _23342_/A sky130_fd_sc_hd__mux2_1
X_20553_ _33941_/Q _33877_/Q _33813_/Q _36117_/Q _18362_/X _18364_/X VGND VGND VPWR
+ VPWR _20553_/X sky130_fd_sc_hd__mux4_1
X_32539_ _35995_/CLK _32539_/D VGND VGND VPWR VPWR _32539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26060_ _24964_/X _33483_/Q _26072_/S VGND VGND VPWR VPWR _26061_/A sky130_fd_sc_hd__mux2_1
X_23272_ _32163_/Q _23271_/X _23290_/S VGND VGND VPWR VPWR _23273_/A sky130_fd_sc_hd__mux2_1
X_35258_ _36026_/CLK _35258_/D VGND VGND VPWR VPWR _35258_/Q sky130_fd_sc_hd__dfxtp_1
X_20484_ _34962_/Q _34898_/Q _34834_/Q _34770_/Q _18383_/X _18385_/X VGND VGND VPWR
+ VPWR _20484_/X sky130_fd_sc_hd__mux4_1
XFILLER_165_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25011_ _24818_/X _32988_/Q _25017_/S VGND VGND VPWR VPWR _25012_/A sky130_fd_sc_hd__mux2_1
X_22223_ _34178_/Q _34114_/Q _34050_/Q _33986_/Q _22046_/X _22047_/X VGND VGND VPWR
+ VPWR _22223_/X sky130_fd_sc_hd__mux4_1
X_34209_ _36128_/CLK _34209_/D VGND VGND VPWR VPWR _34209_/Q sky130_fd_sc_hd__dfxtp_1
X_35189_ _35829_/CLK _35189_/D VGND VGND VPWR VPWR _35189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22154_ _22507_/A VGND VGND VPWR VPWR _22154_/X sky130_fd_sc_hd__buf_4
XFILLER_79_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21105_ _21099_/X _21104_/X _21026_/X VGND VGND VPWR VPWR _21129_/A sky130_fd_sc_hd__o21ba_1
X_29750_ _35135_/Q _29457_/X _29766_/S VGND VGND VPWR VPWR _29751_/A sky130_fd_sc_hd__mux2_1
XTAP_6838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22085_ _22438_/A VGND VGND VPWR VPWR _22085_/X sky130_fd_sc_hd__clkbuf_4
X_26962_ _27031_/S VGND VGND VPWR VPWR _26981_/S sky130_fd_sc_hd__buf_4
XFILLER_102_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_20_CLK clkbuf_6_4__f_CLK/X VGND VGND VPWR VPWR _35554_/CLK sky130_fd_sc_hd__clkbuf_16
X_28701_ _34669_/Q _27106_/X _28713_/S VGND VGND VPWR VPWR _28702_/A sky130_fd_sc_hd__mux2_1
X_25913_ _25913_/A VGND VGND VPWR VPWR _33413_/D sky130_fd_sc_hd__clkbuf_1
X_21036_ _21030_/X _21033_/X _21034_/X _21035_/X VGND VGND VPWR VPWR _21061_/B sky130_fd_sc_hd__o211a_1
XFILLER_43_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29681_ _29681_/A VGND VGND VPWR VPWR _35102_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_1056 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26893_ _26893_/A VGND VGND VPWR VPWR _33875_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28632_ _27813_/X _34637_/Q _28640_/S VGND VGND VPWR VPWR _28633_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25844_ _25844_/A VGND VGND VPWR VPWR _33380_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_1051 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28563_ _27711_/X _34604_/Q _28577_/S VGND VGND VPWR VPWR _28564_/A sky130_fd_sc_hd__mux2_1
X_25775_ _24942_/X _33348_/Q _25781_/S VGND VGND VPWR VPWR _25776_/A sky130_fd_sc_hd__mux2_1
X_22987_ input26/X VGND VGND VPWR VPWR _22987_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_55_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27514_ _34138_/Q _27047_/X _27524_/S VGND VGND VPWR VPWR _27515_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21938_ _33402_/Q _33338_/Q _33274_/Q _33210_/Q _21727_/X _21728_/X VGND VGND VPWR
+ VPWR _21938_/X sky130_fd_sc_hd__mux4_1
X_24726_ _22980_/X _32884_/Q _24744_/S VGND VGND VPWR VPWR _24727_/A sky130_fd_sc_hd__mux2_1
XFILLER_245_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28494_ _28494_/A VGND VGND VPWR VPWR _34571_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_243_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24657_ _23079_/X _32852_/Q _24659_/S VGND VGND VPWR VPWR _24658_/A sky130_fd_sc_hd__mux2_1
X_27445_ _27445_/A VGND VGND VPWR VPWR _34105_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21869_ _33656_/Q _33592_/Q _33528_/Q _33464_/Q _21800_/X _21801_/X VGND VGND VPWR
+ VPWR _21869_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_87_CLK clkbuf_leaf_88_CLK/A VGND VGND VPWR VPWR _35743_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_128_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23608_ _22943_/X _32296_/Q _23610_/S VGND VGND VPWR VPWR _23609_/A sky130_fd_sc_hd__mux2_1
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27376_ _27376_/A VGND VGND VPWR VPWR _34072_/D sky130_fd_sc_hd__clkbuf_1
X_24588_ _22977_/X _32819_/Q _24588_/S VGND VGND VPWR VPWR _24589_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29115_ _29115_/A VGND VGND VPWR VPWR _34864_/D sky130_fd_sc_hd__clkbuf_1
X_26327_ _26327_/A VGND VGND VPWR VPWR _33609_/D sky130_fd_sc_hd__clkbuf_1
X_23539_ _32264_/Q _23453_/X _23557_/S VGND VGND VPWR VPWR _23540_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17060_ _17766_/A VGND VGND VPWR VPWR _17060_/X sky130_fd_sc_hd__clkbuf_4
X_29046_ _34832_/Q _27214_/X _29048_/S VGND VGND VPWR VPWR _29047_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26258_ _24858_/X _33577_/Q _26258_/S VGND VGND VPWR VPWR _26259_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16011_ _17961_/A VGND VGND VPWR VPWR _16011_/X sky130_fd_sc_hd__buf_4
XFILLER_155_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25209_ _33081_/Q _23405_/X _25217_/S VGND VGND VPWR VPWR _25210_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26189_ _24954_/X _33544_/Q _26207_/S VGND VGND VPWR VPWR _26190_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_907 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_6_15__f_CLK clkbuf_5_7_0_CLK/X VGND VGND VPWR VPWR clkbuf_leaf_61_CLK/A sky130_fd_sc_hd__clkbuf_16
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17962_ _35467_/Q _35403_/Q _35339_/Q _35275_/Q _17960_/X _17961_/X VGND VGND VPWR
+ VPWR _17962_/X sky130_fd_sc_hd__mux4_1
X_29948_ _35229_/Q _29351_/X _29952_/S VGND VGND VPWR VPWR _29949_/A sky130_fd_sc_hd__mux2_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_11_CLK clkbuf_6_3__f_CLK/X VGND VGND VPWR VPWR _35177_/CLK sky130_fd_sc_hd__clkbuf_16
X_19701_ _19458_/X _19699_/X _19700_/X _19463_/X VGND VGND VPWR VPWR _19701_/X sky130_fd_sc_hd__a22o_1
X_16913_ _16909_/X _16912_/X _16812_/X VGND VGND VPWR VPWR _16914_/D sky130_fd_sc_hd__o21ba_1
XFILLER_78_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17893_ _33097_/Q _32073_/Q _35849_/Q _35785_/Q _17784_/X _17785_/X VGND VGND VPWR
+ VPWR _17893_/X sky130_fd_sc_hd__mux4_1
XFILLER_61_1438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29879_ _29879_/A VGND VGND VPWR VPWR _35196_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_215_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31910_ _31910_/A VGND VGND VPWR VPWR _36158_/D sky130_fd_sc_hd__clkbuf_1
X_19632_ _19628_/X _19631_/X _19465_/X VGND VGND VPWR VPWR _19633_/D sky130_fd_sc_hd__o21ba_1
XFILLER_226_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16844_ _16844_/A _16844_/B _16844_/C _16844_/D VGND VGND VPWR VPWR _16845_/A sky130_fd_sc_hd__or4_4
XFILLER_65_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32890_ _32890_/CLK _32890_/D VGND VGND VPWR VPWR _32890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31841_ _23255_/X _36126_/Q _31843_/S VGND VGND VPWR VPWR _31842_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_1290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19563_ _34423_/Q _36151_/Q _34295_/Q _34231_/Q _19529_/X _19530_/X VGND VGND VPWR
+ VPWR _19563_/X sky130_fd_sc_hd__mux4_1
XFILLER_81_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16775_ _17834_/A VGND VGND VPWR VPWR _16775_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_111_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18514_ _33882_/Q _33818_/Q _33754_/Q _36058_/Q _18412_/X _18413_/X VGND VGND VPWR
+ VPWR _18514_/X sky130_fd_sc_hd__mux4_1
XFILLER_248_1052 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34560_ _34690_/CLK _34560_/D VGND VGND VPWR VPWR _34560_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31772_ _31772_/A VGND VGND VPWR VPWR _36093_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19494_ _34933_/Q _34869_/Q _34805_/Q _34741_/Q _19460_/X _19461_/X VGND VGND VPWR
+ VPWR _19494_/X sky130_fd_sc_hd__mux4_1
XFILLER_59_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33511_ _36068_/CLK _33511_/D VGND VGND VPWR VPWR _33511_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30723_ _30723_/A VGND VGND VPWR VPWR _35596_/D sky130_fd_sc_hd__clkbuf_1
X_18445_ _20162_/A VGND VGND VPWR VPWR _18445_/X sky130_fd_sc_hd__buf_4
XFILLER_22_907 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34491_ _34685_/CLK _34491_/D VGND VGND VPWR VPWR _34491_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_78_CLK clkbuf_leaf_81_CLK/A VGND VGND VPWR VPWR _35994_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_36230_ _36235_/CLK _36230_/D VGND VGND VPWR VPWR _36230_/Q sky130_fd_sc_hd__dfxtp_1
X_33442_ _33573_/CLK _33442_/D VGND VGND VPWR VPWR _33442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18376_ _18359_/X _18373_/X _18375_/X VGND VGND VPWR VPWR _18406_/C sky130_fd_sc_hd__o21ba_1
XFILLER_159_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30654_ _30654_/A VGND VGND VPWR VPWR _35563_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_222_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_36161_ _36161_/CLK _36161_/D VGND VGND VPWR VPWR _36161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17327_ _35193_/Q _35129_/Q _35065_/Q _32249_/Q _17010_/X _17011_/X VGND VGND VPWR
+ VPWR _17327_/X sky130_fd_sc_hd__mux4_1
X_33373_ _33821_/CLK _33373_/D VGND VGND VPWR VPWR _33373_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30585_ _35531_/Q _29494_/X _30597_/S VGND VGND VPWR VPWR _30586_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35112_ _35176_/CLK _35112_/D VGND VGND VPWR VPWR _35112_/Q sky130_fd_sc_hd__dfxtp_1
X_32324_ _35973_/CLK _32324_/D VGND VGND VPWR VPWR _32324_/Q sky130_fd_sc_hd__dfxtp_1
X_36092_ _36092_/CLK _36092_/D VGND VGND VPWR VPWR _36092_/Q sky130_fd_sc_hd__dfxtp_1
X_17258_ _17003_/X _17256_/X _17257_/X _17006_/X VGND VGND VPWR VPWR _17258_/X sky130_fd_sc_hd__a22o_1
XFILLER_31_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16209_ _16209_/A VGND VGND VPWR VPWR _31961_/D sky130_fd_sc_hd__clkbuf_4
X_35043_ _36210_/CLK _35043_/D VGND VGND VPWR VPWR _35043_/Q sky130_fd_sc_hd__dfxtp_1
X_32255_ _36100_/CLK _32255_/D VGND VGND VPWR VPWR _32255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17189_ _17185_/X _17188_/X _17151_/X VGND VGND VPWR VPWR _17197_/C sky130_fd_sc_hd__o21ba_1
XFILLER_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31206_ _27726_/X _35825_/Q _31210_/S VGND VGND VPWR VPWR _31207_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32186_ _35747_/CLK _32186_/D VGND VGND VPWR VPWR _32186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31137_ _35793_/Q input55/X _31137_/S VGND VGND VPWR VPWR _31138_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31068_ _35760_/Q input19/X _31074_/S VGND VGND VPWR VPWR _31069_/A sky130_fd_sc_hd__mux2_1
X_35945_ _35945_/CLK _35945_/D VGND VGND VPWR VPWR _35945_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_1276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22910_ _22909_/X _32029_/Q _22916_/S VGND VGND VPWR VPWR _22911_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30019_ _30019_/A VGND VGND VPWR VPWR _35262_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23890_ _22953_/X _32491_/Q _23906_/S VGND VGND VPWR VPWR _23891_/A sky130_fd_sc_hd__mux2_1
X_35876_ _35939_/CLK _35876_/D VGND VGND VPWR VPWR _35876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34827_ _34957_/CLK _34827_/D VGND VGND VPWR VPWR _34827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22841_ _35220_/Q _35156_/Q _35092_/Q _32276_/Q _20692_/X _20694_/X VGND VGND VPWR
+ VPWR _22841_/X sky130_fd_sc_hd__mux4_1
XFILLER_216_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25560_ _24824_/X _33246_/Q _25562_/S VGND VGND VPWR VPWR _25561_/A sky130_fd_sc_hd__mux2_1
X_34758_ _36167_/CLK _34758_/D VGND VGND VPWR VPWR _34758_/Q sky130_fd_sc_hd__dfxtp_1
X_22772_ _22768_/X _22771_/X _22446_/A _22447_/A VGND VGND VPWR VPWR _22787_/B sky130_fd_sc_hd__o211a_1
XFILLER_231_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24511_ _24511_/A VGND VGND VPWR VPWR _32782_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_212_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21723_ _21723_/A VGND VGND VPWR VPWR _36211_/D sky130_fd_sc_hd__clkbuf_4
X_33709_ _35693_/CLK _33709_/D VGND VGND VPWR VPWR _33709_/Q sky130_fd_sc_hd__dfxtp_1
X_25491_ _25491_/A VGND VGND VPWR VPWR _33213_/D sky130_fd_sc_hd__clkbuf_1
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34689_ _34690_/CLK _34689_/D VGND VGND VPWR VPWR _34689_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_69_CLK clkbuf_leaf_73_CLK/A VGND VGND VPWR VPWR _32802_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27230_ _34005_/Q _27229_/X _27230_/S VGND VGND VPWR VPWR _27231_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24442_ _24442_/A VGND VGND VPWR VPWR _32749_/D sky130_fd_sc_hd__clkbuf_1
X_21654_ _21446_/X _21652_/X _21653_/X _21451_/X VGND VGND VPWR VPWR _21654_/X sky130_fd_sc_hd__a22o_1
X_20605_ input74/X input73/X VGND VGND VPWR VPWR _22377_/A sky130_fd_sc_hd__nor2b_4
X_27161_ _27161_/A VGND VGND VPWR VPWR _33982_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24373_ _23058_/X _32717_/Q _24381_/S VGND VGND VPWR VPWR _24374_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21585_ _33392_/Q _33328_/Q _33264_/Q _33200_/Q _21374_/X _21375_/X VGND VGND VPWR
+ VPWR _21585_/X sky130_fd_sc_hd__mux4_1
XFILLER_137_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26112_ _26112_/A VGND VGND VPWR VPWR _33507_/D sky130_fd_sc_hd__clkbuf_1
X_23324_ _23324_/A VGND VGND VPWR VPWR _32179_/D sky130_fd_sc_hd__clkbuf_1
X_20536_ _35476_/Q _35412_/Q _35348_/Q _35284_/Q _20260_/X _20261_/X VGND VGND VPWR
+ VPWR _20536_/X sky130_fd_sc_hd__mux4_1
X_27092_ _27092_/A VGND VGND VPWR VPWR _33960_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26043_ _24939_/X _33475_/Q _26051_/S VGND VGND VPWR VPWR _26044_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23255_ input63/X VGND VGND VPWR VPWR _23255_/X sky130_fd_sc_hd__buf_4
XFILLER_4_616 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20467_ _33170_/Q _36050_/Q _33042_/Q _32978_/Q _18332_/X _19461_/A VGND VGND VPWR
+ VPWR _20467_/X sky130_fd_sc_hd__mux4_1
XFILLER_119_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_238_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22206_ _21951_/X _22204_/X _22205_/X _21954_/X VGND VGND VPWR VPWR _22206_/X sky130_fd_sc_hd__a22o_1
XFILLER_106_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23186_ _23027_/X _32131_/Q _23194_/S VGND VGND VPWR VPWR _23187_/A sky130_fd_sc_hd__mux2_1
X_20398_ _20398_/A VGND VGND VPWR VPWR _32463_/D sky130_fd_sc_hd__clkbuf_4
Xclkbuf_5_3_0_CLK clkbuf_5_7_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_3_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XTAP_6602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29802_ _29802_/A VGND VGND VPWR VPWR _35159_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22137_ _35647_/Q _35007_/Q _34367_/Q _33727_/Q _22097_/X _22098_/X VGND VGND VPWR
+ VPWR _22137_/X sky130_fd_sc_hd__mux4_1
XFILLER_134_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27994_ _27994_/A VGND VGND VPWR VPWR _34334_/D sky130_fd_sc_hd__clkbuf_1
Xoutput280 _32414_/Q VGND VGND VPWR VPWR D3[8] sky130_fd_sc_hd__buf_2
XTAP_6646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29733_ _35127_/Q _29432_/X _29745_/S VGND VGND VPWR VPWR _29734_/A sky130_fd_sc_hd__mux2_1
XTAP_6668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26945_ _26945_/A VGND VGND VPWR VPWR _33899_/D sky130_fd_sc_hd__clkbuf_1
X_22068_ _34685_/Q _34621_/Q _34557_/Q _34493_/Q _21892_/X _21893_/X VGND VGND VPWR
+ VPWR _22068_/X sky130_fd_sc_hd__mux4_1
XTAP_6679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21019_ _34144_/Q _34080_/Q _34016_/Q _33952_/Q _20987_/X _20988_/X VGND VGND VPWR
+ VPWR _21019_/X sky130_fd_sc_hd__mux4_1
X_29664_ _35094_/Q _29328_/X _29682_/S VGND VGND VPWR VPWR _29665_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26876_ _33867_/Q _23466_/X _26888_/S VGND VGND VPWR VPWR _26877_/A sky130_fd_sc_hd__mux2_1
XTAP_5978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28615_ _27788_/X _34629_/Q _28619_/S VGND VGND VPWR VPWR _28616_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25827_ _25827_/A VGND VGND VPWR VPWR _33372_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29595_ _29595_/A VGND VGND VPWR VPWR _35061_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28546_ _27686_/X _34596_/Q _28556_/S VGND VGND VPWR VPWR _28547_/A sky130_fd_sc_hd__mux2_1
X_16560_ _16556_/X _16559_/X _16459_/X VGND VGND VPWR VPWR _16561_/D sky130_fd_sc_hd__o21ba_1
XFILLER_210_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25758_ _24917_/X _33340_/Q _25760_/S VGND VGND VPWR VPWR _25759_/A sky130_fd_sc_hd__mux2_1
XFILLER_245_1214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24709_ _22956_/X _32876_/Q _24723_/S VGND VGND VPWR VPWR _24710_/A sky130_fd_sc_hd__mux2_1
X_28477_ _28477_/A VGND VGND VPWR VPWR _34563_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16491_ _16491_/A _16491_/B _16491_/C _16491_/D VGND VGND VPWR VPWR _16492_/A sky130_fd_sc_hd__or4_4
X_25689_ _24815_/X _33307_/Q _25697_/S VGND VGND VPWR VPWR _25690_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_245_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18230_ _32916_/Q _32852_/Q _32788_/Q _32724_/Q _15984_/X _15987_/X VGND VGND VPWR
+ VPWR _18230_/X sky130_fd_sc_hd__mux4_1
XFILLER_54_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27428_ _27428_/A VGND VGND VPWR VPWR _34097_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_0_CLK clkbuf_leaf_2_CLK/A VGND VGND VPWR VPWR _34085_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_19_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18161_ _17905_/X _18159_/X _18160_/X _17910_/X VGND VGND VPWR VPWR _18161_/X sky130_fd_sc_hd__a22o_1
XFILLER_169_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27359_ _34065_/Q _27217_/X _27359_/S VGND VGND VPWR VPWR _27360_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17112_ _33075_/Q _32051_/Q _35827_/Q _35763_/Q _17078_/X _17079_/X VGND VGND VPWR
+ VPWR _17112_/X sky130_fd_sc_hd__mux4_1
X_18092_ _17859_/X _18090_/X _18091_/X _17862_/X VGND VGND VPWR VPWR _18092_/X sky130_fd_sc_hd__a22o_1
X_30370_ _35429_/Q _29376_/X _30378_/S VGND VGND VPWR VPWR _30371_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29029_ _29056_/S VGND VGND VPWR VPWR _29048_/S sky130_fd_sc_hd__buf_4
XFILLER_184_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17043_ _34673_/Q _34609_/Q _34545_/Q _34481_/Q _16939_/X _16940_/X VGND VGND VPWR
+ VPWR _17043_/X sky130_fd_sc_hd__mux4_1
XFILLER_171_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32040_ _35753_/CLK _32040_/D VGND VGND VPWR VPWR _32040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18994_ _34919_/Q _34855_/Q _34791_/Q _34727_/Q _18754_/X _18755_/X VGND VGND VPWR
+ VPWR _18994_/X sky130_fd_sc_hd__mux4_1
XFILLER_225_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17945_ _17905_/X _17943_/X _17944_/X _17910_/X VGND VGND VPWR VPWR _17945_/X sky130_fd_sc_hd__a22o_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33991_ _34185_/CLK _33991_/D VGND VGND VPWR VPWR _33991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35730_ _35730_/CLK _35730_/D VGND VGND VPWR VPWR _35730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32942_ _36015_/CLK _32942_/D VGND VGND VPWR VPWR _32942_/Q sky130_fd_sc_hd__dfxtp_1
X_17876_ _34185_/Q _34121_/Q _34057_/Q _33993_/Q _17799_/X _17800_/X VGND VGND VPWR
+ VPWR _17876_/X sky130_fd_sc_hd__mux4_1
XFILLER_238_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19615_ _19367_/X _19613_/X _19614_/X _19371_/X VGND VGND VPWR VPWR _19615_/X sky130_fd_sc_hd__a22o_1
X_35661_ _35661_/CLK _35661_/D VGND VGND VPWR VPWR _35661_/Q sky130_fd_sc_hd__dfxtp_1
X_16827_ _32875_/Q _32811_/Q _32747_/Q _32683_/Q _16640_/X _16641_/X VGND VGND VPWR
+ VPWR _16827_/X sky130_fd_sc_hd__mux4_1
X_32873_ _32873_/CLK _32873_/D VGND VGND VPWR VPWR _32873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34612_ _34612_/CLK _34612_/D VGND VGND VPWR VPWR _34612_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31824_ _31956_/S VGND VGND VPWR VPWR _31843_/S sky130_fd_sc_hd__buf_4
XFILLER_80_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19546_ _19359_/X _19544_/X _19545_/X _19365_/X VGND VGND VPWR VPWR _19546_/X sky130_fd_sc_hd__a22o_1
X_35592_ _35722_/CLK _35592_/D VGND VGND VPWR VPWR _35592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16758_ _35433_/Q _35369_/Q _35305_/Q _35241_/Q _16548_/X _16549_/X VGND VGND VPWR
+ VPWR _16758_/X sky130_fd_sc_hd__mux4_1
XFILLER_213_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34543_ _36142_/CLK _34543_/D VGND VGND VPWR VPWR _34543_/Q sky130_fd_sc_hd__dfxtp_1
X_31755_ _36085_/Q input25/X _31771_/S VGND VGND VPWR VPWR _31756_/A sky130_fd_sc_hd__mux2_1
X_19477_ _33141_/Q _36021_/Q _33013_/Q _32949_/Q _19362_/X _19363_/X VGND VGND VPWR
+ VPWR _19477_/X sky130_fd_sc_hd__mux4_1
XFILLER_222_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16689_ _16685_/X _16688_/X _16445_/X VGND VGND VPWR VPWR _16697_/C sky130_fd_sc_hd__o21ba_1
XFILLER_224_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_895 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18428_ _33047_/Q _32023_/Q _35799_/Q _35735_/Q _18367_/X _18369_/X VGND VGND VPWR
+ VPWR _18428_/X sky130_fd_sc_hd__mux4_1
XFILLER_179_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30706_ _30706_/A VGND VGND VPWR VPWR _35588_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_1440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34474_ _35180_/CLK _34474_/D VGND VGND VPWR VPWR _34474_/Q sky130_fd_sc_hd__dfxtp_1
X_31686_ _27837_/X _36053_/Q _31686_/S VGND VGND VPWR VPWR _31687_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36213_ _36219_/CLK _36213_/D VGND VGND VPWR VPWR _36213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_912 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33425_ _33425_/CLK _33425_/D VGND VGND VPWR VPWR _33425_/Q sky130_fd_sc_hd__dfxtp_1
X_18359_ _18348_/X _18351_/X _18356_/X _18358_/X VGND VGND VPWR VPWR _18359_/X sky130_fd_sc_hd__a22o_1
X_30637_ _30637_/A VGND VGND VPWR VPWR _35555_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36144_ _36144_/CLK _36144_/D VGND VGND VPWR VPWR _36144_/Q sky130_fd_sc_hd__dfxtp_1
X_33356_ _33420_/CLK _33356_/D VGND VGND VPWR VPWR _33356_/Q sky130_fd_sc_hd__dfxtp_1
X_21370_ _21370_/A VGND VGND VPWR VPWR _36201_/D sky130_fd_sc_hd__clkbuf_1
X_30568_ _35523_/Q _29469_/X _30576_/S VGND VGND VPWR VPWR _30569_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20321_ _20073_/X _20319_/X _20320_/X _20077_/X VGND VGND VPWR VPWR _20321_/X sky130_fd_sc_hd__a22o_1
X_32307_ _35953_/CLK _32307_/D VGND VGND VPWR VPWR _32307_/Q sky130_fd_sc_hd__dfxtp_1
X_36075_ _36075_/CLK _36075_/D VGND VGND VPWR VPWR _36075_/Q sky130_fd_sc_hd__dfxtp_1
X_33287_ _33415_/CLK _33287_/D VGND VGND VPWR VPWR _33287_/Q sky130_fd_sc_hd__dfxtp_1
X_30499_ _35490_/Q _29367_/X _30513_/S VGND VGND VPWR VPWR _30500_/A sky130_fd_sc_hd__mux2_1
X_35026_ _35026_/CLK _35026_/D VGND VGND VPWR VPWR _35026_/Q sky130_fd_sc_hd__dfxtp_1
X_23040_ _23039_/X _32071_/Q _23040_/S VGND VGND VPWR VPWR _23041_/A sky130_fd_sc_hd__mux2_1
X_32238_ _35727_/CLK _32238_/D VGND VGND VPWR VPWR _32238_/Q sky130_fd_sc_hd__dfxtp_1
X_20252_ _20065_/X _20250_/X _20251_/X _20071_/X VGND VGND VPWR VPWR _20252_/X sky130_fd_sc_hd__a22o_1
XFILLER_171_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20183_ _33161_/Q _36041_/Q _33033_/Q _32969_/Q _20068_/X _20069_/X VGND VGND VPWR
+ VPWR _20183_/X sky130_fd_sc_hd__mux4_1
X_32169_ _36137_/CLK _32169_/D VGND VGND VPWR VPWR _32169_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_6_61__f_CLK clkbuf_5_30_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_61__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_24991_ input59/X VGND VGND VPWR VPWR _24991_/X sky130_fd_sc_hd__clkbuf_4
XTAP_4507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26730_ _33798_/Q _23447_/X _26732_/S VGND VGND VPWR VPWR _26731_/A sky130_fd_sc_hd__mux2_1
XTAP_4518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35928_ _35992_/CLK _35928_/D VGND VGND VPWR VPWR _35928_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23942_ _23030_/X _32516_/Q _23948_/S VGND VGND VPWR VPWR _23943_/A sky130_fd_sc_hd__mux2_1
XFILLER_217_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26661_ _33765_/Q _23277_/X _26669_/S VGND VGND VPWR VPWR _26662_/A sky130_fd_sc_hd__mux2_1
X_23873_ _22928_/X _32483_/Q _23885_/S VGND VGND VPWR VPWR _23874_/A sky130_fd_sc_hd__mux2_1
X_35859_ _35859_/CLK _35859_/D VGND VGND VPWR VPWR _35859_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28400_ _27670_/X _34527_/Q _28400_/S VGND VGND VPWR VPWR _28401_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22824_ _20630_/X _22822_/X _22823_/X _20641_/X VGND VGND VPWR VPWR _22824_/X sky130_fd_sc_hd__a22o_1
X_25612_ _25612_/A VGND VGND VPWR VPWR _33270_/D sky130_fd_sc_hd__clkbuf_1
X_29380_ _34982_/Q _29379_/X _29389_/S VGND VGND VPWR VPWR _29381_/A sky130_fd_sc_hd__mux2_1
X_26592_ _26592_/A VGND VGND VPWR VPWR _33734_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28331_ _27766_/X _34494_/Q _28349_/S VGND VGND VPWR VPWR _28332_/A sky130_fd_sc_hd__mux2_1
X_22755_ _22464_/X _22753_/X _22754_/X _22469_/X VGND VGND VPWR VPWR _22755_/X sky130_fd_sc_hd__a22o_1
X_25543_ _25675_/S VGND VGND VPWR VPWR _25562_/S sky130_fd_sc_hd__buf_4
XFILLER_198_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21706_ _21667_/X _21704_/X _21705_/X _21671_/X VGND VGND VPWR VPWR _21706_/X sky130_fd_sc_hd__a22o_1
X_28262_ _28262_/A VGND VGND VPWR VPWR _34461_/D sky130_fd_sc_hd__clkbuf_1
X_25474_ _24896_/X _33205_/Q _25490_/S VGND VGND VPWR VPWR _25475_/A sky130_fd_sc_hd__mux2_1
XFILLER_197_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22686_ _35471_/Q _35407_/Q _35343_/Q _35279_/Q _22560_/X _22561_/X VGND VGND VPWR
+ VPWR _22686_/X sky130_fd_sc_hd__mux4_1
XFILLER_12_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27213_ _27213_/A VGND VGND VPWR VPWR _33999_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_205_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24425_ _24425_/A VGND VGND VPWR VPWR _32741_/D sky130_fd_sc_hd__clkbuf_1
X_21637_ _35633_/Q _34993_/Q _34353_/Q _33713_/Q _21391_/X _21392_/X VGND VGND VPWR
+ VPWR _21637_/X sky130_fd_sc_hd__mux4_1
X_28193_ _27763_/X _34429_/Q _28193_/S VGND VGND VPWR VPWR _28194_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24356_ _23033_/X _32709_/Q _24360_/S VGND VGND VPWR VPWR _24357_/A sky130_fd_sc_hd__mux2_1
X_27144_ _33977_/Q _27143_/X _27156_/S VGND VGND VPWR VPWR _27145_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21568_ _21245_/X _21566_/X _21567_/X _21248_/X VGND VGND VPWR VPWR _21568_/X sky130_fd_sc_hd__a22o_1
XFILLER_5_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23307_ _23307_/A VGND VGND VPWR VPWR _32174_/D sky130_fd_sc_hd__clkbuf_1
X_20519_ _33684_/Q _33620_/Q _33556_/Q _33492_/Q _18324_/X _18325_/X VGND VGND VPWR
+ VPWR _20519_/X sky130_fd_sc_hd__mux4_1
XFILLER_181_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27075_ input5/X VGND VGND VPWR VPWR _27075_/X sky130_fd_sc_hd__buf_4
XFILLER_197_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24287_ _22931_/X _32676_/Q _24297_/S VGND VGND VPWR VPWR _24288_/A sky130_fd_sc_hd__mux2_1
XFILLER_181_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21499_ _35629_/Q _34989_/Q _34349_/Q _33709_/Q _21391_/X _21392_/X VGND VGND VPWR
+ VPWR _21499_/X sky130_fd_sc_hd__mux4_1
XFILLER_101_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23238_ _32152_/Q _23237_/X _23259_/S VGND VGND VPWR VPWR _23239_/A sky130_fd_sc_hd__mux2_1
X_26026_ _24914_/X _33467_/Q _26030_/S VGND VGND VPWR VPWR _26027_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23169_ _23002_/X _32123_/Q _23173_/S VGND VGND VPWR VPWR _23170_/A sky130_fd_sc_hd__mux2_1
XTAP_6421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27977_ _34326_/Q _27033_/X _27995_/S VGND VGND VPWR VPWR _27978_/A sky130_fd_sc_hd__mux2_1
XTAP_5720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15991_ _17910_/A VGND VGND VPWR VPWR _15991_/X sky130_fd_sc_hd__clkbuf_4
XTAP_6476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17730_ _17850_/A VGND VGND VPWR VPWR _17730_/X sky130_fd_sc_hd__buf_4
XFILLER_134_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29716_ _35119_/Q _29407_/X _29724_/S VGND VGND VPWR VPWR _29717_/A sky130_fd_sc_hd__mux2_1
XTAP_6498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26928_ _26928_/A VGND VGND VPWR VPWR _33891_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_236_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29647_ _29647_/A VGND VGND VPWR VPWR _35086_/D sky130_fd_sc_hd__clkbuf_1
X_17661_ _17559_/X _17659_/X _17660_/X _17562_/X VGND VGND VPWR VPWR _17661_/X sky130_fd_sc_hd__a22o_1
XFILLER_236_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26859_ _33859_/Q _23438_/X _26867_/S VGND VGND VPWR VPWR _26860_/A sky130_fd_sc_hd__mux2_1
X_19400_ _19396_/X _19399_/X _19079_/X VGND VGND VPWR VPWR _19422_/A sky130_fd_sc_hd__o21ba_1
XFILLER_35_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16612_ _17800_/A VGND VGND VPWR VPWR _16612_/X sky130_fd_sc_hd__buf_4
X_17592_ _17552_/X _17590_/X _17591_/X _17557_/X VGND VGND VPWR VPWR _17592_/X sky130_fd_sc_hd__a22o_1
X_29578_ _29578_/A VGND VGND VPWR VPWR _35053_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19331_ _19006_/X _19329_/X _19330_/X _19012_/X VGND VGND VPWR VPWR _19331_/X sky130_fd_sc_hd__a22o_1
XFILLER_95_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28529_ _27661_/X _34588_/Q _28535_/S VGND VGND VPWR VPWR _28530_/A sky130_fd_sc_hd__mux2_1
X_16543_ _16361_/X _16541_/X _16542_/X _16365_/X VGND VGND VPWR VPWR _16543_/X sky130_fd_sc_hd__a22o_1
XFILLER_203_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31540_ _31540_/A VGND VGND VPWR VPWR _35983_/D sky130_fd_sc_hd__clkbuf_1
X_19262_ _19014_/X _19260_/X _19261_/X _19018_/X VGND VGND VPWR VPWR _19262_/X sky130_fd_sc_hd__a22o_1
XFILLER_108_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16474_ _32865_/Q _32801_/Q _32737_/Q _32673_/Q _16287_/X _16288_/X VGND VGND VPWR
+ VPWR _16474_/X sky130_fd_sc_hd__mux4_1
XFILLER_93_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18213_ _34451_/Q _36179_/Q _34323_/Q _34259_/Q _17935_/X _17936_/X VGND VGND VPWR
+ VPWR _18213_/X sky130_fd_sc_hd__mux4_1
XFILLER_19_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19193_ _19006_/X _19191_/X _19192_/X _19012_/X VGND VGND VPWR VPWR _19193_/X sky130_fd_sc_hd__a22o_1
X_31471_ _31471_/A VGND VGND VPWR VPWR _35950_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33210_ _33914_/CLK _33210_/D VGND VGND VPWR VPWR _33210_/Q sky130_fd_sc_hd__dfxtp_1
X_18144_ _35665_/Q _35025_/Q _34385_/Q _33745_/Q _17850_/X _17851_/X VGND VGND VPWR
+ VPWR _18144_/X sky130_fd_sc_hd__mux4_1
X_30422_ _30470_/S VGND VGND VPWR VPWR _30441_/S sky130_fd_sc_hd__buf_6
X_34190_ _34192_/CLK _34190_/D VGND VGND VPWR VPWR _34190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33141_ _34485_/CLK _33141_/D VGND VGND VPWR VPWR _33141_/Q sky130_fd_sc_hd__dfxtp_1
X_18075_ _18071_/X _18074_/X _17838_/X VGND VGND VPWR VPWR _18097_/A sky130_fd_sc_hd__o21ba_2
X_30353_ _35421_/Q _29351_/X _30357_/S VGND VGND VPWR VPWR _30354_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17026_ _33905_/Q _33841_/Q _33777_/Q _36081_/Q _17024_/X _17025_/X VGND VGND VPWR
+ VPWR _17026_/X sky130_fd_sc_hd__mux4_1
X_33072_ _36019_/CLK _33072_/D VGND VGND VPWR VPWR _33072_/Q sky130_fd_sc_hd__dfxtp_1
X_30284_ _30284_/A VGND VGND VPWR VPWR _35388_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_217_1102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32023_ _36119_/CLK _32023_/D VGND VGND VPWR VPWR _32023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18977_ _33127_/Q _36007_/Q _32999_/Q _32935_/Q _18656_/X _18657_/X VGND VGND VPWR
+ VPWR _18977_/X sky130_fd_sc_hd__mux4_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17928_ _35466_/Q _35402_/Q _35338_/Q _35274_/Q _17607_/X _17608_/X VGND VGND VPWR
+ VPWR _17928_/X sky130_fd_sc_hd__mux4_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33974_ _34166_/CLK _33974_/D VGND VGND VPWR VPWR _33974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32925_ _36054_/CLK _32925_/D VGND VGND VPWR VPWR _32925_/Q sky130_fd_sc_hd__dfxtp_1
X_35713_ _35713_/CLK _35713_/D VGND VGND VPWR VPWR _35713_/Q sky130_fd_sc_hd__dfxtp_1
X_17859_ _17859_/A VGND VGND VPWR VPWR _17859_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_113_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20870_ _34395_/Q _36123_/Q _34267_/Q _34203_/Q _20770_/X _20771_/X VGND VGND VPWR
+ VPWR _20870_/X sky130_fd_sc_hd__mux4_1
X_32856_ _32856_/CLK _32856_/D VGND VGND VPWR VPWR _32856_/Q sky130_fd_sc_hd__dfxtp_1
X_35644_ _35644_/CLK _35644_/D VGND VGND VPWR VPWR _35644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31807_ _36110_/Q input52/X _31813_/S VGND VGND VPWR VPWR _31808_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19529_ _20235_/A VGND VGND VPWR VPWR _19529_/X sky130_fd_sc_hd__buf_8
X_35575_ _35703_/CLK _35575_/D VGND VGND VPWR VPWR _35575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_1415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32787_ _35922_/CLK _32787_/D VGND VGND VPWR VPWR _32787_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22540_ _22534_/X _22539_/X _22471_/X VGND VGND VPWR VPWR _22541_/D sky130_fd_sc_hd__o21ba_1
X_34526_ _36229_/CLK _34526_/D VGND VGND VPWR VPWR _34526_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31738_ _36077_/Q input16/X _31750_/S VGND VGND VPWR VPWR _31739_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34457_ _34903_/CLK _34457_/D VGND VGND VPWR VPWR _34457_/Q sky130_fd_sc_hd__dfxtp_1
X_22471_ _22471_/A VGND VGND VPWR VPWR _22471_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_887 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31669_ _31669_/A VGND VGND VPWR VPWR _36044_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24210_ _32641_/Q _23432_/X _24222_/S VGND VGND VPWR VPWR _24211_/A sky130_fd_sc_hd__mux2_1
X_33408_ _33921_/CLK _33408_/D VGND VGND VPWR VPWR _33408_/Q sky130_fd_sc_hd__dfxtp_1
X_21422_ _21418_/X _21421_/X _21379_/X VGND VGND VPWR VPWR _21444_/A sky130_fd_sc_hd__o21ba_1
X_25190_ _33072_/Q _23340_/X _25196_/S VGND VGND VPWR VPWR _25191_/A sky130_fd_sc_hd__mux2_1
X_34388_ _35733_/CLK _34388_/D VGND VGND VPWR VPWR _34388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36127_ _36127_/CLK _36127_/D VGND VGND VPWR VPWR _36127_/Q sky130_fd_sc_hd__dfxtp_1
X_24141_ _32608_/Q _23261_/X _24159_/S VGND VGND VPWR VPWR _24142_/A sky130_fd_sc_hd__mux2_1
X_33339_ _36092_/CLK _33339_/D VGND VGND VPWR VPWR _33339_/Q sky130_fd_sc_hd__dfxtp_1
X_21353_ _21314_/X _21351_/X _21352_/X _21318_/X VGND VGND VPWR VPWR _21353_/X sky130_fd_sc_hd__a22o_1
XFILLER_194_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20304_ _34956_/Q _34892_/Q _34828_/Q _34764_/Q _20166_/X _20167_/X VGND VGND VPWR
+ VPWR _20304_/X sky130_fd_sc_hd__mux4_1
XFILLER_200_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36058_ _36058_/CLK _36058_/D VGND VGND VPWR VPWR _36058_/Q sky130_fd_sc_hd__dfxtp_1
X_24072_ _23021_/X _32577_/Q _24084_/S VGND VGND VPWR VPWR _24073_/A sky130_fd_sc_hd__mux2_1
X_21284_ _35623_/Q _34983_/Q _34343_/Q _33703_/Q _21038_/X _21039_/X VGND VGND VPWR
+ VPWR _21284_/X sky130_fd_sc_hd__mux4_1
XFILLER_116_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35009_ _36096_/CLK _35009_/D VGND VGND VPWR VPWR _35009_/Q sky130_fd_sc_hd__dfxtp_1
X_23023_ _23023_/A VGND VGND VPWR VPWR _32065_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27900_ _27729_/X _34290_/Q _27902_/S VGND VGND VPWR VPWR _27901_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20235_ _20235_/A VGND VGND VPWR VPWR _20235_/X sky130_fd_sc_hd__buf_6
X_28880_ _34753_/Q _27168_/X _28892_/S VGND VGND VPWR VPWR _28881_/A sky130_fd_sc_hd__mux2_1
XFILLER_131_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27831_ input58/X VGND VGND VPWR VPWR _27831_/X sky130_fd_sc_hd__clkbuf_4
XTAP_5005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20166_ _20166_/A VGND VGND VPWR VPWR _20166_/X sky130_fd_sc_hd__buf_4
XTAP_5016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27762_ _27762_/A VGND VGND VPWR VPWR _34236_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20097_ _20097_/A VGND VGND VPWR VPWR _32454_/D sky130_fd_sc_hd__clkbuf_4
X_24974_ _24973_/X _32974_/Q _24983_/S VGND VGND VPWR VPWR _24975_/A sky130_fd_sc_hd__mux2_1
XTAP_4326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29501_ _35021_/Q _29500_/X _29513_/S VGND VGND VPWR VPWR _29502_/A sky130_fd_sc_hd__mux2_1
XTAP_4337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26713_ _26761_/S VGND VGND VPWR VPWR _26732_/S sky130_fd_sc_hd__buf_6
XTAP_4348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23925_ _23005_/X _32508_/Q _23927_/S VGND VGND VPWR VPWR _23926_/A sky130_fd_sc_hd__mux2_1
XTAP_3625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27693_ _27692_/X _34214_/Q _27702_/S VGND VGND VPWR VPWR _27694_/A sky130_fd_sc_hd__mux2_1
XTAP_3636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29432_ input27/X VGND VGND VPWR VPWR _29432_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26644_ _33757_/Q _23252_/X _26648_/S VGND VGND VPWR VPWR _26645_/A sky130_fd_sc_hd__mux2_1
XTAP_3658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23856_ _22903_/X _32475_/Q _23864_/S VGND VGND VPWR VPWR _23857_/A sky130_fd_sc_hd__mux2_1
XTAP_3669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_840 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22807_ _33107_/Q _32083_/Q _35859_/Q _35795_/Q _20679_/X _20680_/X VGND VGND VPWR
+ VPWR _22807_/X sky130_fd_sc_hd__mux4_1
X_29363_ _29363_/A VGND VGND VPWR VPWR _34976_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26575_ _24923_/X _33726_/Q _26593_/S VGND VGND VPWR VPWR _26576_/A sky130_fd_sc_hd__mux2_1
XTAP_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20999_ _32863_/Q _32799_/Q _32735_/Q _32671_/Q _20887_/X _20888_/X VGND VGND VPWR
+ VPWR _20999_/X sky130_fd_sc_hd__mux4_1
XFILLER_53_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23787_ _23787_/A VGND VGND VPWR VPWR _32379_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_207_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28314_ _27742_/X _34486_/Q _28328_/S VGND VGND VPWR VPWR _28315_/A sky130_fd_sc_hd__mux2_1
X_25526_ _24973_/X _33230_/Q _25532_/S VGND VGND VPWR VPWR _25527_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29294_ _29294_/A VGND VGND VPWR VPWR _34949_/D sky130_fd_sc_hd__clkbuf_1
X_22738_ _21753_/A _22736_/X _22737_/X _21756_/A VGND VGND VPWR VPWR _22738_/X sky130_fd_sc_hd__a22o_1
XFILLER_246_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28245_ _31418_/B _31823_/B VGND VGND VPWR VPWR _28378_/S sky130_fd_sc_hd__nand2_8
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22669_ _33679_/Q _33615_/Q _33551_/Q _33487_/Q _22506_/X _22507_/X VGND VGND VPWR
+ VPWR _22669_/X sky130_fd_sc_hd__mux4_1
X_25457_ _24871_/X _33197_/Q _25469_/S VGND VGND VPWR VPWR _25458_/A sky130_fd_sc_hd__mux2_1
XFILLER_197_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24408_ _24408_/A VGND VGND VPWR VPWR _32733_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_199_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16190_ _16030_/X _16188_/X _16189_/X _16041_/X VGND VGND VPWR VPWR _16190_/X sky130_fd_sc_hd__a22o_1
XFILLER_187_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28176_ _28176_/A VGND VGND VPWR VPWR _34420_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_205_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25388_ _25388_/A VGND VGND VPWR VPWR _33165_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27127_ input24/X VGND VGND VPWR VPWR _27127_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_51_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24339_ _23008_/X _32701_/Q _24339_/S VGND VGND VPWR VPWR _24340_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_778 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27058_ _27058_/A VGND VGND VPWR VPWR _33949_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18900_ _33381_/Q _33317_/Q _33253_/Q _33189_/Q _18721_/X _18722_/X VGND VGND VPWR
+ VPWR _18900_/X sky130_fd_sc_hd__mux4_1
X_26009_ _24889_/X _33459_/Q _26009_/S VGND VGND VPWR VPWR _26010_/A sky130_fd_sc_hd__mux2_1
X_19880_ _35200_/Q _35136_/Q _35072_/Q _32256_/Q _19663_/X _19664_/X VGND VGND VPWR
+ VPWR _19880_/X sky130_fd_sc_hd__mux4_1
XFILLER_49_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18831_ _33635_/Q _33571_/Q _33507_/Q _33443_/Q _18794_/X _18795_/X VGND VGND VPWR
+ VPWR _18831_/X sky130_fd_sc_hd__mux4_1
XTAP_6240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18762_ _18762_/A VGND VGND VPWR VPWR _32416_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17713_ _17709_/X _17710_/X _17711_/X _17712_/X VGND VGND VPWR VPWR _17713_/X sky130_fd_sc_hd__a22o_1
XFILLER_48_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30971_ _35714_/Q input39/X _30981_/S VGND VGND VPWR VPWR _30972_/A sky130_fd_sc_hd__mux2_1
X_18693_ _18447_/X _18691_/X _18692_/X _18450_/X VGND VGND VPWR VPWR _18693_/X sky130_fd_sc_hd__a22o_1
XFILLER_23_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_291_CLK clkbuf_6_56__f_CLK/X VGND VGND VPWR VPWR _35969_/CLK sky130_fd_sc_hd__clkbuf_16
X_32710_ _32905_/CLK _32710_/D VGND VGND VPWR VPWR _32710_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17644_ _17640_/X _17643_/X _17504_/X VGND VGND VPWR VPWR _17654_/C sky130_fd_sc_hd__o21ba_1
X_33690_ _35610_/CLK _33690_/D VGND VGND VPWR VPWR _33690_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32641_ _36033_/CLK _32641_/D VGND VGND VPWR VPWR _32641_/Q sky130_fd_sc_hd__dfxtp_1
X_17575_ _35456_/Q _35392_/Q _35328_/Q _35264_/Q _17254_/X _17255_/X VGND VGND VPWR
+ VPWR _17575_/X sky130_fd_sc_hd__mux4_1
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19314_ _34416_/Q _36144_/Q _34288_/Q _34224_/Q _19176_/X _19177_/X VGND VGND VPWR
+ VPWR _19314_/X sky130_fd_sc_hd__mux4_1
XFILLER_189_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16526_ _34914_/Q _34850_/Q _34786_/Q _34722_/Q _16454_/X _16455_/X VGND VGND VPWR
+ VPWR _16526_/X sky130_fd_sc_hd__mux4_1
X_35360_ _36005_/CLK _35360_/D VGND VGND VPWR VPWR _35360_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_911 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32572_ _35965_/CLK _32572_/D VGND VGND VPWR VPWR _32572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34311_ _34698_/CLK _34311_/D VGND VGND VPWR VPWR _34311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31523_ _31523_/A VGND VGND VPWR VPWR _35975_/D sky130_fd_sc_hd__clkbuf_1
X_19245_ _34926_/Q _34862_/Q _34798_/Q _34734_/Q _19107_/X _19108_/X VGND VGND VPWR
+ VPWR _19245_/X sky130_fd_sc_hd__mux4_1
XFILLER_231_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35291_ _35802_/CLK _35291_/D VGND VGND VPWR VPWR _35291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16457_ _17163_/A VGND VGND VPWR VPWR _16457_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34242_ _34690_/CLK _34242_/D VGND VGND VPWR VPWR _34242_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19176_ _20016_/A VGND VGND VPWR VPWR _19176_/X sky130_fd_sc_hd__buf_4
X_31454_ _31454_/A VGND VGND VPWR VPWR _35942_/D sky130_fd_sc_hd__clkbuf_1
X_16388_ _17961_/A VGND VGND VPWR VPWR _16388_/X sky130_fd_sc_hd__buf_4
XFILLER_185_870 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18127_ _18127_/A _18127_/B _18127_/C _18127_/D VGND VGND VPWR VPWR _18128_/A sky130_fd_sc_hd__or4_2
X_30405_ _30405_/A VGND VGND VPWR VPWR _35445_/D sky130_fd_sc_hd__clkbuf_1
X_34173_ _34877_/CLK _34173_/D VGND VGND VPWR VPWR _34173_/Q sky130_fd_sc_hd__dfxtp_1
X_31385_ _27791_/X _35910_/Q _31387_/S VGND VGND VPWR VPWR _31386_/A sky130_fd_sc_hd__mux2_1
XFILLER_247_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33124_ _36005_/CLK _33124_/D VGND VGND VPWR VPWR _33124_/Q sky130_fd_sc_hd__dfxtp_1
X_18058_ _16001_/X _18056_/X _18057_/X _16007_/X VGND VGND VPWR VPWR _18058_/X sky130_fd_sc_hd__a22o_1
X_30336_ _30336_/A VGND VGND VPWR VPWR _35413_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17009_ _34672_/Q _34608_/Q _34544_/Q _34480_/Q _16939_/X _16940_/X VGND VGND VPWR
+ VPWR _17009_/X sky130_fd_sc_hd__mux4_1
X_33055_ _35807_/CLK _33055_/D VGND VGND VPWR VPWR _33055_/Q sky130_fd_sc_hd__dfxtp_1
X_30267_ _35380_/Q _29422_/X _30285_/S VGND VGND VPWR VPWR _30268_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20020_ _34436_/Q _36164_/Q _34308_/Q _34244_/Q _19882_/X _19883_/X VGND VGND VPWR
+ VPWR _20020_/X sky130_fd_sc_hd__mux4_1
X_32006_ _36209_/CLK _32006_/D VGND VGND VPWR VPWR _32006_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_876 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30198_ _35348_/Q _29521_/X _30200_/S VGND VGND VPWR VPWR _30199_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_246_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21971_ _21971_/A _21971_/B _21971_/C _21971_/D VGND VGND VPWR VPWR _21972_/A sky130_fd_sc_hd__or4_4
XFILLER_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33957_ _34085_/CLK _33957_/D VGND VGND VPWR VPWR _33957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_282_CLK clkbuf_6_58__f_CLK/X VGND VGND VPWR VPWR _35646_/CLK sky130_fd_sc_hd__clkbuf_16
X_23710_ _23710_/A VGND VGND VPWR VPWR _32342_/D sky130_fd_sc_hd__clkbuf_1
X_20922_ _20916_/X _20921_/X _20615_/X VGND VGND VPWR VPWR _20944_/A sky130_fd_sc_hd__o21ba_1
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24690_ _22928_/X _32867_/Q _24702_/S VGND VGND VPWR VPWR _24691_/A sky130_fd_sc_hd__mux2_1
X_32908_ _32909_/CLK _32908_/D VGND VGND VPWR VPWR _32908_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33888_ _35618_/CLK _33888_/D VGND VGND VPWR VPWR _33888_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20853_ _20618_/X _20851_/X _20852_/X _20627_/X VGND VGND VPWR VPWR _20853_/X sky130_fd_sc_hd__a22o_1
X_32839_ _32903_/CLK _32839_/D VGND VGND VPWR VPWR _32839_/Q sky130_fd_sc_hd__dfxtp_1
X_35627_ _35627_/CLK _35627_/D VGND VGND VPWR VPWR _35627_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23641_ _23641_/A VGND VGND VPWR VPWR _32311_/D sky130_fd_sc_hd__clkbuf_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23572_ _23572_/A VGND VGND VPWR VPWR _32278_/D sky130_fd_sc_hd__clkbuf_1
X_26360_ _26360_/A VGND VGND VPWR VPWR _33624_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20784_ _20780_/X _20783_/X _20615_/X VGND VGND VPWR VPWR _20808_/A sky130_fd_sc_hd__o21ba_1
X_35558_ _35559_/CLK _35558_/D VGND VGND VPWR VPWR _35558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22523_ _22373_/X _22521_/X _22522_/X _22377_/X VGND VGND VPWR VPWR _22523_/X sky130_fd_sc_hd__a22o_1
X_25311_ _33129_/Q _23289_/X _25311_/S VGND VGND VPWR VPWR _25312_/A sky130_fd_sc_hd__mux2_1
XFILLER_222_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34509_ _35213_/CLK _34509_/D VGND VGND VPWR VPWR _34509_/Q sky130_fd_sc_hd__dfxtp_1
X_26291_ _26291_/A VGND VGND VPWR VPWR _33592_/D sky130_fd_sc_hd__clkbuf_1
X_35489_ _35490_/CLK _35489_/D VGND VGND VPWR VPWR _35489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28030_ _28030_/A VGND VGND VPWR VPWR _34351_/D sky130_fd_sc_hd__clkbuf_1
X_22454_ _35464_/Q _35400_/Q _35336_/Q _35272_/Q _22207_/X _22208_/X VGND VGND VPWR
+ VPWR _22454_/X sky130_fd_sc_hd__mux4_1
X_25242_ _25242_/A VGND VGND VPWR VPWR _33096_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21405_ _21758_/A VGND VGND VPWR VPWR _21405_/X sky130_fd_sc_hd__buf_2
XFILLER_182_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25173_ _33064_/Q _23286_/X _25175_/S VGND VGND VPWR VPWR _25174_/A sky130_fd_sc_hd__mux2_1
X_22385_ _22536_/A VGND VGND VPWR VPWR _22385_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_175_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24124_ _32600_/Q _23237_/X _24138_/S VGND VGND VPWR VPWR _24125_/A sky130_fd_sc_hd__mux2_1
X_21336_ _21332_/X _21335_/X _21059_/X VGND VGND VPWR VPWR _21337_/D sky130_fd_sc_hd__o21ba_1
X_29981_ _29981_/A VGND VGND VPWR VPWR _35244_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28932_ _28932_/A VGND VGND VPWR VPWR _34777_/D sky130_fd_sc_hd__clkbuf_1
X_24055_ _22996_/X _32569_/Q _24063_/S VGND VGND VPWR VPWR _24056_/A sky130_fd_sc_hd__mux2_1
X_21267_ _33639_/Q _33575_/Q _33511_/Q _33447_/Q _21094_/X _21095_/X VGND VGND VPWR
+ VPWR _21267_/X sky130_fd_sc_hd__mux4_1
XFILLER_235_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23006_ _23005_/X _32060_/Q _23009_/S VGND VGND VPWR VPWR _23007_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20218_ _32650_/Q _32586_/Q _32522_/Q _35978_/Q _19929_/X _20066_/X VGND VGND VPWR
+ VPWR _20218_/X sky130_fd_sc_hd__mux4_1
XFILLER_235_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28863_ _34745_/Q _27143_/X _28871_/S VGND VGND VPWR VPWR _28864_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21198_ _34149_/Q _34085_/Q _34021_/Q _33957_/Q _20987_/X _20988_/X VGND VGND VPWR
+ VPWR _21198_/X sky130_fd_sc_hd__mux4_1
XFILLER_89_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27814_ _27813_/X _34253_/Q _27826_/S VGND VGND VPWR VPWR _27815_/A sky130_fd_sc_hd__mux2_1
X_20149_ _35720_/Q _32230_/Q _35592_/Q _35528_/Q _19970_/X _19971_/X VGND VGND VPWR
+ VPWR _20149_/X sky130_fd_sc_hd__mux4_1
XTAP_4101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28794_ _34712_/Q _27041_/X _28808_/S VGND VGND VPWR VPWR _28795_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27745_ input27/X VGND VGND VPWR VPWR _27745_/X sky130_fd_sc_hd__buf_2
XTAP_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24957_ _24957_/A VGND VGND VPWR VPWR _32968_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_273_CLK clkbuf_6_57__f_CLK/X VGND VGND VPWR VPWR _35458_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23908_ _23977_/S VGND VGND VPWR VPWR _23927_/S sky130_fd_sc_hd__buf_4
XTAP_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27676_ _27676_/A VGND VGND VPWR VPWR _34208_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24888_ _24888_/A VGND VGND VPWR VPWR _32946_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29415_ _29415_/A VGND VGND VPWR VPWR _34993_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26627_ _26627_/A VGND VGND VPWR VPWR _31688_/B sky130_fd_sc_hd__buf_12
XTAP_3488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23839_ _23839_/A VGND VGND VPWR VPWR _32404_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29346_ _34971_/Q _29345_/X _29358_/S VGND VGND VPWR VPWR _29347_/A sky130_fd_sc_hd__mux2_1
X_17360_ _17356_/X _17357_/X _17358_/X _17359_/X VGND VGND VPWR VPWR _17360_/X sky130_fd_sc_hd__a22o_1
XFILLER_92_1334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_843 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26558_ _24899_/X _33718_/Q _26572_/S VGND VGND VPWR VPWR _26559_/A sky130_fd_sc_hd__mux2_1
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16311_ _16307_/X _16310_/X _16104_/X VGND VGND VPWR VPWR _16312_/D sky130_fd_sc_hd__o21ba_1
XFILLER_201_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25509_ _24948_/X _33222_/Q _25511_/S VGND VGND VPWR VPWR _25510_/A sky130_fd_sc_hd__mux2_1
X_17291_ _17287_/X _17290_/X _17151_/X VGND VGND VPWR VPWR _17301_/C sky130_fd_sc_hd__o21ba_1
X_29277_ _29277_/A VGND VGND VPWR VPWR _34941_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26489_ _26489_/A VGND VGND VPWR VPWR _26622_/S sky130_fd_sc_hd__buf_12
XFILLER_224_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19030_ _34664_/Q _34600_/Q _34536_/Q _34472_/Q _18886_/X _18887_/X VGND VGND VPWR
+ VPWR _19030_/X sky130_fd_sc_hd__mux4_1
X_28228_ _28228_/A VGND VGND VPWR VPWR _34445_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_224_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16242_ _16242_/A _16242_/B _16242_/C _16242_/D VGND VGND VPWR VPWR _16243_/A sky130_fd_sc_hd__or4_1
XFILLER_185_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16173_ _34904_/Q _34840_/Q _34776_/Q _34712_/Q _16096_/X _16098_/X VGND VGND VPWR
+ VPWR _16173_/X sky130_fd_sc_hd__mux4_1
XFILLER_220_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28159_ _28159_/A VGND VGND VPWR VPWR _34412_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput109 _31985_/Q VGND VGND VPWR VPWR D1[27] sky130_fd_sc_hd__buf_2
X_31170_ _31281_/S VGND VGND VPWR VPWR _31189_/S sky130_fd_sc_hd__buf_4
XFILLER_56_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30121_ _35311_/Q _29407_/X _30129_/S VGND VGND VPWR VPWR _30122_/A sky130_fd_sc_hd__mux2_1
X_19932_ _19712_/X _19930_/X _19931_/X _19718_/X VGND VGND VPWR VPWR _19932_/X sky130_fd_sc_hd__a22o_1
XFILLER_141_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_218_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19863_ _19859_/X _19860_/X _19861_/X _19862_/X VGND VGND VPWR VPWR _19863_/X sky130_fd_sc_hd__a22o_1
X_30052_ _30052_/A VGND VGND VPWR VPWR _35278_/D sky130_fd_sc_hd__clkbuf_1
Xoutput91 _31968_/Q VGND VGND VPWR VPWR D1[10] sky130_fd_sc_hd__buf_2
XFILLER_214_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18814_ _35618_/Q _34978_/Q _34338_/Q _33698_/Q _18738_/X _18739_/X VGND VGND VPWR
+ VPWR _18814_/X sky130_fd_sc_hd__mux4_1
XTAP_6070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19794_ _20147_/A VGND VGND VPWR VPWR _19794_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34860_ _35183_/CLK _34860_/D VGND VGND VPWR VPWR _34860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33811_ _36179_/CLK _33811_/D VGND VGND VPWR VPWR _33811_/Q sky130_fd_sc_hd__dfxtp_1
X_18745_ _20157_/A VGND VGND VPWR VPWR _18745_/X sky130_fd_sc_hd__buf_2
XTAP_5380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34791_ _34920_/CLK _34791_/D VGND VGND VPWR VPWR _34791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_264_CLK clkbuf_6_62__f_CLK/X VGND VGND VPWR VPWR _35071_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_188_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33742_ _35663_/CLK _33742_/D VGND VGND VPWR VPWR _33742_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18676_ _18670_/X _18675_/X _18375_/X VGND VGND VPWR VPWR _18684_/C sky130_fd_sc_hd__o21ba_1
X_30954_ _35706_/Q input30/X _30960_/S VGND VGND VPWR VPWR _30955_/A sky130_fd_sc_hd__mux2_1
XTAP_4690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_1267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17627_ _17559_/X _17625_/X _17626_/X _17562_/X VGND VGND VPWR VPWR _17627_/X sky130_fd_sc_hd__a22o_1
X_33673_ _33673_/CLK _33673_/D VGND VGND VPWR VPWR _33673_/Q sky130_fd_sc_hd__dfxtp_1
X_30885_ _35673_/Q input34/X _30897_/S VGND VGND VPWR VPWR _30886_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35412_ _35668_/CLK _35412_/D VGND VGND VPWR VPWR _35412_/Q sky130_fd_sc_hd__dfxtp_1
X_32624_ _36016_/CLK _32624_/D VGND VGND VPWR VPWR _32624_/Q sky130_fd_sc_hd__dfxtp_1
X_17558_ _17552_/X _17555_/X _17556_/X _17557_/X VGND VGND VPWR VPWR _17558_/X sky130_fd_sc_hd__a22o_1
XFILLER_211_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35343_ _35599_/CLK _35343_/D VGND VGND VPWR VPWR _35343_/Q sky130_fd_sc_hd__dfxtp_1
X_16509_ _32098_/Q _32290_/Q _32354_/Q _35874_/Q _16221_/X _16362_/X VGND VGND VPWR
+ VPWR _16509_/X sky130_fd_sc_hd__mux4_1
XFILLER_20_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32555_ _35947_/CLK _32555_/D VGND VGND VPWR VPWR _32555_/Q sky130_fd_sc_hd__dfxtp_1
X_17489_ _17412_/X _17487_/X _17488_/X _17418_/X VGND VGND VPWR VPWR _17489_/X sky130_fd_sc_hd__a22o_1
XFILLER_108_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31506_ _27770_/X _35967_/Q _31522_/S VGND VGND VPWR VPWR _31507_/A sky130_fd_sc_hd__mux2_1
X_19228_ _32110_/Q _32302_/Q _32366_/Q _35886_/Q _19227_/X _19015_/X VGND VGND VPWR
+ VPWR _19228_/X sky130_fd_sc_hd__mux4_1
X_35274_ _35723_/CLK _35274_/D VGND VGND VPWR VPWR _35274_/Q sky130_fd_sc_hd__dfxtp_1
X_32486_ _35944_/CLK _32486_/D VGND VGND VPWR VPWR _32486_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34225_ _36144_/CLK _34225_/D VGND VGND VPWR VPWR _34225_/Q sky130_fd_sc_hd__dfxtp_1
X_31437_ _31437_/A VGND VGND VPWR VPWR _35934_/D sky130_fd_sc_hd__clkbuf_1
X_19159_ _32620_/Q _32556_/Q _32492_/Q _35948_/Q _18870_/X _19007_/X VGND VGND VPWR
+ VPWR _19159_/X sky130_fd_sc_hd__mux4_1
XFILLER_157_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22170_ _22020_/X _22168_/X _22169_/X _22024_/X VGND VGND VPWR VPWR _22170_/X sky130_fd_sc_hd__a22o_1
XFILLER_121_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34156_ _35627_/CLK _34156_/D VGND VGND VPWR VPWR _34156_/Q sky130_fd_sc_hd__dfxtp_1
X_31368_ _31416_/S VGND VGND VPWR VPWR _31387_/S sky130_fd_sc_hd__buf_4
XFILLER_219_1027 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33107_ _35859_/CLK _33107_/D VGND VGND VPWR VPWR _33107_/Q sky130_fd_sc_hd__dfxtp_1
X_21121_ _35170_/Q _35106_/Q _35042_/Q _32162_/Q _20904_/X _20905_/X VGND VGND VPWR
+ VPWR _21121_/X sky130_fd_sc_hd__mux4_1
X_30319_ _35405_/Q _29500_/X _30327_/S VGND VGND VPWR VPWR _30320_/A sky130_fd_sc_hd__mux2_1
X_34087_ _34146_/CLK _34087_/D VGND VGND VPWR VPWR _34087_/Q sky130_fd_sc_hd__dfxtp_1
X_31299_ _27664_/X _35869_/Q _31303_/S VGND VGND VPWR VPWR _31300_/A sky130_fd_sc_hd__mux2_1
X_33038_ _36047_/CLK _33038_/D VGND VGND VPWR VPWR _33038_/Q sky130_fd_sc_hd__dfxtp_1
X_21052_ _21758_/A VGND VGND VPWR VPWR _21052_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_232_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20003_ _19997_/X _20002_/X _19793_/X _19794_/X VGND VGND VPWR VPWR _20024_/B sky130_fd_sc_hd__o211a_1
XFILLER_219_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25860_ _24868_/X _33388_/Q _25874_/S VGND VGND VPWR VPWR _25861_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24811_ _24811_/A VGND VGND VPWR VPWR _32921_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25791_ _25791_/A VGND VGND VPWR VPWR _33355_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34989_ _35693_/CLK _34989_/D VGND VGND VPWR VPWR _34989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_255_CLK clkbuf_6_63__f_CLK/X VGND VGND VPWR VPWR _34180_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_189_1159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27530_ _27530_/A VGND VGND VPWR VPWR _34145_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_215_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24742_ _23005_/X _32892_/Q _24744_/S VGND VGND VPWR VPWR _24743_/A sky130_fd_sc_hd__mux2_1
X_21954_ _22462_/A VGND VGND VPWR VPWR _21954_/X sky130_fd_sc_hd__buf_6
XFILLER_227_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27461_ _34113_/Q _27168_/X _27473_/S VGND VGND VPWR VPWR _27462_/A sky130_fd_sc_hd__mux2_1
X_20905_ _21611_/A VGND VGND VPWR VPWR _20905_/X sky130_fd_sc_hd__buf_6
XFILLER_27_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24673_ _22903_/X _32859_/Q _24681_/S VGND VGND VPWR VPWR _24674_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21885_ _35704_/Q _32213_/Q _35576_/Q _35512_/Q _21564_/X _21565_/X VGND VGND VPWR
+ VPWR _21885_/X sky130_fd_sc_hd__mux4_1
XFILLER_243_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29200_ _29200_/A VGND VGND VPWR VPWR _34904_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_242_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26412_ _26412_/A VGND VGND VPWR VPWR _33649_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20836_ _35162_/Q _35098_/Q _35034_/Q _32154_/Q _20683_/X _20685_/X VGND VGND VPWR
+ VPWR _20836_/X sky130_fd_sc_hd__mux4_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23624_ _23624_/A VGND VGND VPWR VPWR _32303_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_247_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27392_ _34080_/Q _27065_/X _27410_/S VGND VGND VPWR VPWR _27393_/A sky130_fd_sc_hd__mux2_1
XFILLER_242_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29131_ _34872_/Q _27140_/X _29141_/S VGND VGND VPWR VPWR _29132_/A sky130_fd_sc_hd__mux2_1
X_26343_ _26343_/A VGND VGND VPWR VPWR _33617_/D sky130_fd_sc_hd__clkbuf_1
X_20767_ _34648_/Q _34584_/Q _34520_/Q _34456_/Q _20679_/X _20680_/X VGND VGND VPWR
+ VPWR _20767_/X sky130_fd_sc_hd__mux4_1
X_23555_ _32272_/Q _23481_/X _23557_/S VGND VGND VPWR VPWR _23556_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29062_ _34839_/Q _27038_/X _29078_/S VGND VGND VPWR VPWR _29063_/A sky130_fd_sc_hd__mux2_1
X_22506_ _22506_/A VGND VGND VPWR VPWR _22506_/X sky130_fd_sc_hd__buf_6
XFILLER_211_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1018 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23486_ _23486_/A VGND VGND VPWR VPWR _32240_/D sky130_fd_sc_hd__clkbuf_1
X_26274_ _26274_/A VGND VGND VPWR VPWR _33584_/D sky130_fd_sc_hd__clkbuf_1
X_20698_ _21761_/A VGND VGND VPWR VPWR _20698_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_183_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28013_ _28013_/A VGND VGND VPWR VPWR _34343_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22437_ _22159_/X _22435_/X _22436_/X _22162_/X VGND VGND VPWR VPWR _22437_/X sky130_fd_sc_hd__a22o_1
X_25225_ _25225_/A VGND VGND VPWR VPWR _33088_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_1463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22368_ _22586_/A VGND VGND VPWR VPWR _22368_/X sky130_fd_sc_hd__buf_4
XFILLER_136_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25156_ _25267_/S VGND VGND VPWR VPWR _25175_/S sky130_fd_sc_hd__buf_4
XFILLER_174_1406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24107_ _23073_/X _32594_/Q _24113_/S VGND VGND VPWR VPWR _24108_/A sky130_fd_sc_hd__mux2_1
X_21319_ _21314_/X _21316_/X _21317_/X _21318_/X VGND VGND VPWR VPWR _21319_/X sky130_fd_sc_hd__a22o_1
XFILLER_151_534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25087_ _24930_/X _33024_/Q _25101_/S VGND VGND VPWR VPWR _25088_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1081 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29964_ _29964_/A VGND VGND VPWR VPWR _35236_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22299_ _22433_/A VGND VGND VPWR VPWR _22299_/X sky130_fd_sc_hd__buf_4
XFILLER_105_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28915_ _34770_/Q _27220_/X _28921_/S VGND VGND VPWR VPWR _28916_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24038_ _22971_/X _32561_/Q _24042_/S VGND VGND VPWR VPWR _24039_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29895_ _35204_/Q _29472_/X _29901_/S VGND VGND VPWR VPWR _29896_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_494_CLK clkbuf_6_3__f_CLK/X VGND VGND VPWR VPWR _35559_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_77_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28846_ _34737_/Q _27118_/X _28850_/S VGND VGND VPWR VPWR _28847_/A sky130_fd_sc_hd__mux2_1
X_16860_ _33132_/Q _36012_/Q _33004_/Q _32940_/Q _16709_/X _16710_/X VGND VGND VPWR
+ VPWR _16860_/X sky130_fd_sc_hd__mux4_1
XFILLER_172_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28777_ _28777_/A VGND VGND VPWR VPWR _34705_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16791_ _17998_/A VGND VGND VPWR VPWR _16791_/X sky130_fd_sc_hd__buf_6
XFILLER_93_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_924 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25989_ _25989_/A VGND VGND VPWR VPWR _33449_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_246_CLK clkbuf_6_61__f_CLK/X VGND VGND VPWR VPWR _34186_/CLK sky130_fd_sc_hd__clkbuf_16
X_18530_ _33050_/Q _32026_/Q _35802_/Q _35738_/Q _18367_/X _18369_/X VGND VGND VPWR
+ VPWR _18530_/X sky130_fd_sc_hd__mux4_1
XFILLER_150_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27728_ _27728_/A VGND VGND VPWR VPWR _34225_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_776 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18461_ _35608_/Q _34968_/Q _34328_/Q _33688_/Q _18353_/X _18355_/X VGND VGND VPWR
+ VPWR _18461_/X sky130_fd_sc_hd__mux4_1
XFILLER_94_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27659_ _27658_/X _34203_/Q _27671_/S VGND VGND VPWR VPWR _27660_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17412_ _17905_/A VGND VGND VPWR VPWR _17412_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18392_ _20016_/A VGND VGND VPWR VPWR _18392_/X sky130_fd_sc_hd__clkbuf_8
X_30670_ _30670_/A VGND VGND VPWR VPWR _35571_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29329_ _31147_/A _29662_/B VGND VGND VPWR VPWR _29525_/S sky130_fd_sc_hd__nor2_8
Xclkbuf_6_38__f_CLK clkbuf_5_19_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_38__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_17343_ _33146_/Q _36026_/Q _33018_/Q _32954_/Q _17062_/X _17063_/X VGND VGND VPWR
+ VPWR _17343_/X sky130_fd_sc_hd__mux4_1
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32340_ _35989_/CLK _32340_/D VGND VGND VPWR VPWR _32340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17274_ _17206_/X _17272_/X _17273_/X _17209_/X VGND VGND VPWR VPWR _17274_/X sky130_fd_sc_hd__a22o_1
XFILLER_186_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19013_ _19006_/X _19008_/X _19011_/X _19012_/X VGND VGND VPWR VPWR _19013_/X sky130_fd_sc_hd__a22o_1
X_16225_ _16220_/X _16224_/X _16044_/X _16046_/X VGND VGND VPWR VPWR _16242_/B sky130_fd_sc_hd__o211a_1
XFILLER_228_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32271_ _34705_/CLK _32271_/D VGND VGND VPWR VPWR _32271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34010_ _36219_/CLK _34010_/D VGND VGND VPWR VPWR _34010_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31222_ _31222_/A VGND VGND VPWR VPWR _35832_/D sky130_fd_sc_hd__clkbuf_1
X_16156_ _32088_/Q _32280_/Q _32344_/Q _35864_/Q _16032_/X _17867_/A VGND VGND VPWR
+ VPWR _16156_/X sky130_fd_sc_hd__mux4_1
XFILLER_220_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31153_ _31153_/A VGND VGND VPWR VPWR _35799_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16087_ _17771_/A VGND VGND VPWR VPWR _17156_/A sky130_fd_sc_hd__buf_8
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30104_ _35303_/Q _29382_/X _30108_/S VGND VGND VPWR VPWR _30105_/A sky130_fd_sc_hd__mux2_1
X_19915_ _19806_/X _19913_/X _19914_/X _19809_/X VGND VGND VPWR VPWR _19915_/X sky130_fd_sc_hd__a22o_1
XFILLER_114_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31084_ _31084_/A VGND VGND VPWR VPWR _35767_/D sky130_fd_sc_hd__clkbuf_1
X_35961_ _35961_/CLK _35961_/D VGND VGND VPWR VPWR _35961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_485_CLK _35560_/CLK VGND VGND VPWR VPWR _34153_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_29_1386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30035_ _30035_/A VGND VGND VPWR VPWR _35270_/D sky130_fd_sc_hd__clkbuf_1
X_34912_ _34915_/CLK _34912_/D VGND VGND VPWR VPWR _34912_/Q sky130_fd_sc_hd__dfxtp_1
X_19846_ _34431_/Q _36159_/Q _34303_/Q _34239_/Q _19529_/X _19530_/X VGND VGND VPWR
+ VPWR _19846_/X sky130_fd_sc_hd__mux4_1
XFILLER_229_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35892_ _35956_/CLK _35892_/D VGND VGND VPWR VPWR _35892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34843_ _34907_/CLK _34843_/D VGND VGND VPWR VPWR _34843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19777_ _33662_/Q _33598_/Q _33534_/Q _33470_/Q _19500_/X _19501_/X VGND VGND VPWR
+ VPWR _19777_/X sky130_fd_sc_hd__mux4_1
X_16989_ _32624_/Q _32560_/Q _32496_/Q _35952_/Q _16923_/X _16707_/X VGND VGND VPWR
+ VPWR _16989_/X sky130_fd_sc_hd__mux4_1
XFILLER_83_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_237_CLK clkbuf_6_54__f_CLK/X VGND VGND VPWR VPWR _34694_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18728_ _32608_/Q _32544_/Q _32480_/Q _35936_/Q _18517_/X _18654_/X VGND VGND VPWR
+ VPWR _18728_/X sky130_fd_sc_hd__mux4_1
XFILLER_36_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34774_ _34904_/CLK _34774_/D VGND VGND VPWR VPWR _34774_/Q sky130_fd_sc_hd__dfxtp_1
X_31986_ _34914_/CLK _31986_/D VGND VGND VPWR VPWR _31986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18659_ _20210_/A VGND VGND VPWR VPWR _18659_/X sky130_fd_sc_hd__clkbuf_4
X_30937_ _35698_/Q input21/X _30939_/S VGND VGND VPWR VPWR _30938_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33725_ _35645_/CLK _33725_/D VGND VGND VPWR VPWR _33725_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1056 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21670_ _32882_/Q _32818_/Q _32754_/Q _32690_/Q _21593_/X _21594_/X VGND VGND VPWR
+ VPWR _21670_/X sky130_fd_sc_hd__mux4_1
X_30868_ _30868_/A VGND VGND VPWR VPWR _35665_/D sky130_fd_sc_hd__clkbuf_1
X_33656_ _35641_/CLK _33656_/D VGND VGND VPWR VPWR _33656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20621_ _20663_/A VGND VGND VPWR VPWR _22366_/A sky130_fd_sc_hd__buf_12
XFILLER_178_943 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32607_ _35999_/CLK _32607_/D VGND VGND VPWR VPWR _32607_/Q sky130_fd_sc_hd__dfxtp_1
X_33587_ _36082_/CLK _33587_/D VGND VGND VPWR VPWR _33587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30799_ _30799_/A VGND VGND VPWR VPWR _35632_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23340_ input19/X VGND VGND VPWR VPWR _23340_/X sky130_fd_sc_hd__buf_4
X_20552_ _33429_/Q _33365_/Q _33301_/Q _33237_/Q _18337_/X _18339_/X VGND VGND VPWR
+ VPWR _20552_/X sky130_fd_sc_hd__mux4_1
X_32538_ _35995_/CLK _32538_/D VGND VGND VPWR VPWR _32538_/Q sky130_fd_sc_hd__dfxtp_1
X_35326_ _35454_/CLK _35326_/D VGND VGND VPWR VPWR _35326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23271_ input5/X VGND VGND VPWR VPWR _23271_/X sky130_fd_sc_hd__buf_6
X_20483_ _34450_/Q _36178_/Q _34322_/Q _34258_/Q _20235_/X _20236_/X VGND VGND VPWR
+ VPWR _20483_/X sky130_fd_sc_hd__mux4_1
X_32469_ _36076_/CLK _32469_/D VGND VGND VPWR VPWR _32469_/Q sky130_fd_sc_hd__dfxtp_1
X_35257_ _35449_/CLK _35257_/D VGND VGND VPWR VPWR _35257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22222_ _33666_/Q _33602_/Q _33538_/Q _33474_/Q _22153_/X _22154_/X VGND VGND VPWR
+ VPWR _22222_/X sky130_fd_sc_hd__mux4_1
X_25010_ _25010_/A VGND VGND VPWR VPWR _32987_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34208_ _36128_/CLK _34208_/D VGND VGND VPWR VPWR _34208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35188_ _35829_/CLK _35188_/D VGND VGND VPWR VPWR _35188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22153_ _22506_/A VGND VGND VPWR VPWR _22153_/X sky130_fd_sc_hd__buf_4
XFILLER_218_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34139_ _36212_/CLK _34139_/D VGND VGND VPWR VPWR _34139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21104_ _21100_/X _21101_/X _21102_/X _21103_/X VGND VGND VPWR VPWR _21104_/X sky130_fd_sc_hd__a22o_1
XTAP_6817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22084_ _21806_/X _22082_/X _22083_/X _21809_/X VGND VGND VPWR VPWR _22084_/X sky130_fd_sc_hd__a22o_1
XFILLER_121_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26961_ _26961_/A VGND VGND VPWR VPWR _33907_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_476_CLK clkbuf_6_10__f_CLK/X VGND VGND VPWR VPWR _36079_/CLK sky130_fd_sc_hd__clkbuf_16
X_28700_ _28700_/A VGND VGND VPWR VPWR _34668_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_248_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25912_ _24945_/X _33413_/Q _25916_/S VGND VGND VPWR VPWR _25913_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21035_ _22447_/A VGND VGND VPWR VPWR _21035_/X sky130_fd_sc_hd__clkbuf_4
X_29680_ _35102_/Q _29354_/X _29682_/S VGND VGND VPWR VPWR _29681_/A sky130_fd_sc_hd__mux2_1
XFILLER_134_1445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26892_ _33875_/Q _23492_/X _26896_/S VGND VGND VPWR VPWR _26893_/A sky130_fd_sc_hd__mux2_1
XFILLER_232_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28631_ _28631_/A VGND VGND VPWR VPWR _34636_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25843_ _24843_/X _33380_/Q _25853_/S VGND VGND VPWR VPWR _25844_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_228_CLK clkbuf_6_55__f_CLK/X VGND VGND VPWR VPWR _34192_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_216_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28562_ _28562_/A VGND VGND VPWR VPWR _34603_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_234_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25774_ _25774_/A VGND VGND VPWR VPWR _33347_/D sky130_fd_sc_hd__clkbuf_1
X_22986_ _22986_/A VGND VGND VPWR VPWR _32053_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27513_ _27513_/A VGND VGND VPWR VPWR _34137_/D sky130_fd_sc_hd__clkbuf_1
X_24725_ _24794_/S VGND VGND VPWR VPWR _24744_/S sky130_fd_sc_hd__buf_4
XFILLER_55_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28493_ _27807_/X _34571_/Q _28505_/S VGND VGND VPWR VPWR _28494_/A sky130_fd_sc_hd__mux2_1
X_21937_ _21799_/X _21935_/X _21936_/X _21804_/X VGND VGND VPWR VPWR _21937_/X sky130_fd_sc_hd__a22o_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_1254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27444_ _34105_/Q _27143_/X _27452_/S VGND VGND VPWR VPWR _27445_/A sky130_fd_sc_hd__mux2_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24656_ _24656_/A VGND VGND VPWR VPWR _32851_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21868_ _21868_/A VGND VGND VPWR VPWR _36215_/D sky130_fd_sc_hd__buf_6
XFILLER_187_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23607_ _23607_/A VGND VGND VPWR VPWR _32295_/D sky130_fd_sc_hd__clkbuf_1
X_27375_ _34072_/Q _27041_/X _27389_/S VGND VGND VPWR VPWR _27376_/A sky130_fd_sc_hd__mux2_1
X_20819_ _33114_/Q _35994_/Q _32986_/Q _32922_/Q _20624_/X _20625_/X VGND VGND VPWR
+ VPWR _20819_/X sky130_fd_sc_hd__mux4_1
XFILLER_179_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21799_ _22505_/A VGND VGND VPWR VPWR _21799_/X sky130_fd_sc_hd__buf_6
X_24587_ _24587_/A VGND VGND VPWR VPWR _32818_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_1164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_400_CLK clkbuf_6_35__f_CLK/X VGND VGND VPWR VPWR _35446_/CLK sky130_fd_sc_hd__clkbuf_16
X_29114_ _34864_/Q _27115_/X _29120_/S VGND VGND VPWR VPWR _29115_/A sky130_fd_sc_hd__mux2_1
X_26326_ _24958_/X _33609_/Q _26342_/S VGND VGND VPWR VPWR _26327_/A sky130_fd_sc_hd__mux2_1
X_23538_ _23565_/S VGND VGND VPWR VPWR _23557_/S sky130_fd_sc_hd__buf_4
XFILLER_168_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29045_ _29045_/A VGND VGND VPWR VPWR _34831_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26257_ _26257_/A VGND VGND VPWR VPWR _33576_/D sky130_fd_sc_hd__clkbuf_1
X_23469_ input50/X VGND VGND VPWR VPWR _23469_/X sky130_fd_sc_hd__buf_4
XFILLER_195_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16010_ _16063_/A VGND VGND VPWR VPWR _17961_/A sky130_fd_sc_hd__buf_12
XFILLER_155_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25208_ _25208_/A VGND VGND VPWR VPWR _33080_/D sky130_fd_sc_hd__clkbuf_1
X_26188_ _26215_/S VGND VGND VPWR VPWR _26207_/S sky130_fd_sc_hd__buf_4
XFILLER_137_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25139_ _25139_/A VGND VGND VPWR VPWR _33047_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17961_ _17961_/A VGND VGND VPWR VPWR _17961_/X sky130_fd_sc_hd__buf_4
XFILLER_69_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29947_ _29947_/A VGND VGND VPWR VPWR _35228_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19700_ _34939_/Q _34875_/Q _34811_/Q _34747_/Q _19460_/X _19461_/X VGND VGND VPWR
+ VPWR _19700_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_467_CLK clkbuf_6_11__f_CLK/X VGND VGND VPWR VPWR _35183_/CLK sky130_fd_sc_hd__clkbuf_16
X_16912_ _16805_/X _16910_/X _16911_/X _16810_/X VGND VGND VPWR VPWR _16912_/X sky130_fd_sc_hd__a22o_1
X_17892_ _35465_/Q _35401_/Q _35337_/Q _35273_/Q _17607_/X _17608_/X VGND VGND VPWR
+ VPWR _17892_/X sky130_fd_sc_hd__mux4_1
XFILLER_215_1266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29878_ _35196_/Q _29447_/X _29880_/S VGND VGND VPWR VPWR _29879_/A sky130_fd_sc_hd__mux2_1
X_19631_ _19458_/X _19629_/X _19630_/X _19463_/X VGND VGND VPWR VPWR _19631_/X sky130_fd_sc_hd__a22o_1
X_16843_ _16839_/X _16842_/X _16812_/X VGND VGND VPWR VPWR _16844_/D sky130_fd_sc_hd__o21ba_1
X_28829_ _34729_/Q _27093_/X _28829_/S VGND VGND VPWR VPWR _28830_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_219_CLK clkbuf_6_53__f_CLK/X VGND VGND VPWR VPWR _36171_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31840_ _31840_/A VGND VGND VPWR VPWR _36125_/D sky130_fd_sc_hd__clkbuf_1
X_19562_ _19453_/X _19560_/X _19561_/X _19456_/X VGND VGND VPWR VPWR _19562_/X sky130_fd_sc_hd__a22o_1
X_16774_ _17833_/A VGND VGND VPWR VPWR _16774_/X sky130_fd_sc_hd__buf_4
XFILLER_225_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18513_ _33370_/Q _33306_/Q _33242_/Q _33178_/Q _18302_/X _18303_/X VGND VGND VPWR
+ VPWR _18513_/X sky130_fd_sc_hd__mux4_1
XTAP_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31771_ _36093_/Q input33/X _31771_/S VGND VGND VPWR VPWR _31772_/A sky130_fd_sc_hd__mux2_1
X_19493_ _34421_/Q _36149_/Q _34293_/Q _34229_/Q _19176_/X _19177_/X VGND VGND VPWR
+ VPWR _19493_/X sky130_fd_sc_hd__mux4_1
XFILLER_111_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1075 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18444_ _34136_/Q _34072_/Q _34008_/Q _33944_/Q _18309_/X _18311_/X VGND VGND VPWR
+ VPWR _18444_/X sky130_fd_sc_hd__mux4_1
X_30722_ _35596_/Q _29497_/X _30732_/S VGND VGND VPWR VPWR _30723_/A sky130_fd_sc_hd__mux2_1
X_33510_ _34146_/CLK _33510_/D VGND VGND VPWR VPWR _33510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34490_ _35194_/CLK _34490_/D VGND VGND VPWR VPWR _34490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_221_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33441_ _34593_/CLK _33441_/D VGND VGND VPWR VPWR _33441_/Q sky130_fd_sc_hd__dfxtp_1
X_18375_ _20157_/A VGND VGND VPWR VPWR _18375_/X sky130_fd_sc_hd__clkbuf_4
X_30653_ _35563_/Q _29395_/X _30669_/S VGND VGND VPWR VPWR _30654_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1081 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17326_ _34681_/Q _34617_/Q _34553_/Q _34489_/Q _17292_/X _17293_/X VGND VGND VPWR
+ VPWR _17326_/X sky130_fd_sc_hd__mux4_1
X_36160_ _36161_/CLK _36160_/D VGND VGND VPWR VPWR _36160_/Q sky130_fd_sc_hd__dfxtp_1
X_33372_ _36060_/CLK _33372_/D VGND VGND VPWR VPWR _33372_/Q sky130_fd_sc_hd__dfxtp_1
X_30584_ _30584_/A VGND VGND VPWR VPWR _35530_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32323_ _35907_/CLK _32323_/D VGND VGND VPWR VPWR _32323_/Q sky130_fd_sc_hd__dfxtp_1
X_35111_ _35367_/CLK _35111_/D VGND VGND VPWR VPWR _35111_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36091_ _36092_/CLK _36091_/D VGND VGND VPWR VPWR _36091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17257_ _33079_/Q _32055_/Q _35831_/Q _35767_/Q _17078_/X _17079_/X VGND VGND VPWR
+ VPWR _17257_/X sky130_fd_sc_hd__mux4_1
XFILLER_146_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16208_ _16208_/A _16208_/B _16208_/C _16208_/D VGND VGND VPWR VPWR _16209_/A sky130_fd_sc_hd__or4_1
X_35042_ _36197_/CLK _35042_/D VGND VGND VPWR VPWR _35042_/Q sky130_fd_sc_hd__dfxtp_1
X_32254_ _36100_/CLK _32254_/D VGND VGND VPWR VPWR _32254_/Q sky130_fd_sc_hd__dfxtp_1
X_17188_ _17003_/X _17186_/X _17187_/X _17006_/X VGND VGND VPWR VPWR _17188_/X sky130_fd_sc_hd__a22o_1
XFILLER_157_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31205_ _31205_/A VGND VGND VPWR VPWR _35824_/D sky130_fd_sc_hd__clkbuf_1
X_16139_ _16139_/A VGND VGND VPWR VPWR _31959_/D sky130_fd_sc_hd__buf_4
X_32185_ _36129_/CLK _32185_/D VGND VGND VPWR VPWR _32185_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31136_ _31136_/A VGND VGND VPWR VPWR _35792_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_458_CLK clkbuf_leaf_49_CLK/A VGND VGND VPWR VPWR _35754_/CLK sky130_fd_sc_hd__clkbuf_16
X_31067_ _31067_/A VGND VGND VPWR VPWR _35759_/D sky130_fd_sc_hd__clkbuf_1
X_35944_ _35944_/CLK _35944_/D VGND VGND VPWR VPWR _35944_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30018_ _35262_/Q _29453_/X _30036_/S VGND VGND VPWR VPWR _30019_/A sky130_fd_sc_hd__mux2_1
X_19829_ _32639_/Q _32575_/Q _32511_/Q _35967_/Q _19576_/X _19713_/X VGND VGND VPWR
+ VPWR _19829_/X sky130_fd_sc_hd__mux4_1
XFILLER_97_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35875_ _35875_/CLK _35875_/D VGND VGND VPWR VPWR _35875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34826_ _34956_/CLK _34826_/D VGND VGND VPWR VPWR _34826_/Q sky130_fd_sc_hd__dfxtp_1
X_22840_ _34708_/Q _34644_/Q _34580_/Q _34516_/Q _22598_/X _22599_/X VGND VGND VPWR
+ VPWR _22840_/X sky130_fd_sc_hd__mux4_1
XFILLER_83_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34757_ _34949_/CLK _34757_/D VGND VGND VPWR VPWR _34757_/Q sky130_fd_sc_hd__dfxtp_1
X_22771_ _21758_/A _22769_/X _22770_/X _21763_/A VGND VGND VPWR VPWR _22771_/X sky130_fd_sc_hd__a22o_1
XFILLER_65_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31969_ _34085_/CLK _31969_/D VGND VGND VPWR VPWR _31969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24510_ _23061_/X _32782_/Q _24516_/S VGND VGND VPWR VPWR _24511_/A sky130_fd_sc_hd__mux2_1
X_33708_ _35627_/CLK _33708_/D VGND VGND VPWR VPWR _33708_/Q sky130_fd_sc_hd__dfxtp_1
X_21722_ _21722_/A _21722_/B _21722_/C _21722_/D VGND VGND VPWR VPWR _21723_/A sky130_fd_sc_hd__or4_4
X_25490_ _24920_/X _33213_/Q _25490_/S VGND VGND VPWR VPWR _25491_/A sky130_fd_sc_hd__mux2_1
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34688_ _34690_/CLK _34688_/D VGND VGND VPWR VPWR _34688_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21653_ _34162_/Q _34098_/Q _34034_/Q _33970_/Q _21340_/X _21341_/X VGND VGND VPWR
+ VPWR _21653_/X sky130_fd_sc_hd__mux4_1
X_24441_ _22959_/X _32749_/Q _24453_/S VGND VGND VPWR VPWR _24442_/A sky130_fd_sc_hd__mux2_1
X_33639_ _36073_/CLK _33639_/D VGND VGND VPWR VPWR _33639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_21__f_CLK clkbuf_5_10_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_21__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_184_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20604_ _33366_/Q _33302_/Q _33238_/Q _33174_/Q _20602_/X _20603_/X VGND VGND VPWR
+ VPWR _20604_/X sky130_fd_sc_hd__mux4_1
XFILLER_138_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27160_ _33982_/Q _27158_/X _27187_/S VGND VGND VPWR VPWR _27161_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24372_ _24372_/A VGND VGND VPWR VPWR _32716_/D sky130_fd_sc_hd__clkbuf_1
X_21584_ _21446_/X _21582_/X _21583_/X _21451_/X VGND VGND VPWR VPWR _21584_/X sky130_fd_sc_hd__a22o_1
XFILLER_220_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26111_ _24840_/X _33507_/Q _26123_/S VGND VGND VPWR VPWR _26112_/A sky130_fd_sc_hd__mux2_1
X_23323_ _32179_/Q _23240_/X _23335_/S VGND VGND VPWR VPWR _23324_/A sky130_fd_sc_hd__mux2_1
X_20535_ _18281_/X _20533_/X _20534_/X _18291_/X VGND VGND VPWR VPWR _20535_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35309_ _35694_/CLK _35309_/D VGND VGND VPWR VPWR _35309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27091_ _33960_/Q _27090_/X _27094_/S VGND VGND VPWR VPWR _27092_/A sky130_fd_sc_hd__mux2_1
XFILLER_197_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26042_ _26042_/A VGND VGND VPWR VPWR _33474_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23254_ _23254_/A VGND VGND VPWR VPWR _32157_/D sky130_fd_sc_hd__clkbuf_1
X_20466_ _32658_/Q _32594_/Q _32530_/Q _35986_/Q _20282_/X _19177_/A VGND VGND VPWR
+ VPWR _20466_/X sky130_fd_sc_hd__mux4_1
XFILLER_140_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_238_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22205_ _35649_/Q _35009_/Q _34369_/Q _33729_/Q _22097_/X _22098_/X VGND VGND VPWR
+ VPWR _22205_/X sky130_fd_sc_hd__mux4_1
XFILLER_152_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23185_ _23185_/A VGND VGND VPWR VPWR _32130_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20397_ _20397_/A _20397_/B _20397_/C _20397_/D VGND VGND VPWR VPWR _20398_/A sky130_fd_sc_hd__or4_1
XFILLER_134_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29801_ _35159_/Q _29333_/X _29817_/S VGND VGND VPWR VPWR _29802_/A sky130_fd_sc_hd__mux2_1
X_22136_ _35711_/Q _32221_/Q _35583_/Q _35519_/Q _21917_/X _21918_/X VGND VGND VPWR
+ VPWR _22136_/X sky130_fd_sc_hd__mux4_1
XTAP_6614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27993_ _34334_/Q _27059_/X _27995_/S VGND VGND VPWR VPWR _27994_/A sky130_fd_sc_hd__mux2_1
Xoutput270 _32463_/Q VGND VGND VPWR VPWR D3[57] sky130_fd_sc_hd__buf_2
XTAP_6636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput281 _32415_/Q VGND VGND VPWR VPWR D3[9] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_449_CLK clkbuf_6_14__f_CLK/X VGND VGND VPWR VPWR _36013_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_6647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26944_ _33899_/Q _23296_/X _26960_/S VGND VGND VPWR VPWR _26945_/A sky130_fd_sc_hd__mux2_1
X_29732_ _29732_/A VGND VGND VPWR VPWR _35126_/D sky130_fd_sc_hd__clkbuf_1
X_22067_ _22063_/X _22066_/X _21751_/X VGND VGND VPWR VPWR _22075_/C sky130_fd_sc_hd__o21ba_1
XTAP_6669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21018_ _33632_/Q _33568_/Q _33504_/Q _33440_/Q _20741_/X _20742_/X VGND VGND VPWR
+ VPWR _21018_/X sky130_fd_sc_hd__mux4_1
XTAP_5957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29663_ _29795_/S VGND VGND VPWR VPWR _29682_/S sky130_fd_sc_hd__buf_6
XFILLER_181_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26875_ _26875_/A VGND VGND VPWR VPWR _33866_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28614_ _28614_/A VGND VGND VPWR VPWR _34628_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25826_ _24818_/X _33372_/Q _25832_/S VGND VGND VPWR VPWR _25827_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29594_ _35061_/Q _29426_/X _29610_/S VGND VGND VPWR VPWR _29595_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28545_ _28545_/A VGND VGND VPWR VPWR _34595_/D sky130_fd_sc_hd__clkbuf_1
X_25757_ _25757_/A VGND VGND VPWR VPWR _33339_/D sky130_fd_sc_hd__clkbuf_1
X_22969_ _22968_/X _32048_/Q _22978_/S VGND VGND VPWR VPWR _22970_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24708_ _24708_/A VGND VGND VPWR VPWR _32875_/D sky130_fd_sc_hd__clkbuf_1
X_28476_ _27782_/X _34563_/Q _28484_/S VGND VGND VPWR VPWR _28477_/A sky130_fd_sc_hd__mux2_1
X_16490_ _16486_/X _16489_/X _16459_/X VGND VGND VPWR VPWR _16491_/D sky130_fd_sc_hd__o21ba_1
X_25688_ _25688_/A VGND VGND VPWR VPWR _33306_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_203_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1057 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27427_ _34097_/Q _27118_/X _27431_/S VGND VGND VPWR VPWR _27428_/A sky130_fd_sc_hd__mux2_1
X_24639_ _23052_/X _32843_/Q _24651_/S VGND VGND VPWR VPWR _24640_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_941 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18160_ _34194_/Q _34130_/Q _34066_/Q _34002_/Q _16049_/X _16050_/X VGND VGND VPWR
+ VPWR _18160_/X sky130_fd_sc_hd__mux4_1
XFILLER_54_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27358_ _27358_/A VGND VGND VPWR VPWR _34064_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17111_ _35443_/Q _35379_/Q _35315_/Q _35251_/Q _16901_/X _16902_/X VGND VGND VPWR
+ VPWR _17111_/X sky130_fd_sc_hd__mux4_1
X_26309_ _24933_/X _33601_/Q _26321_/S VGND VGND VPWR VPWR _26310_/A sky130_fd_sc_hd__mux2_1
X_18091_ _35215_/Q _35151_/Q _35087_/Q _32271_/Q _16092_/X _16094_/X VGND VGND VPWR
+ VPWR _18091_/X sky130_fd_sc_hd__mux4_1
XFILLER_89_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27289_ _27289_/A VGND VGND VPWR VPWR _34031_/D sky130_fd_sc_hd__clkbuf_1
X_29028_ _29028_/A VGND VGND VPWR VPWR _34823_/D sky130_fd_sc_hd__clkbuf_1
X_17042_ _17038_/X _17041_/X _16798_/X VGND VGND VPWR VPWR _17050_/C sky130_fd_sc_hd__o21ba_1
XFILLER_137_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18993_ _34407_/Q _36135_/Q _34279_/Q _34215_/Q _18823_/X _18824_/X VGND VGND VPWR
+ VPWR _18993_/X sky130_fd_sc_hd__mux4_1
XFILLER_112_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17944_ _34187_/Q _34123_/Q _34059_/Q _33995_/Q _17799_/X _17800_/X VGND VGND VPWR
+ VPWR _17944_/X sky130_fd_sc_hd__mux4_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33990_ _34182_/CLK _33990_/D VGND VGND VPWR VPWR _33990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17875_ _33673_/Q _33609_/Q _33545_/Q _33481_/Q _17553_/X _17554_/X VGND VGND VPWR
+ VPWR _17875_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32941_ _36013_/CLK _32941_/D VGND VGND VPWR VPWR _32941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_215_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_226_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19614_ _32889_/Q _32825_/Q _32761_/Q _32697_/Q _19293_/X _19294_/X VGND VGND VPWR
+ VPWR _19614_/X sky130_fd_sc_hd__mux4_1
X_35660_ _35661_/CLK _35660_/D VGND VGND VPWR VPWR _35660_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16826_ _32107_/Q _32299_/Q _32363_/Q _35883_/Q _16574_/X _16715_/X VGND VGND VPWR
+ VPWR _16826_/X sky130_fd_sc_hd__mux4_1
X_32872_ _32914_/CLK _32872_/D VGND VGND VPWR VPWR _32872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34611_ _34611_/CLK _34611_/D VGND VGND VPWR VPWR _34611_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31823_ _31823_/A _31823_/B VGND VGND VPWR VPWR _31956_/S sky130_fd_sc_hd__nand2_8
X_16757_ _16645_/X _16755_/X _16756_/X _16648_/X VGND VGND VPWR VPWR _16757_/X sky130_fd_sc_hd__a22o_1
XFILLER_59_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19545_ _33143_/Q _36023_/Q _33015_/Q _32951_/Q _19362_/X _19363_/X VGND VGND VPWR
+ VPWR _19545_/X sky130_fd_sc_hd__mux4_1
X_35591_ _35721_/CLK _35591_/D VGND VGND VPWR VPWR _35591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31754_ _31754_/A VGND VGND VPWR VPWR _36084_/D sky130_fd_sc_hd__clkbuf_1
X_34542_ _34926_/CLK _34542_/D VGND VGND VPWR VPWR _34542_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16688_ _16650_/X _16686_/X _16687_/X _16653_/X VGND VGND VPWR VPWR _16688_/X sky130_fd_sc_hd__a22o_1
X_19476_ _32629_/Q _32565_/Q _32501_/Q _35957_/Q _19223_/X _19360_/X VGND VGND VPWR
+ VPWR _19476_/X sky130_fd_sc_hd__mux4_1
XFILLER_206_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30705_ _35588_/Q _29472_/X _30711_/S VGND VGND VPWR VPWR _30706_/A sky130_fd_sc_hd__mux2_1
X_18427_ _35415_/Q _35351_/Q _35287_/Q _35223_/Q _18362_/X _18364_/X VGND VGND VPWR
+ VPWR _18427_/X sky130_fd_sc_hd__mux4_1
XFILLER_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31685_ _31685_/A VGND VGND VPWR VPWR _36052_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34473_ _34913_/CLK _34473_/D VGND VGND VPWR VPWR _34473_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36212_ _36212_/CLK _36212_/D VGND VGND VPWR VPWR _36212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33424_ _34186_/CLK _33424_/D VGND VGND VPWR VPWR _33424_/Q sky130_fd_sc_hd__dfxtp_1
X_18358_ _20162_/A VGND VGND VPWR VPWR _18358_/X sky130_fd_sc_hd__clkbuf_4
X_30636_ _35555_/Q _29370_/X _30648_/S VGND VGND VPWR VPWR _30637_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_5_19_0_CLK clkbuf_2_2_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_19_0_CLK/X sky130_fd_sc_hd__clkbuf_8
X_17309_ _17305_/X _17308_/X _17132_/X VGND VGND VPWR VPWR _17333_/A sky130_fd_sc_hd__o21ba_1
X_33355_ _33420_/CLK _33355_/D VGND VGND VPWR VPWR _33355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36143_ _36143_/CLK _36143_/D VGND VGND VPWR VPWR _36143_/Q sky130_fd_sc_hd__dfxtp_1
X_30567_ _30567_/A VGND VGND VPWR VPWR _35522_/D sky130_fd_sc_hd__clkbuf_1
X_18289_ input79/X input80/X VGND VGND VPWR VPWR _20071_/A sky130_fd_sc_hd__nor2_4
XFILLER_148_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20320_ _32909_/Q _32845_/Q _32781_/Q _32717_/Q _19999_/X _20000_/X VGND VGND VPWR
+ VPWR _20320_/X sky130_fd_sc_hd__mux4_1
X_32306_ _35955_/CLK _32306_/D VGND VGND VPWR VPWR _32306_/Q sky130_fd_sc_hd__dfxtp_1
X_33286_ _33415_/CLK _33286_/D VGND VGND VPWR VPWR _33286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36074_ _36075_/CLK _36074_/D VGND VGND VPWR VPWR _36074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30498_ _30498_/A VGND VGND VPWR VPWR _35489_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35025_ _35731_/CLK _35025_/D VGND VGND VPWR VPWR _35025_/Q sky130_fd_sc_hd__dfxtp_1
X_32237_ _35728_/CLK _32237_/D VGND VGND VPWR VPWR _32237_/Q sky130_fd_sc_hd__dfxtp_1
X_20251_ _33163_/Q _36043_/Q _33035_/Q _32971_/Q _20068_/X _20069_/X VGND VGND VPWR
+ VPWR _20251_/X sky130_fd_sc_hd__mux4_1
XFILLER_190_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20182_ _32649_/Q _32585_/Q _32521_/Q _35977_/Q _19929_/X _20066_/X VGND VGND VPWR
+ VPWR _20182_/X sky130_fd_sc_hd__mux4_1
X_32168_ _36137_/CLK _32168_/D VGND VGND VPWR VPWR _32168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31119_ _35784_/Q input46/X _31137_/S VGND VGND VPWR VPWR _31120_/A sky130_fd_sc_hd__mux2_1
X_24990_ _24990_/A VGND VGND VPWR VPWR _32979_/D sky130_fd_sc_hd__clkbuf_1
X_32099_ _32552_/CLK _32099_/D VGND VGND VPWR VPWR _32099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35927_ _35929_/CLK _35927_/D VGND VGND VPWR VPWR _35927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23941_ _23941_/A VGND VGND VPWR VPWR _32515_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_131_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26660_ _26660_/A VGND VGND VPWR VPWR _33764_/D sky130_fd_sc_hd__clkbuf_1
X_35858_ _35858_/CLK _35858_/D VGND VGND VPWR VPWR _35858_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23872_ _23872_/A VGND VGND VPWR VPWR _32482_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25611_ _24899_/X _33270_/Q _25625_/S VGND VGND VPWR VPWR _25612_/A sky130_fd_sc_hd__mux2_1
X_22823_ _33940_/Q _33876_/Q _33812_/Q _36116_/Q _20662_/X _20664_/X VGND VGND VPWR
+ VPWR _22823_/X sky130_fd_sc_hd__mux4_1
X_34809_ _35769_/CLK _34809_/D VGND VGND VPWR VPWR _34809_/Q sky130_fd_sc_hd__dfxtp_1
X_26591_ _24948_/X _33734_/Q _26593_/S VGND VGND VPWR VPWR _26592_/A sky130_fd_sc_hd__mux2_1
X_35789_ _35852_/CLK _35789_/D VGND VGND VPWR VPWR _35789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_232_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28330_ _28378_/S VGND VGND VPWR VPWR _28349_/S sky130_fd_sc_hd__buf_4
XFILLER_53_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25542_ _27840_/A _26352_/B VGND VGND VPWR VPWR _25675_/S sky130_fd_sc_hd__nand2_8
XFILLER_25_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22754_ _34961_/Q _34897_/Q _34833_/Q _34769_/Q _22466_/X _22467_/X VGND VGND VPWR
+ VPWR _22754_/X sky130_fd_sc_hd__mux4_1
XFILLER_225_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28261_ _27664_/X _34461_/Q _28265_/S VGND VGND VPWR VPWR _28262_/A sky130_fd_sc_hd__mux2_1
X_21705_ _32883_/Q _32819_/Q _32755_/Q _32691_/Q _21593_/X _21594_/X VGND VGND VPWR
+ VPWR _21705_/X sky130_fd_sc_hd__mux4_1
X_25473_ _25473_/A VGND VGND VPWR VPWR _33204_/D sky130_fd_sc_hd__clkbuf_1
X_22685_ _20581_/X _22683_/X _22684_/X _20591_/X VGND VGND VPWR VPWR _22685_/X sky130_fd_sc_hd__a22o_1
XFILLER_200_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27212_ _33999_/Q _27211_/X _27218_/S VGND VGND VPWR VPWR _27213_/A sky130_fd_sc_hd__mux2_1
XFILLER_197_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24424_ _22934_/X _32741_/Q _24432_/S VGND VGND VPWR VPWR _24425_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21636_ _35697_/Q _32205_/Q _35569_/Q _35505_/Q _21564_/X _21565_/X VGND VGND VPWR
+ VPWR _21636_/X sky130_fd_sc_hd__mux4_1
X_28192_ _28192_/A VGND VGND VPWR VPWR _34428_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27143_ input29/X VGND VGND VPWR VPWR _27143_/X sky130_fd_sc_hd__buf_2
XFILLER_51_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24355_ _24355_/A VGND VGND VPWR VPWR _32708_/D sky130_fd_sc_hd__clkbuf_1
X_21567_ _35631_/Q _34991_/Q _34351_/Q _33711_/Q _21391_/X _21392_/X VGND VGND VPWR
+ VPWR _21567_/X sky130_fd_sc_hd__mux4_1
XFILLER_20_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23306_ _32174_/Q _23305_/X _23424_/S VGND VGND VPWR VPWR _23307_/A sky130_fd_sc_hd__mux2_1
X_20518_ _20518_/A VGND VGND VPWR VPWR _32467_/D sky130_fd_sc_hd__clkbuf_4
X_27074_ _27074_/A VGND VGND VPWR VPWR _33954_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_1271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24286_ _24286_/A VGND VGND VPWR VPWR _32675_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21498_ _35693_/Q _32201_/Q _35565_/Q _35501_/Q _21211_/X _21212_/X VGND VGND VPWR
+ VPWR _21498_/X sky130_fd_sc_hd__mux4_1
XFILLER_107_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26025_ _26025_/A VGND VGND VPWR VPWR _33466_/D sky130_fd_sc_hd__clkbuf_1
X_23237_ input23/X VGND VGND VPWR VPWR _23237_/X sky130_fd_sc_hd__clkbuf_4
X_20449_ _20445_/X _20448_/X _20157_/X VGND VGND VPWR VPWR _20457_/C sky130_fd_sc_hd__o21ba_1
XTAP_7101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23168_ _23168_/A VGND VGND VPWR VPWR _32122_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22119_ _22110_/X _22117_/X _22118_/X VGND VGND VPWR VPWR _22120_/D sky130_fd_sc_hd__o21ba_1
XTAP_5710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23099_ _23099_/A VGND VGND VPWR VPWR _32089_/D sky130_fd_sc_hd__clkbuf_1
X_15990_ _17771_/A VGND VGND VPWR VPWR _17910_/A sky130_fd_sc_hd__buf_12
X_27976_ _28108_/S VGND VGND VPWR VPWR _27995_/S sky130_fd_sc_hd__buf_4
XTAP_6455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26927_ _33891_/Q _23271_/X _26939_/S VGND VGND VPWR VPWR _26928_/A sky130_fd_sc_hd__mux2_1
X_29715_ _29715_/A VGND VGND VPWR VPWR _35118_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_890 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17660_ _33923_/Q _33859_/Q _33795_/Q _36099_/Q _17377_/X _17378_/X VGND VGND VPWR
+ VPWR _17660_/X sky130_fd_sc_hd__mux4_1
XTAP_5798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29646_ _35086_/Q _29503_/X _29652_/S VGND VGND VPWR VPWR _29647_/A sky130_fd_sc_hd__mux2_1
X_26858_ _26858_/A VGND VGND VPWR VPWR _33858_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16611_ _17799_/A VGND VGND VPWR VPWR _16611_/X sky130_fd_sc_hd__buf_4
X_25809_ _25809_/A VGND VGND VPWR VPWR _33364_/D sky130_fd_sc_hd__clkbuf_1
X_17591_ _34177_/Q _34113_/Q _34049_/Q _33985_/Q _17446_/X _17447_/X VGND VGND VPWR
+ VPWR _17591_/X sky130_fd_sc_hd__mux4_1
X_29577_ _35053_/Q _29401_/X _29589_/S VGND VGND VPWR VPWR _29578_/A sky130_fd_sc_hd__mux2_1
XFILLER_223_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_972 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26789_ _26789_/A VGND VGND VPWR VPWR _33825_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28528_ _28528_/A VGND VGND VPWR VPWR _34587_/D sky130_fd_sc_hd__clkbuf_1
X_16542_ _32867_/Q _32803_/Q _32739_/Q _32675_/Q _16287_/X _16288_/X VGND VGND VPWR
+ VPWR _16542_/X sky130_fd_sc_hd__mux4_1
X_19330_ _33137_/Q _36017_/Q _33009_/Q _32945_/Q _19009_/X _19010_/X VGND VGND VPWR
+ VPWR _19330_/X sky130_fd_sc_hd__mux4_1
XFILLER_16_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19261_ _32879_/Q _32815_/Q _32751_/Q _32687_/Q _18940_/X _18941_/X VGND VGND VPWR
+ VPWR _19261_/X sky130_fd_sc_hd__mux4_1
X_16473_ _32097_/Q _32289_/Q _32353_/Q _35873_/Q _16221_/X _16362_/X VGND VGND VPWR
+ VPWR _16473_/X sky130_fd_sc_hd__mux4_1
X_28459_ _27757_/X _34555_/Q _28463_/S VGND VGND VPWR VPWR _28460_/A sky130_fd_sc_hd__mux2_1
XFILLER_232_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18212_ _16048_/X _18210_/X _18211_/X _16058_/X VGND VGND VPWR VPWR _18212_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19192_ _33133_/Q _36013_/Q _33005_/Q _32941_/Q _19009_/X _19010_/X VGND VGND VPWR
+ VPWR _19192_/X sky130_fd_sc_hd__mux4_1
X_31470_ _27717_/X _35950_/Q _31480_/S VGND VGND VPWR VPWR _31471_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18143_ _35729_/Q _32240_/Q _35601_/Q _35537_/Q _15993_/X _15995_/X VGND VGND VPWR
+ VPWR _18143_/X sky130_fd_sc_hd__mux4_1
XFILLER_141_1032 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30421_ _30421_/A VGND VGND VPWR VPWR _35453_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33140_ _36021_/CLK _33140_/D VGND VGND VPWR VPWR _33140_/Q sky130_fd_sc_hd__dfxtp_1
X_18074_ _17912_/X _18072_/X _18073_/X _17915_/X VGND VGND VPWR VPWR _18074_/X sky130_fd_sc_hd__a22o_1
X_30352_ _30352_/A VGND VGND VPWR VPWR _35420_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17025_ _17851_/A VGND VGND VPWR VPWR _17025_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_67_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_908 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33071_ _36144_/CLK _33071_/D VGND VGND VPWR VPWR _33071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_236_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30283_ _35388_/Q _29447_/X _30285_/S VGND VGND VPWR VPWR _30284_/A sky130_fd_sc_hd__mux2_1
X_32022_ _36119_/CLK _32022_/D VGND VGND VPWR VPWR _32022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18976_ _32615_/Q _32551_/Q _32487_/Q _35943_/Q _18870_/X _18654_/X VGND VGND VPWR
+ VPWR _18976_/X sky130_fd_sc_hd__mux4_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17927_ _17704_/X _17925_/X _17926_/X _17707_/X VGND VGND VPWR VPWR _17927_/X sky130_fd_sc_hd__a22o_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33973_ _34101_/CLK _33973_/D VGND VGND VPWR VPWR _33973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35712_ _35713_/CLK _35712_/D VGND VGND VPWR VPWR _35712_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32924_ _36054_/CLK _32924_/D VGND VGND VPWR VPWR _32924_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17858_ _17853_/X _17856_/X _17857_/X VGND VGND VPWR VPWR _17873_/C sky130_fd_sc_hd__o21ba_1
XFILLER_226_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16809_ _34922_/Q _34858_/Q _34794_/Q _34730_/Q _16807_/X _16808_/X VGND VGND VPWR
+ VPWR _16809_/X sky130_fd_sc_hd__mux4_1
XFILLER_54_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35643_ _35644_/CLK _35643_/D VGND VGND VPWR VPWR _35643_/Q sky130_fd_sc_hd__dfxtp_1
X_32855_ _35221_/CLK _32855_/D VGND VGND VPWR VPWR _32855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17789_ _34694_/Q _34630_/Q _34566_/Q _34502_/Q _17645_/X _17646_/X VGND VGND VPWR
+ VPWR _17789_/X sky130_fd_sc_hd__mux4_1
XFILLER_35_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31806_ _31806_/A VGND VGND VPWR VPWR _36109_/D sky130_fd_sc_hd__clkbuf_1
X_19528_ _19453_/X _19526_/X _19527_/X _19456_/X VGND VGND VPWR VPWR _19528_/X sky130_fd_sc_hd__a22o_1
X_35574_ _35701_/CLK _35574_/D VGND VGND VPWR VPWR _35574_/Q sky130_fd_sc_hd__dfxtp_1
X_32786_ _32914_/CLK _32786_/D VGND VGND VPWR VPWR _32786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_5_2_0_CLK clkbuf_5_7_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_2_0_CLK/X sky130_fd_sc_hd__clkbuf_8
X_34525_ _36229_/CLK _34525_/D VGND VGND VPWR VPWR _34525_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31737_ _31737_/A VGND VGND VPWR VPWR _36076_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19459_ _34420_/Q _36148_/Q _34292_/Q _34228_/Q _19176_/X _19177_/X VGND VGND VPWR
+ VPWR _19459_/X sky130_fd_sc_hd__mux4_1
XFILLER_34_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34456_ _34903_/CLK _34456_/D VGND VGND VPWR VPWR _34456_/Q sky130_fd_sc_hd__dfxtp_1
X_22470_ _22464_/X _22465_/X _22468_/X _22469_/X VGND VGND VPWR VPWR _22470_/X sky130_fd_sc_hd__a22o_1
XFILLER_195_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31668_ _27810_/X _36044_/Q _31678_/S VGND VGND VPWR VPWR _31669_/A sky130_fd_sc_hd__mux2_1
X_33407_ _35648_/CLK _33407_/D VGND VGND VPWR VPWR _33407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21421_ _21100_/X _21419_/X _21420_/X _21103_/X VGND VGND VPWR VPWR _21421_/X sky130_fd_sc_hd__a22o_1
X_30619_ _35547_/Q _29345_/X _30627_/S VGND VGND VPWR VPWR _30620_/A sky130_fd_sc_hd__mux2_1
X_34387_ _35730_/CLK _34387_/D VGND VGND VPWR VPWR _34387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31599_ _27708_/X _36011_/Q _31615_/S VGND VGND VPWR VPWR _31600_/A sky130_fd_sc_hd__mux2_1
XFILLER_202_1449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36126_ _36229_/CLK _36126_/D VGND VGND VPWR VPWR _36126_/Q sky130_fd_sc_hd__dfxtp_1
X_24140_ _24251_/S VGND VGND VPWR VPWR _24159_/S sky130_fd_sc_hd__buf_4
X_21352_ _32873_/Q _32809_/Q _32745_/Q _32681_/Q _21240_/X _21241_/X VGND VGND VPWR
+ VPWR _21352_/X sky130_fd_sc_hd__mux4_1
X_33338_ _33914_/CLK _33338_/D VGND VGND VPWR VPWR _33338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20303_ _34444_/Q _36172_/Q _34316_/Q _34252_/Q _20235_/X _20236_/X VGND VGND VPWR
+ VPWR _20303_/X sky130_fd_sc_hd__mux4_1
XFILLER_147_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36057_ _36057_/CLK _36057_/D VGND VGND VPWR VPWR _36057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24071_ _24071_/A VGND VGND VPWR VPWR _32576_/D sky130_fd_sc_hd__clkbuf_1
X_21283_ _35687_/Q _32194_/Q _35559_/Q _35495_/Q _21211_/X _21212_/X VGND VGND VPWR
+ VPWR _21283_/X sky130_fd_sc_hd__mux4_1
X_33269_ _34100_/CLK _33269_/D VGND VGND VPWR VPWR _33269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20234_ _20159_/X _20232_/X _20233_/X _20162_/X VGND VGND VPWR VPWR _20234_/X sky130_fd_sc_hd__a22o_1
X_35008_ _36096_/CLK _35008_/D VGND VGND VPWR VPWR _35008_/Q sky130_fd_sc_hd__dfxtp_1
X_23022_ _23021_/X _32065_/Q _23040_/S VGND VGND VPWR VPWR _23023_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_1023 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27830_ _27830_/A VGND VGND VPWR VPWR _34258_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20165_ _34440_/Q _36168_/Q _34312_/Q _34248_/Q _19882_/X _19883_/X VGND VGND VPWR
+ VPWR _20165_/X sky130_fd_sc_hd__mux4_1
XTAP_5006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27761_ _27760_/X _34236_/Q _27764_/S VGND VGND VPWR VPWR _27762_/A sky130_fd_sc_hd__mux2_1
X_24973_ input52/X VGND VGND VPWR VPWR _24973_/X sky130_fd_sc_hd__buf_4
X_20096_ _20096_/A _20096_/B _20096_/C _20096_/D VGND VGND VPWR VPWR _20097_/A sky130_fd_sc_hd__or4_1
XTAP_4305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29500_ input51/X VGND VGND VPWR VPWR _29500_/X sky130_fd_sc_hd__buf_2
XTAP_4338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26712_ _26712_/A VGND VGND VPWR VPWR _33789_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23924_ _23924_/A VGND VGND VPWR VPWR _32507_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27692_ input8/X VGND VGND VPWR VPWR _27692_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_85_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29431_ _29431_/A VGND VGND VPWR VPWR _34998_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26643_ _26643_/A VGND VGND VPWR VPWR _33756_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23855_ _23855_/A VGND VGND VPWR VPWR _32474_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22806_ _35475_/Q _35411_/Q _35347_/Q _35283_/Q _22560_/X _22561_/X VGND VGND VPWR
+ VPWR _22806_/X sky130_fd_sc_hd__mux4_1
XFILLER_26_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29362_ _34976_/Q _29360_/X _29389_/S VGND VGND VPWR VPWR _29363_/A sky130_fd_sc_hd__mux2_1
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_791 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26574_ _26622_/S VGND VGND VPWR VPWR _26593_/S sky130_fd_sc_hd__buf_4
XTAP_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23786_ _23002_/X _32379_/Q _23790_/S VGND VGND VPWR VPWR _23787_/A sky130_fd_sc_hd__mux2_1
X_20998_ _32095_/Q _32287_/Q _32351_/Q _35871_/Q _20821_/X _20962_/X VGND VGND VPWR
+ VPWR _20998_/X sky130_fd_sc_hd__mux4_1
XFILLER_77_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28313_ _28313_/A VGND VGND VPWR VPWR _34485_/D sky130_fd_sc_hd__clkbuf_1
X_25525_ _25525_/A VGND VGND VPWR VPWR _33229_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_246_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_750 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29293_ _34949_/Q _27180_/X _29297_/S VGND VGND VPWR VPWR _29294_/A sky130_fd_sc_hd__mux2_1
X_22737_ _33169_/Q _36049_/Q _33041_/Q _32977_/Q _20632_/X _21761_/A VGND VGND VPWR
+ VPWR _22737_/X sky130_fd_sc_hd__mux4_1
XFILLER_40_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28244_ _28244_/A VGND VGND VPWR VPWR _34453_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25456_ _25456_/A VGND VGND VPWR VPWR _33196_/D sky130_fd_sc_hd__clkbuf_1
X_22668_ _22668_/A VGND VGND VPWR VPWR _36238_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24407_ _22909_/X _32733_/Q _24411_/S VGND VGND VPWR VPWR _24408_/A sky130_fd_sc_hd__mux2_1
X_21619_ _21619_/A VGND VGND VPWR VPWR _36208_/D sky130_fd_sc_hd__clkbuf_1
X_28175_ _27735_/X _34420_/Q _28193_/S VGND VGND VPWR VPWR _28176_/A sky130_fd_sc_hd__mux2_1
X_25387_ _33165_/Q _23472_/X _25395_/S VGND VGND VPWR VPWR _25388_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22599_ _22599_/A VGND VGND VPWR VPWR _22599_/X sky130_fd_sc_hd__buf_4
XFILLER_16_1377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27126_ _27126_/A VGND VGND VPWR VPWR _33971_/D sky130_fd_sc_hd__clkbuf_1
X_24338_ _24338_/A VGND VGND VPWR VPWR _32700_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27057_ _33949_/Q _27056_/X _27063_/S VGND VGND VPWR VPWR _27058_/A sky130_fd_sc_hd__mux2_1
X_24269_ _24269_/A VGND VGND VPWR VPWR _32667_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26008_ _26008_/A VGND VGND VPWR VPWR _33458_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_941 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18830_ _18830_/A VGND VGND VPWR VPWR _32418_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1036 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18761_ _18761_/A _18761_/B _18761_/C _18761_/D VGND VGND VPWR VPWR _18762_/A sky130_fd_sc_hd__or4_2
X_27959_ _27816_/X _34318_/Q _27965_/S VGND VGND VPWR VPWR _27960_/A sky130_fd_sc_hd__mux2_1
XTAP_6285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17712_ _17869_/A VGND VGND VPWR VPWR _17712_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_248_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30970_ _30970_/A VGND VGND VPWR VPWR _35713_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_903 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_222_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18692_ _33887_/Q _33823_/Q _33759_/Q _36063_/Q _18618_/X _18619_/X VGND VGND VPWR
+ VPWR _18692_/X sky130_fd_sc_hd__mux4_1
XFILLER_114_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29629_ _35078_/Q _29478_/X _29631_/S VGND VGND VPWR VPWR _29630_/A sky130_fd_sc_hd__mux2_1
XTAP_4883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17643_ _17356_/X _17641_/X _17642_/X _17359_/X VGND VGND VPWR VPWR _17643_/X sky130_fd_sc_hd__a22o_1
XFILLER_184_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17574_ _17351_/X _17572_/X _17573_/X _17354_/X VGND VGND VPWR VPWR _17574_/X sky130_fd_sc_hd__a22o_1
X_32640_ _36030_/CLK _32640_/D VGND VGND VPWR VPWR _32640_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19313_ _19100_/X _19309_/X _19312_/X _19103_/X VGND VGND VPWR VPWR _19313_/X sky130_fd_sc_hd__a22o_1
X_16525_ _34402_/Q _36130_/Q _34274_/Q _34210_/Q _16523_/X _16524_/X VGND VGND VPWR
+ VPWR _16525_/X sky130_fd_sc_hd__mux4_1
XFILLER_95_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32571_ _36027_/CLK _32571_/D VGND VGND VPWR VPWR _32571_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34310_ _34694_/CLK _34310_/D VGND VGND VPWR VPWR _34310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31522_ _27794_/X _35975_/Q _31522_/S VGND VGND VPWR VPWR _31523_/A sky130_fd_sc_hd__mux2_1
X_16456_ _34912_/Q _34848_/Q _34784_/Q _34720_/Q _16454_/X _16455_/X VGND VGND VPWR
+ VPWR _16456_/X sky130_fd_sc_hd__mux4_1
X_19244_ _34414_/Q _36142_/Q _34286_/Q _34222_/Q _19176_/X _19177_/X VGND VGND VPWR
+ VPWR _19244_/X sky130_fd_sc_hd__mux4_1
X_35290_ _35802_/CLK _35290_/D VGND VGND VPWR VPWR _35290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34241_ _34690_/CLK _34241_/D VGND VGND VPWR VPWR _34241_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19175_ _19100_/X _19173_/X _19174_/X _19103_/X VGND VGND VPWR VPWR _19175_/X sky130_fd_sc_hd__a22o_1
X_31453_ _27692_/X _35942_/Q _31459_/S VGND VGND VPWR VPWR _31454_/A sky130_fd_sc_hd__mux2_1
X_16387_ _17960_/A VGND VGND VPWR VPWR _16387_/X sky130_fd_sc_hd__buf_6
XFILLER_121_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18126_ _18122_/X _18125_/X _17871_/X VGND VGND VPWR VPWR _18127_/D sky130_fd_sc_hd__o21ba_1
XFILLER_160_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30404_ _35445_/Q _29426_/X _30420_/S VGND VGND VPWR VPWR _30405_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34172_ _34172_/CLK _34172_/D VGND VGND VPWR VPWR _34172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31384_ _31384_/A VGND VGND VPWR VPWR _35909_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30335_ _35413_/Q _29524_/X _30335_/S VGND VGND VPWR VPWR _30336_/A sky130_fd_sc_hd__mux2_1
X_18057_ _33102_/Q _32078_/Q _35854_/Q _35790_/Q _17784_/X _17785_/X VGND VGND VPWR
+ VPWR _18057_/X sky130_fd_sc_hd__mux4_1
X_33123_ _36003_/CLK _33123_/D VGND VGND VPWR VPWR _33123_/Q sky130_fd_sc_hd__dfxtp_1
X_17008_ _17002_/X _17007_/X _16798_/X VGND VGND VPWR VPWR _17018_/C sky130_fd_sc_hd__o21ba_1
XFILLER_67_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33054_ _33119_/CLK _33054_/D VGND VGND VPWR VPWR _33054_/Q sky130_fd_sc_hd__dfxtp_1
X_30266_ _30335_/S VGND VGND VPWR VPWR _30285_/S sky130_fd_sc_hd__buf_6
XFILLER_116_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32005_ _36202_/CLK _32005_/D VGND VGND VPWR VPWR _32005_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30197_ _30197_/A VGND VGND VPWR VPWR _35347_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18959_ _35174_/Q _35110_/Q _35046_/Q _32166_/Q _18957_/X _18958_/X VGND VGND VPWR
+ VPWR _18959_/X sky130_fd_sc_hd__mux4_1
XFILLER_100_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33956_ _34148_/CLK _33956_/D VGND VGND VPWR VPWR _33956_/Q sky130_fd_sc_hd__dfxtp_1
X_21970_ _21966_/X _21969_/X _21765_/X VGND VGND VPWR VPWR _21971_/D sky130_fd_sc_hd__o21ba_1
XFILLER_239_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20921_ _20747_/X _20917_/X _20920_/X _20750_/X VGND VGND VPWR VPWR _20921_/X sky130_fd_sc_hd__a22o_1
X_32907_ _32907_/CLK _32907_/D VGND VGND VPWR VPWR _32907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33887_ _35551_/CLK _33887_/D VGND VGND VPWR VPWR _33887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35626_ _35693_/CLK _35626_/D VGND VGND VPWR VPWR _35626_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23640_ _22990_/X _32311_/Q _23652_/S VGND VGND VPWR VPWR _23641_/A sky130_fd_sc_hd__mux2_1
X_20852_ _33115_/Q _35995_/Q _32987_/Q _32923_/Q _20624_/X _20625_/X VGND VGND VPWR
+ VPWR _20852_/X sky130_fd_sc_hd__mux4_1
X_32838_ _32905_/CLK _32838_/D VGND VGND VPWR VPWR _32838_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23571_ _22879_/X _32278_/Q _23589_/S VGND VGND VPWR VPWR _23572_/A sky130_fd_sc_hd__mux2_1
X_35557_ _35625_/CLK _35557_/D VGND VGND VPWR VPWR _35557_/Q sky130_fd_sc_hd__dfxtp_1
X_20783_ _20747_/X _20781_/X _20782_/X _20750_/X VGND VGND VPWR VPWR _20783_/X sky130_fd_sc_hd__a22o_1
X_32769_ _35902_/CLK _32769_/D VGND VGND VPWR VPWR _32769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25310_ _25310_/A VGND VGND VPWR VPWR _33128_/D sky130_fd_sc_hd__clkbuf_1
X_34508_ _35147_/CLK _34508_/D VGND VGND VPWR VPWR _34508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22522_ _32906_/Q _32842_/Q _32778_/Q _32714_/Q _22299_/X _22300_/X VGND VGND VPWR
+ VPWR _22522_/X sky130_fd_sc_hd__mux4_1
X_26290_ _24905_/X _33592_/Q _26300_/S VGND VGND VPWR VPWR _26291_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35488_ _35747_/CLK _35488_/D VGND VGND VPWR VPWR _35488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25241_ _33096_/Q _23453_/X _25259_/S VGND VGND VPWR VPWR _25242_/A sky130_fd_sc_hd__mux2_1
X_34439_ _36167_/CLK _34439_/D VGND VGND VPWR VPWR _34439_/Q sky130_fd_sc_hd__dfxtp_1
X_22453_ _22304_/X _22449_/X _22452_/X _22307_/X VGND VGND VPWR VPWR _22453_/X sky130_fd_sc_hd__a22o_1
X_21404_ _21400_/X _21401_/X _21402_/X _21403_/X VGND VGND VPWR VPWR _21404_/X sky130_fd_sc_hd__a22o_1
X_25172_ _25172_/A VGND VGND VPWR VPWR _33063_/D sky130_fd_sc_hd__clkbuf_1
X_22384_ _22535_/A VGND VGND VPWR VPWR _22384_/X sky130_fd_sc_hd__buf_6
XFILLER_191_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36109_ _36109_/CLK _36109_/D VGND VGND VPWR VPWR _36109_/Q sky130_fd_sc_hd__dfxtp_1
X_24123_ _24123_/A VGND VGND VPWR VPWR _32599_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21335_ _21052_/X _21333_/X _21334_/X _21057_/X VGND VGND VPWR VPWR _21335_/X sky130_fd_sc_hd__a22o_1
XFILLER_203_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29980_ _35244_/Q _29398_/X _29994_/S VGND VGND VPWR VPWR _29981_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28931_ _34777_/Q _27044_/X _28943_/S VGND VGND VPWR VPWR _28932_/A sky130_fd_sc_hd__mux2_1
X_24054_ _24054_/A VGND VGND VPWR VPWR _32568_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21266_ _21266_/A VGND VGND VPWR VPWR _36198_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_1326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23005_ input32/X VGND VGND VPWR VPWR _23005_/X sky130_fd_sc_hd__buf_2
X_20217_ _20211_/X _20216_/X _20138_/X VGND VGND VPWR VPWR _20241_/A sky130_fd_sc_hd__o21ba_2
XFILLER_172_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21197_ _33637_/Q _33573_/Q _33509_/Q _33445_/Q _21094_/X _21095_/X VGND VGND VPWR
+ VPWR _21197_/X sky130_fd_sc_hd__mux4_1
X_28862_ _28862_/A VGND VGND VPWR VPWR _34744_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27813_ input51/X VGND VGND VPWR VPWR _27813_/X sky130_fd_sc_hd__clkbuf_4
X_20148_ _20142_/X _20145_/X _20146_/X _20147_/X VGND VGND VPWR VPWR _20173_/B sky130_fd_sc_hd__o211a_1
X_28793_ _28793_/A VGND VGND VPWR VPWR _34711_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24956_ _24954_/X _32968_/Q _24983_/S VGND VGND VPWR VPWR _24957_/A sky130_fd_sc_hd__mux2_1
X_20079_ _20072_/X _20078_/X _19793_/X _19794_/X VGND VGND VPWR VPWR _20096_/B sky130_fd_sc_hd__o211a_1
XTAP_4135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27744_ _27744_/A VGND VGND VPWR VPWR _34230_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23907_ _23907_/A VGND VGND VPWR VPWR _32499_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27675_ _27673_/X _34208_/Q _27702_/S VGND VGND VPWR VPWR _27676_/A sky130_fd_sc_hd__mux2_1
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24887_ _24886_/X _32946_/Q _24890_/S VGND VGND VPWR VPWR _24888_/A sky130_fd_sc_hd__mux2_1
XTAP_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26626_ input87/X input86/X input88/X VGND VGND VPWR VPWR _26627_/A sky130_fd_sc_hd__or3b_1
XTAP_3478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29414_ _34993_/Q _29413_/X _29420_/S VGND VGND VPWR VPWR _29415_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23838_ _23079_/X _32404_/Q _23840_/S VGND VGND VPWR VPWR _23839_/A sky130_fd_sc_hd__mux2_1
XTAP_3489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29345_ input56/X VGND VGND VPWR VPWR _29345_/X sky130_fd_sc_hd__clkbuf_4
X_26557_ _26557_/A VGND VGND VPWR VPWR _33717_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23769_ _22977_/X _32371_/Q _23769_/S VGND VGND VPWR VPWR _23770_/A sky130_fd_sc_hd__mux2_1
XFILLER_202_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16310_ _16091_/X _16308_/X _16309_/X _16101_/X VGND VGND VPWR VPWR _16310_/X sky130_fd_sc_hd__a22o_1
XFILLER_198_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25508_ _25508_/A VGND VGND VPWR VPWR _33221_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17290_ _17003_/X _17288_/X _17289_/X _17006_/X VGND VGND VPWR VPWR _17290_/X sky130_fd_sc_hd__a22o_1
X_29276_ _34941_/Q _27155_/X _29276_/S VGND VGND VPWR VPWR _29277_/A sky130_fd_sc_hd__mux2_1
X_26488_ _31147_/A _30472_/A VGND VGND VPWR VPWR _26489_/A sky130_fd_sc_hd__or2_1
XFILLER_158_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28227_ _27813_/X _34445_/Q _28235_/S VGND VGND VPWR VPWR _28228_/A sky130_fd_sc_hd__mux2_1
X_16241_ _16237_/X _16240_/X _16104_/X VGND VGND VPWR VPWR _16242_/D sky130_fd_sc_hd__o21ba_1
X_25439_ _25439_/A VGND VGND VPWR VPWR _33188_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16172_ _34392_/Q _36120_/Q _34264_/Q _34200_/Q _16170_/X _16171_/X VGND VGND VPWR
+ VPWR _16172_/X sky130_fd_sc_hd__mux4_1
XFILLER_16_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28158_ _27711_/X _34412_/Q _28172_/S VGND VGND VPWR VPWR _28159_/A sky130_fd_sc_hd__mux2_1
XFILLER_220_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27109_ input17/X VGND VGND VPWR VPWR _27109_/X sky130_fd_sc_hd__buf_2
XFILLER_103_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28089_ _28089_/A VGND VGND VPWR VPWR _34379_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30120_ _30120_/A VGND VGND VPWR VPWR _35310_/D sky130_fd_sc_hd__clkbuf_1
X_19931_ _33154_/Q _36034_/Q _33026_/Q _32962_/Q _19715_/X _19716_/X VGND VGND VPWR
+ VPWR _19931_/X sky130_fd_sc_hd__mux4_1
X_30051_ _35278_/Q _29503_/X _30057_/S VGND VGND VPWR VPWR _30052_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19862_ _20215_/A VGND VGND VPWR VPWR _19862_/X sky130_fd_sc_hd__buf_4
XFILLER_190_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput92 _31969_/Q VGND VGND VPWR VPWR D1[11] sky130_fd_sc_hd__buf_2
X_18813_ _35682_/Q _32189_/Q _35554_/Q _35490_/Q _18558_/X _18559_/X VGND VGND VPWR
+ VPWR _18813_/X sky130_fd_sc_hd__mux4_1
XTAP_6060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_847 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19793_ _20146_/A VGND VGND VPWR VPWR _19793_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_68_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33810_ _36179_/CLK _33810_/D VGND VGND VPWR VPWR _33810_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18744_ _18597_/X _18742_/X _18743_/X _18600_/X VGND VGND VPWR VPWR _18744_/X sky130_fd_sc_hd__a22o_1
XTAP_5370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34790_ _34790_/CLK _34790_/D VGND VGND VPWR VPWR _34790_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33741_ _35661_/CLK _33741_/D VGND VGND VPWR VPWR _33741_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18675_ _18597_/X _18671_/X _18674_/X _18600_/X VGND VGND VPWR VPWR _18675_/X sky130_fd_sc_hd__a22o_1
XFILLER_23_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30953_ _30953_/A VGND VGND VPWR VPWR _35705_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_237_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17626_ _33922_/Q _33858_/Q _33794_/Q _36098_/Q _17377_/X _17378_/X VGND VGND VPWR
+ VPWR _17626_/X sky130_fd_sc_hd__mux4_1
XFILLER_36_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33672_ _33673_/CLK _33672_/D VGND VGND VPWR VPWR _33672_/Q sky130_fd_sc_hd__dfxtp_1
X_30884_ _30884_/A VGND VGND VPWR VPWR _35672_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35411_ _35666_/CLK _35411_/D VGND VGND VPWR VPWR _35411_/Q sky130_fd_sc_hd__dfxtp_1
X_32623_ _36015_/CLK _32623_/D VGND VGND VPWR VPWR _32623_/Q sky130_fd_sc_hd__dfxtp_1
X_17557_ _17910_/A VGND VGND VPWR VPWR _17557_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_211_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35342_ _35855_/CLK _35342_/D VGND VGND VPWR VPWR _35342_/Q sky130_fd_sc_hd__dfxtp_1
X_16508_ _16353_/X _16506_/X _16507_/X _16359_/X VGND VGND VPWR VPWR _16508_/X sky130_fd_sc_hd__a22o_1
X_17488_ _33150_/Q _36030_/Q _33022_/Q _32958_/Q _17415_/X _17416_/X VGND VGND VPWR
+ VPWR _17488_/X sky130_fd_sc_hd__mux4_1
X_32554_ _35883_/CLK _32554_/D VGND VGND VPWR VPWR _32554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31505_ _31505_/A VGND VGND VPWR VPWR _35966_/D sky130_fd_sc_hd__clkbuf_1
X_19227_ _20286_/A VGND VGND VPWR VPWR _19227_/X sky130_fd_sc_hd__buf_4
XFILLER_220_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35273_ _35466_/CLK _35273_/D VGND VGND VPWR VPWR _35273_/Q sky130_fd_sc_hd__dfxtp_1
X_16439_ _17999_/A VGND VGND VPWR VPWR _16439_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_34_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32485_ _35943_/CLK _32485_/D VGND VGND VPWR VPWR _32485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34224_ _36144_/CLK _34224_/D VGND VGND VPWR VPWR _34224_/Q sky130_fd_sc_hd__dfxtp_1
X_31436_ _27667_/X _35934_/Q _31438_/S VGND VGND VPWR VPWR _31437_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19158_ _19152_/X _19157_/X _19079_/X VGND VGND VPWR VPWR _19182_/A sky130_fd_sc_hd__o21ba_1
XFILLER_173_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18109_ _32144_/Q _32336_/Q _32400_/Q _35920_/Q _17986_/X _17011_/A VGND VGND VPWR
+ VPWR _18109_/X sky130_fd_sc_hd__mux4_1
X_34155_ _35627_/CLK _34155_/D VGND VGND VPWR VPWR _34155_/Q sky130_fd_sc_hd__dfxtp_1
X_31367_ _31367_/A VGND VGND VPWR VPWR _35901_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_219_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19089_ _19083_/X _19086_/X _19087_/X _19088_/X VGND VGND VPWR VPWR _19114_/B sky130_fd_sc_hd__o211a_1
XFILLER_219_1039 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30318_ _30318_/A VGND VGND VPWR VPWR _35404_/D sky130_fd_sc_hd__clkbuf_1
X_33106_ _35859_/CLK _33106_/D VGND VGND VPWR VPWR _33106_/Q sky130_fd_sc_hd__dfxtp_1
X_21120_ _34658_/Q _34594_/Q _34530_/Q _34466_/Q _20833_/X _20834_/X VGND VGND VPWR
+ VPWR _21120_/X sky130_fd_sc_hd__mux4_1
XFILLER_156_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31298_ _31298_/A VGND VGND VPWR VPWR _35868_/D sky130_fd_sc_hd__clkbuf_1
X_34086_ _34790_/CLK _34086_/D VGND VGND VPWR VPWR _34086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21051_ _21047_/X _21048_/X _21049_/X _21050_/X VGND VGND VPWR VPWR _21051_/X sky130_fd_sc_hd__a22o_1
X_33037_ _35853_/CLK _33037_/D VGND VGND VPWR VPWR _33037_/Q sky130_fd_sc_hd__dfxtp_1
X_30249_ _30249_/A VGND VGND VPWR VPWR _35371_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20002_ _19720_/X _19998_/X _20001_/X _19724_/X VGND VGND VPWR VPWR _20002_/X sky130_fd_sc_hd__a22o_1
XFILLER_8_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24810_ _24809_/X _32921_/Q _24828_/S VGND VGND VPWR VPWR _24811_/A sky130_fd_sc_hd__mux2_1
X_25790_ _24964_/X _33355_/Q _25802_/S VGND VGND VPWR VPWR _25791_/A sky130_fd_sc_hd__mux2_1
X_34988_ _35692_/CLK _34988_/D VGND VGND VPWR VPWR _34988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24741_ _24741_/A VGND VGND VPWR VPWR _32891_/D sky130_fd_sc_hd__clkbuf_1
X_33939_ _36177_/CLK _33939_/D VGND VGND VPWR VPWR _33939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21953_ _35642_/Q _35002_/Q _34362_/Q _33722_/Q _21744_/X _21745_/X VGND VGND VPWR
+ VPWR _21953_/X sky130_fd_sc_hd__mux4_1
XFILLER_28_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27460_ _27460_/A VGND VGND VPWR VPWR _34112_/D sky130_fd_sc_hd__clkbuf_1
X_20904_ _22316_/A VGND VGND VPWR VPWR _20904_/X sky130_fd_sc_hd__buf_6
X_24672_ _24672_/A VGND VGND VPWR VPWR _32858_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21884_ _21879_/X _21883_/X _21740_/X _21741_/X VGND VGND VPWR VPWR _21901_/B sky130_fd_sc_hd__o211a_1
XFILLER_203_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26411_ _33649_/Q _23364_/X _26415_/S VGND VGND VPWR VPWR _26412_/A sky130_fd_sc_hd__mux2_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35609_ _35609_/CLK _35609_/D VGND VGND VPWR VPWR _35609_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23623_ _22965_/X _32303_/Q _23631_/S VGND VGND VPWR VPWR _23624_/A sky130_fd_sc_hd__mux2_1
X_20835_ _34650_/Q _34586_/Q _34522_/Q _34458_/Q _20833_/X _20834_/X VGND VGND VPWR
+ VPWR _20835_/X sky130_fd_sc_hd__mux4_1
X_27391_ _27502_/S VGND VGND VPWR VPWR _27410_/S sky130_fd_sc_hd__buf_6
XFILLER_153_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29130_ _29130_/A VGND VGND VPWR VPWR _34871_/D sky130_fd_sc_hd__clkbuf_1
X_26342_ _24982_/X _33617_/Q _26342_/S VGND VGND VPWR VPWR _26343_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23554_ _23554_/A VGND VGND VPWR VPWR _32271_/D sky130_fd_sc_hd__clkbuf_1
X_20766_ _20762_/X _20765_/X _20675_/X VGND VGND VPWR VPWR _20776_/C sky130_fd_sc_hd__o21ba_1
XFILLER_11_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29061_ _29061_/A VGND VGND VPWR VPWR _34838_/D sky130_fd_sc_hd__clkbuf_1
X_22505_ _22505_/A VGND VGND VPWR VPWR _22505_/X sky130_fd_sc_hd__buf_4
X_26273_ _24880_/X _33584_/Q _26279_/S VGND VGND VPWR VPWR _26274_/A sky130_fd_sc_hd__mux2_1
X_23485_ _32240_/Q _23484_/X _23485_/S VGND VGND VPWR VPWR _23486_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20697_ _22374_/A VGND VGND VPWR VPWR _21761_/A sky130_fd_sc_hd__buf_12
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28012_ _34343_/Q _27087_/X _28016_/S VGND VGND VPWR VPWR _28013_/A sky130_fd_sc_hd__mux2_1
XFILLER_202_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25224_ _33088_/Q _23429_/X _25238_/S VGND VGND VPWR VPWR _25225_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22436_ _33928_/Q _33864_/Q _33800_/Q _36104_/Q _22330_/X _22331_/X VGND VGND VPWR
+ VPWR _22436_/X sky130_fd_sc_hd__mux4_1
XFILLER_104_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25155_ _25155_/A VGND VGND VPWR VPWR _33055_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_191_CLK clkbuf_6_48__f_CLK/X VGND VGND VPWR VPWR _36045_/CLK sky130_fd_sc_hd__clkbuf_16
X_22367_ _32646_/Q _32582_/Q _32518_/Q _35974_/Q _22229_/X _22366_/X VGND VGND VPWR
+ VPWR _22367_/X sky130_fd_sc_hd__mux4_1
XFILLER_191_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24106_ _24106_/A VGND VGND VPWR VPWR _32593_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21318_ _22515_/A VGND VGND VPWR VPWR _21318_/X sky130_fd_sc_hd__clkbuf_4
X_25086_ _25086_/A VGND VGND VPWR VPWR _33023_/D sky130_fd_sc_hd__clkbuf_1
X_29963_ _35236_/Q _29373_/X _29973_/S VGND VGND VPWR VPWR _29964_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22298_ _32132_/Q _32324_/Q _32388_/Q _35908_/Q _22233_/X _22021_/X VGND VGND VPWR
+ VPWR _22298_/X sky130_fd_sc_hd__mux4_1
XFILLER_11_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28914_ _28914_/A VGND VGND VPWR VPWR _34769_/D sky130_fd_sc_hd__clkbuf_1
X_24037_ _24037_/A VGND VGND VPWR VPWR _32560_/D sky130_fd_sc_hd__clkbuf_1
X_21249_ _21245_/X _21246_/X _21247_/X _21248_/X VGND VGND VPWR VPWR _21249_/X sky130_fd_sc_hd__a22o_1
X_29894_ _29894_/A VGND VGND VPWR VPWR _35203_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_836 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28845_ _28845_/A VGND VGND VPWR VPWR _34736_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16790_ _35690_/Q _32197_/Q _35562_/Q _35498_/Q _16611_/X _16612_/X VGND VGND VPWR
+ VPWR _16790_/X sky130_fd_sc_hd__mux4_1
X_28776_ _34705_/Q _27217_/X _28776_/S VGND VGND VPWR VPWR _28777_/A sky130_fd_sc_hd__mux2_1
X_25988_ _24858_/X _33449_/Q _25988_/S VGND VGND VPWR VPWR _25989_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_936 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24939_ input40/X VGND VGND VPWR VPWR _24939_/X sky130_fd_sc_hd__buf_4
X_27727_ _27726_/X _34225_/Q _27733_/S VGND VGND VPWR VPWR _27728_/A sky130_fd_sc_hd__mux2_1
XTAP_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18460_ _35672_/Q _32178_/Q _35544_/Q _35480_/Q _18349_/X _18350_/X VGND VGND VPWR
+ VPWR _18460_/X sky130_fd_sc_hd__mux4_1
XFILLER_61_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27658_ input56/X VGND VGND VPWR VPWR _27658_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_46_788 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17411_ _17407_/X _17410_/X _17132_/X VGND VGND VPWR VPWR _17443_/A sky130_fd_sc_hd__o21ba_1
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18391_ _19458_/A VGND VGND VPWR VPWR _18391_/X sky130_fd_sc_hd__clkbuf_4
X_26609_ _26609_/A VGND VGND VPWR VPWR _33742_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27589_ _27637_/S VGND VGND VPWR VPWR _27608_/S sky130_fd_sc_hd__buf_6
XFILLER_221_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ _32634_/Q _32570_/Q _32506_/Q _35962_/Q _17276_/X _17060_/X VGND VGND VPWR
+ VPWR _17342_/X sky130_fd_sc_hd__mux4_1
X_29328_ input1/X VGND VGND VPWR VPWR _29328_/X sky130_fd_sc_hd__buf_2
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17273_ _33912_/Q _33848_/Q _33784_/Q _36088_/Q _17024_/X _17025_/X VGND VGND VPWR
+ VPWR _17273_/X sky130_fd_sc_hd__mux4_1
XFILLER_144_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29259_ _29259_/A VGND VGND VPWR VPWR _34932_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16224_ _16030_/X _16222_/X _16223_/X _16041_/X VGND VGND VPWR VPWR _16224_/X sky130_fd_sc_hd__a22o_1
X_19012_ _20210_/A VGND VGND VPWR VPWR _19012_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_201_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32270_ _36114_/CLK _32270_/D VGND VGND VPWR VPWR _32270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_1165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31221_ _27748_/X _35832_/Q _31231_/S VGND VGND VPWR VPWR _31222_/A sky130_fd_sc_hd__mux2_1
X_16155_ _16018_/X _16153_/X _16154_/X _16027_/X VGND VGND VPWR VPWR _16155_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_182_CLK clkbuf_6_27__f_CLK/X VGND VGND VPWR VPWR _35855_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_6_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31152_ _27646_/X _35799_/Q _31168_/S VGND VGND VPWR VPWR _31153_/A sky130_fd_sc_hd__mux2_1
X_16086_ _35158_/Q _35094_/Q _35030_/Q _32150_/Q _16083_/X _16085_/X VGND VGND VPWR
+ VPWR _16086_/X sky130_fd_sc_hd__mux4_1
XFILLER_154_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1086 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30103_ _30103_/A VGND VGND VPWR VPWR _35302_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19914_ _35201_/Q _35137_/Q _35073_/Q _32257_/Q _19663_/X _19664_/X VGND VGND VPWR
+ VPWR _19914_/X sky130_fd_sc_hd__mux4_1
XFILLER_64_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31083_ _35767_/Q input27/X _31095_/S VGND VGND VPWR VPWR _31084_/A sky130_fd_sc_hd__mux2_1
X_35960_ _35961_/CLK _35960_/D VGND VGND VPWR VPWR _35960_/Q sky130_fd_sc_hd__dfxtp_1
X_34911_ _34911_/CLK _34911_/D VGND VGND VPWR VPWR _34911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_218_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30034_ _35270_/Q _29478_/X _30036_/S VGND VGND VPWR VPWR _30035_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19845_ _19806_/X _19843_/X _19844_/X _19809_/X VGND VGND VPWR VPWR _19845_/X sky130_fd_sc_hd__a22o_1
XFILLER_64_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35891_ _35953_/CLK _35891_/D VGND VGND VPWR VPWR _35891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34842_ _36245_/CLK _34842_/D VGND VGND VPWR VPWR _34842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19776_ _19776_/A VGND VGND VPWR VPWR _32445_/D sky130_fd_sc_hd__clkbuf_4
X_16988_ _16984_/X _16987_/X _16779_/X VGND VGND VPWR VPWR _17018_/A sky130_fd_sc_hd__o21ba_1
X_18727_ _18720_/X _18725_/X _18726_/X VGND VGND VPWR VPWR _18761_/A sky130_fd_sc_hd__o21ba_1
XFILLER_110_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34773_ _34773_/CLK _34773_/D VGND VGND VPWR VPWR _34773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_823 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31985_ _34918_/CLK _31985_/D VGND VGND VPWR VPWR _31985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_1002 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_917 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33724_ _35645_/CLK _33724_/D VGND VGND VPWR VPWR _33724_/Q sky130_fd_sc_hd__dfxtp_1
X_18658_ _33118_/Q _35998_/Q _32990_/Q _32926_/Q _18656_/X _18657_/X VGND VGND VPWR
+ VPWR _18658_/X sky130_fd_sc_hd__mux4_1
X_30936_ _30936_/A VGND VGND VPWR VPWR _35697_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17609_ _35457_/Q _35393_/Q _35329_/Q _35265_/Q _17607_/X _17608_/X VGND VGND VPWR
+ VPWR _17609_/X sky130_fd_sc_hd__mux4_1
XFILLER_52_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33655_ _34166_/CLK _33655_/D VGND VGND VPWR VPWR _33655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30867_ _35665_/Q input55/X _30867_/S VGND VGND VPWR VPWR _30868_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18589_ _32860_/Q _32796_/Q _32732_/Q _32668_/Q _18587_/X _18588_/X VGND VGND VPWR
+ VPWR _18589_/X sky130_fd_sc_hd__mux4_1
XFILLER_51_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32606_ _35999_/CLK _32606_/D VGND VGND VPWR VPWR _32606_/Q sky130_fd_sc_hd__dfxtp_1
X_20620_ _22582_/A VGND VGND VPWR VPWR _22466_/A sky130_fd_sc_hd__buf_12
XFILLER_189_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33586_ _34098_/CLK _33586_/D VGND VGND VPWR VPWR _33586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30798_ _35632_/Q input19/X _30804_/S VGND VGND VPWR VPWR _30799_/A sky130_fd_sc_hd__mux2_1
X_35325_ _36029_/CLK _35325_/D VGND VGND VPWR VPWR _35325_/Q sky130_fd_sc_hd__dfxtp_1
X_20551_ _18318_/X _20549_/X _20550_/X _18327_/X VGND VGND VPWR VPWR _20551_/X sky130_fd_sc_hd__a22o_1
X_32537_ _35929_/CLK _32537_/D VGND VGND VPWR VPWR _32537_/Q sky130_fd_sc_hd__dfxtp_1
X_35256_ _35320_/CLK _35256_/D VGND VGND VPWR VPWR _35256_/Q sky130_fd_sc_hd__dfxtp_1
X_23270_ _23270_/A VGND VGND VPWR VPWR _32162_/D sky130_fd_sc_hd__clkbuf_1
X_20482_ _18348_/X _20480_/X _20481_/X _18358_/X VGND VGND VPWR VPWR _20482_/X sky130_fd_sc_hd__a22o_1
XFILLER_197_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32468_ _36076_/CLK _32468_/D VGND VGND VPWR VPWR _32468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34207_ _36121_/CLK _34207_/D VGND VGND VPWR VPWR _34207_/Q sky130_fd_sc_hd__dfxtp_1
X_22221_ _22221_/A VGND VGND VPWR VPWR _36225_/D sky130_fd_sc_hd__clkbuf_1
X_31419_ _31551_/S VGND VGND VPWR VPWR _31438_/S sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_173_CLK clkbuf_6_28__f_CLK/X VGND VGND VPWR VPWR _34070_/CLK sky130_fd_sc_hd__clkbuf_16
X_35187_ _35187_/CLK _35187_/D VGND VGND VPWR VPWR _35187_/Q sky130_fd_sc_hd__dfxtp_1
X_32399_ _35983_/CLK _32399_/D VGND VGND VPWR VPWR _32399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22152_ _22505_/A VGND VGND VPWR VPWR _22152_/X sky130_fd_sc_hd__clkbuf_4
X_34138_ _36219_/CLK _34138_/D VGND VGND VPWR VPWR _34138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_218_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21103_ _22469_/A VGND VGND VPWR VPWR _21103_/X sky130_fd_sc_hd__buf_4
XFILLER_47_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34069_ _36181_/CLK _34069_/D VGND VGND VPWR VPWR _34069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22083_ _33918_/Q _33854_/Q _33790_/Q _36094_/Q _21977_/X _21978_/X VGND VGND VPWR
+ VPWR _22083_/X sky130_fd_sc_hd__mux4_1
X_26960_ _33907_/Q _23384_/X _26960_/S VGND VGND VPWR VPWR _26961_/A sky130_fd_sc_hd__mux2_1
XTAP_6829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25911_ _25911_/A VGND VGND VPWR VPWR _33412_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21034_ _22446_/A VGND VGND VPWR VPWR _21034_/X sky130_fd_sc_hd__clkbuf_4
X_26891_ _26891_/A VGND VGND VPWR VPWR _33874_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_248_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28630_ _27810_/X _34636_/Q _28640_/S VGND VGND VPWR VPWR _28631_/A sky130_fd_sc_hd__mux2_1
X_25842_ _25842_/A VGND VGND VPWR VPWR _33379_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_6_44__f_CLK clkbuf_5_22_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_44__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_59_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25773_ _24939_/X _33347_/Q _25781_/S VGND VGND VPWR VPWR _25774_/A sky130_fd_sc_hd__mux2_1
X_28561_ _27708_/X _34603_/Q _28577_/S VGND VGND VPWR VPWR _28562_/A sky130_fd_sc_hd__mux2_1
X_22985_ _22984_/X _32053_/Q _23009_/S VGND VGND VPWR VPWR _22986_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27512_ _34137_/Q _27044_/X _27524_/S VGND VGND VPWR VPWR _27513_/A sky130_fd_sc_hd__mux2_1
X_24724_ _24724_/A VGND VGND VPWR VPWR _32883_/D sky130_fd_sc_hd__clkbuf_1
X_28492_ _28492_/A VGND VGND VPWR VPWR _34570_/D sky130_fd_sc_hd__clkbuf_1
X_21936_ _34170_/Q _34106_/Q _34042_/Q _33978_/Q _21693_/X _21694_/X VGND VGND VPWR
+ VPWR _21936_/X sky130_fd_sc_hd__mux4_1
XFILLER_15_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27443_ _27443_/A VGND VGND VPWR VPWR _34104_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24655_ _23076_/X _32851_/Q _24659_/S VGND VGND VPWR VPWR _24656_/A sky130_fd_sc_hd__mux2_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21867_ _21867_/A _21867_/B _21867_/C _21867_/D VGND VGND VPWR VPWR _21868_/A sky130_fd_sc_hd__or4_1
XFILLER_243_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23606_ _22940_/X _32295_/Q _23610_/S VGND VGND VPWR VPWR _23607_/A sky130_fd_sc_hd__mux2_1
X_27374_ _27374_/A VGND VGND VPWR VPWR _34071_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_179_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20818_ _32602_/Q _32538_/Q _32474_/Q _35930_/Q _20817_/X _22317_/A VGND VGND VPWR
+ VPWR _20818_/X sky130_fd_sc_hd__mux4_1
XFILLER_169_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24586_ _22974_/X _32818_/Q _24588_/S VGND VGND VPWR VPWR _24587_/A sky130_fd_sc_hd__mux2_1
X_21798_ _21798_/A VGND VGND VPWR VPWR _36213_/D sky130_fd_sc_hd__buf_6
XFILLER_169_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26325_ _26325_/A VGND VGND VPWR VPWR _33608_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29113_ _29113_/A VGND VGND VPWR VPWR _34863_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23537_ _23537_/A VGND VGND VPWR VPWR _32263_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20749_ _33880_/Q _33816_/Q _33752_/Q _36056_/Q _20712_/X _20713_/X VGND VGND VPWR
+ VPWR _20749_/X sky130_fd_sc_hd__mux4_1
XFILLER_156_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29044_ _34831_/Q _27211_/X _29048_/S VGND VGND VPWR VPWR _29045_/A sky130_fd_sc_hd__mux2_1
X_26256_ _24855_/X _33576_/Q _26258_/S VGND VGND VPWR VPWR _26257_/A sky130_fd_sc_hd__mux2_1
X_23468_ _23468_/A VGND VGND VPWR VPWR _32234_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_221_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25207_ _33080_/Q _23402_/X _25217_/S VGND VGND VPWR VPWR _25208_/A sky130_fd_sc_hd__mux2_1
X_22419_ _22309_/X _22417_/X _22418_/X _22312_/X VGND VGND VPWR VPWR _22419_/X sky130_fd_sc_hd__a22o_1
X_26187_ _26187_/A VGND VGND VPWR VPWR _33543_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_164_CLK clkbuf_6_30__f_CLK/X VGND VGND VPWR VPWR _35664_/CLK sky130_fd_sc_hd__clkbuf_16
X_23399_ input27/X VGND VGND VPWR VPWR _23399_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_136_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25138_ _33047_/Q _23234_/X _25154_/S VGND VGND VPWR VPWR _25139_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17960_ _17960_/A VGND VGND VPWR VPWR _17960_/X sky130_fd_sc_hd__buf_4
X_29946_ _35228_/Q _29348_/X _29952_/S VGND VGND VPWR VPWR _29947_/A sky130_fd_sc_hd__mux2_1
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25069_ _25069_/A VGND VGND VPWR VPWR _33015_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16911_ _34925_/Q _34861_/Q _34797_/Q _34733_/Q _16807_/X _16808_/X VGND VGND VPWR
+ VPWR _16911_/X sky130_fd_sc_hd__mux4_1
XFILLER_77_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17891_ _17704_/X _17889_/X _17890_/X _17707_/X VGND VGND VPWR VPWR _17891_/X sky130_fd_sc_hd__a22o_1
XFILLER_120_730 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29877_ _29877_/A VGND VGND VPWR VPWR _35195_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19630_ _34937_/Q _34873_/Q _34809_/Q _34745_/Q _19460_/X _19461_/X VGND VGND VPWR
+ VPWR _19630_/X sky130_fd_sc_hd__mux4_1
XFILLER_238_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28828_ _28828_/A VGND VGND VPWR VPWR _34728_/D sky130_fd_sc_hd__clkbuf_1
X_16842_ _16805_/X _16840_/X _16841_/X _16810_/X VGND VGND VPWR VPWR _16842_/X sky130_fd_sc_hd__a22o_1
XFILLER_77_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19561_ _35191_/Q _35127_/Q _35063_/Q _32247_/Q _19310_/X _19311_/X VGND VGND VPWR
+ VPWR _19561_/X sky130_fd_sc_hd__mux4_1
XFILLER_92_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28759_ _28759_/A VGND VGND VPWR VPWR _34696_/D sky130_fd_sc_hd__clkbuf_1
X_16773_ _16493_/X _16771_/X _16772_/X _16498_/X VGND VGND VPWR VPWR _16773_/X sky130_fd_sc_hd__a22o_1
XFILLER_168_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18512_ _18440_/X _18510_/X _18511_/X _18445_/X VGND VGND VPWR VPWR _18512_/X sky130_fd_sc_hd__a22o_1
XFILLER_230_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31770_ _31770_/A VGND VGND VPWR VPWR _36092_/D sky130_fd_sc_hd__clkbuf_1
X_19492_ _19453_/X _19490_/X _19491_/X _19456_/X VGND VGND VPWR VPWR _19492_/X sky130_fd_sc_hd__a22o_1
XTAP_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18443_ _33624_/Q _33560_/Q _33496_/Q _33432_/Q _18441_/X _18442_/X VGND VGND VPWR
+ VPWR _18443_/X sky130_fd_sc_hd__mux4_1
X_30721_ _30721_/A VGND VGND VPWR VPWR _35595_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_1377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33440_ _36202_/CLK _33440_/D VGND VGND VPWR VPWR _33440_/Q sky130_fd_sc_hd__dfxtp_1
X_18374_ input81/X input82/X VGND VGND VPWR VPWR _20157_/A sky130_fd_sc_hd__or2_4
XFILLER_21_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30652_ _30652_/A VGND VGND VPWR VPWR _35562_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17325_ _17321_/X _17324_/X _17151_/X VGND VGND VPWR VPWR _17333_/C sky130_fd_sc_hd__o21ba_1
XFILLER_105_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30583_ _35530_/Q _29491_/X _30597_/S VGND VGND VPWR VPWR _30584_/A sky130_fd_sc_hd__mux2_1
X_33371_ _36059_/CLK _33371_/D VGND VGND VPWR VPWR _33371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35110_ _35625_/CLK _35110_/D VGND VGND VPWR VPWR _35110_/Q sky130_fd_sc_hd__dfxtp_1
X_32322_ _35970_/CLK _32322_/D VGND VGND VPWR VPWR _32322_/Q sky130_fd_sc_hd__dfxtp_1
X_36090_ _36090_/CLK _36090_/D VGND VGND VPWR VPWR _36090_/Q sky130_fd_sc_hd__dfxtp_1
X_17256_ _35447_/Q _35383_/Q _35319_/Q _35255_/Q _17254_/X _17255_/X VGND VGND VPWR
+ VPWR _17256_/X sky130_fd_sc_hd__mux4_1
XFILLER_128_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16207_ _16203_/X _16206_/X _16104_/X VGND VGND VPWR VPWR _16208_/D sky130_fd_sc_hd__o21ba_1
XFILLER_174_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35041_ _35168_/CLK _35041_/D VGND VGND VPWR VPWR _35041_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_155_CLK clkbuf_6_31__f_CLK/X VGND VGND VPWR VPWR _34963_/CLK sky130_fd_sc_hd__clkbuf_16
X_17187_ _33077_/Q _32053_/Q _35829_/Q _35765_/Q _17078_/X _17079_/X VGND VGND VPWR
+ VPWR _17187_/X sky130_fd_sc_hd__mux4_1
X_32253_ _35194_/CLK _32253_/D VGND VGND VPWR VPWR _32253_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16138_ _16138_/A _16138_/B _16138_/C _16138_/D VGND VGND VPWR VPWR _16139_/A sky130_fd_sc_hd__or4_2
X_31204_ _27723_/X _35824_/Q _31210_/S VGND VGND VPWR VPWR _31205_/A sky130_fd_sc_hd__mux2_1
X_32184_ _36002_/CLK _32184_/D VGND VGND VPWR VPWR _32184_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16069_ _17936_/A VGND VGND VPWR VPWR _16069_/X sky130_fd_sc_hd__buf_4
X_31135_ _35792_/Q input54/X _31137_/S VGND VGND VPWR VPWR _31136_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_1359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31066_ _35759_/Q input18/X _31074_/S VGND VGND VPWR VPWR _31067_/A sky130_fd_sc_hd__mux2_1
X_35943_ _35943_/CLK _35943_/D VGND VGND VPWR VPWR _35943_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30017_ _30065_/S VGND VGND VPWR VPWR _30036_/S sky130_fd_sc_hd__buf_6
X_19828_ _19824_/X _19827_/X _19785_/X VGND VGND VPWR VPWR _19850_/A sky130_fd_sc_hd__o21ba_1
XFILLER_69_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35874_ _35875_/CLK _35874_/D VGND VGND VPWR VPWR _35874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34825_ _34957_/CLK _34825_/D VGND VGND VPWR VPWR _34825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19759_ _19720_/X _19757_/X _19758_/X _19724_/X VGND VGND VPWR VPWR _19759_/X sky130_fd_sc_hd__a22o_1
XFILLER_42_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34756_ _34949_/CLK _34756_/D VGND VGND VPWR VPWR _34756_/Q sky130_fd_sc_hd__dfxtp_1
X_22770_ _32914_/Q _32850_/Q _32786_/Q _32722_/Q _20584_/X _20587_/X VGND VGND VPWR
+ VPWR _22770_/X sky130_fd_sc_hd__mux4_1
X_31968_ _34085_/CLK _31968_/D VGND VGND VPWR VPWR _31968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33707_ _34987_/CLK _33707_/D VGND VGND VPWR VPWR _33707_/Q sky130_fd_sc_hd__dfxtp_1
X_21721_ _21717_/X _21720_/X _21412_/X VGND VGND VPWR VPWR _21722_/D sky130_fd_sc_hd__o21ba_1
X_30919_ _30919_/A VGND VGND VPWR VPWR _35689_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34687_ _35071_/CLK _34687_/D VGND VGND VPWR VPWR _34687_/Q sky130_fd_sc_hd__dfxtp_1
X_31899_ _31899_/A VGND VGND VPWR VPWR _36153_/D sky130_fd_sc_hd__clkbuf_1
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24440_ _24440_/A VGND VGND VPWR VPWR _32748_/D sky130_fd_sc_hd__clkbuf_1
X_33638_ _34146_/CLK _33638_/D VGND VGND VPWR VPWR _33638_/Q sky130_fd_sc_hd__dfxtp_1
X_21652_ _33650_/Q _33586_/Q _33522_/Q _33458_/Q _21447_/X _21448_/X VGND VGND VPWR
+ VPWR _21652_/X sky130_fd_sc_hd__mux4_1
XFILLER_244_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20603_ _22400_/A VGND VGND VPWR VPWR _20603_/X sky130_fd_sc_hd__buf_4
X_24371_ _23055_/X _32716_/Q _24381_/S VGND VGND VPWR VPWR _24372_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21583_ _34160_/Q _34096_/Q _34032_/Q _33968_/Q _21340_/X _21341_/X VGND VGND VPWR
+ VPWR _21583_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_394_CLK clkbuf_6_40__f_CLK/X VGND VGND VPWR VPWR _35704_/CLK sky130_fd_sc_hd__clkbuf_16
X_33569_ _34593_/CLK _33569_/D VGND VGND VPWR VPWR _33569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26110_ _26110_/A VGND VGND VPWR VPWR _33506_/D sky130_fd_sc_hd__clkbuf_1
X_23322_ _23322_/A VGND VGND VPWR VPWR _32178_/D sky130_fd_sc_hd__clkbuf_1
X_35308_ _35691_/CLK _35308_/D VGND VGND VPWR VPWR _35308_/Q sky130_fd_sc_hd__dfxtp_1
X_20534_ _35668_/Q _35028_/Q _34388_/Q _33748_/Q _18412_/X _18413_/X VGND VGND VPWR
+ VPWR _20534_/X sky130_fd_sc_hd__mux4_1
X_27090_ input10/X VGND VGND VPWR VPWR _27090_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_137_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26041_ _24936_/X _33474_/Q _26051_/S VGND VGND VPWR VPWR _26042_/A sky130_fd_sc_hd__mux2_1
X_23253_ _32157_/Q _23252_/X _23259_/S VGND VGND VPWR VPWR _23254_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35239_ _35367_/CLK _35239_/D VGND VGND VPWR VPWR _35239_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_146_CLK clkbuf_6_29__f_CLK/X VGND VGND VPWR VPWR _33941_/CLK sky130_fd_sc_hd__clkbuf_16
X_20465_ _20461_/X _20464_/X _20138_/A VGND VGND VPWR VPWR _20487_/A sky130_fd_sc_hd__o21ba_1
XFILLER_180_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22204_ _35713_/Q _32223_/Q _35585_/Q _35521_/Q _21917_/X _21918_/X VGND VGND VPWR
+ VPWR _22204_/X sky130_fd_sc_hd__mux4_1
XFILLER_106_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23184_ _23024_/X _32130_/Q _23194_/S VGND VGND VPWR VPWR _23185_/A sky130_fd_sc_hd__mux2_1
X_20396_ _20392_/X _20395_/X _20171_/X VGND VGND VPWR VPWR _20397_/D sky130_fd_sc_hd__o21ba_1
X_29800_ _29800_/A VGND VGND VPWR VPWR _35158_/D sky130_fd_sc_hd__clkbuf_1
X_22135_ _22131_/X _22134_/X _22093_/X _22094_/X VGND VGND VPWR VPWR _22150_/B sky130_fd_sc_hd__o211a_1
XTAP_6604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27992_ _27992_/A VGND VGND VPWR VPWR _34333_/D sky130_fd_sc_hd__clkbuf_1
Xoutput260 _32454_/Q VGND VGND VPWR VPWR D3[48] sky130_fd_sc_hd__buf_2
XTAP_6626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput271 _32464_/Q VGND VGND VPWR VPWR D3[58] sky130_fd_sc_hd__buf_2
XTAP_6637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29731_ _35126_/Q _29429_/X _29745_/S VGND VGND VPWR VPWR _29732_/A sky130_fd_sc_hd__mux2_1
X_26943_ _26943_/A VGND VGND VPWR VPWR _33898_/D sky130_fd_sc_hd__clkbuf_1
X_22066_ _21956_/X _22064_/X _22065_/X _21959_/X VGND VGND VPWR VPWR _22066_/X sky130_fd_sc_hd__a22o_1
XTAP_6659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21017_ _21017_/A VGND VGND VPWR VPWR _36191_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_212_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29662_ _29797_/A _29662_/B VGND VGND VPWR VPWR _29795_/S sky130_fd_sc_hd__nor2_8
XFILLER_87_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26874_ _33866_/Q _23463_/X _26888_/S VGND VGND VPWR VPWR _26875_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28613_ _27785_/X _34628_/Q _28619_/S VGND VGND VPWR VPWR _28614_/A sky130_fd_sc_hd__mux2_1
XFILLER_235_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25825_ _25825_/A VGND VGND VPWR VPWR _33371_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29593_ _29593_/A VGND VGND VPWR VPWR _35060_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_216_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25756_ _24914_/X _33339_/Q _25760_/S VGND VGND VPWR VPWR _25757_/A sky130_fd_sc_hd__mux2_1
X_28544_ _27683_/X _34595_/Q _28556_/S VGND VGND VPWR VPWR _28545_/A sky130_fd_sc_hd__mux2_1
X_22968_ input19/X VGND VGND VPWR VPWR _22968_/X sky130_fd_sc_hd__buf_2
XFILLER_231_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21919_ _35705_/Q _32214_/Q _35577_/Q _35513_/Q _21917_/X _21918_/X VGND VGND VPWR
+ VPWR _21919_/X sky130_fd_sc_hd__mux4_2
X_24707_ _22953_/X _32875_/Q _24723_/S VGND VGND VPWR VPWR _24708_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28475_ _28475_/A VGND VGND VPWR VPWR _34562_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25687_ _24812_/X _33306_/Q _25697_/S VGND VGND VPWR VPWR _25688_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22899_ _22899_/A VGND VGND VPWR VPWR _32025_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24638_ _24638_/A VGND VGND VPWR VPWR _32842_/D sky130_fd_sc_hd__clkbuf_1
X_27426_ _27426_/A VGND VGND VPWR VPWR _34096_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1069 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27357_ _34064_/Q _27214_/X _27359_/S VGND VGND VPWR VPWR _27358_/A sky130_fd_sc_hd__mux2_1
XFILLER_208_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24569_ _24659_/S VGND VGND VPWR VPWR _24588_/S sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_385_CLK clkbuf_6_42__f_CLK/X VGND VGND VPWR VPWR _33913_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_12_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17110_ _16998_/X _17108_/X _17109_/X _17001_/X VGND VGND VPWR VPWR _17110_/X sky130_fd_sc_hd__a22o_1
X_26308_ _26308_/A VGND VGND VPWR VPWR _33600_/D sky130_fd_sc_hd__clkbuf_1
X_18090_ _34703_/Q _34639_/Q _34575_/Q _34511_/Q _17998_/X _17999_/X VGND VGND VPWR
+ VPWR _18090_/X sky130_fd_sc_hd__mux4_1
XFILLER_168_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27288_ _34031_/Q _27112_/X _27296_/S VGND VGND VPWR VPWR _27289_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17041_ _17003_/X _17039_/X _17040_/X _17006_/X VGND VGND VPWR VPWR _17041_/X sky130_fd_sc_hd__a22o_1
XFILLER_239_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29027_ _34823_/Q _27186_/X _29027_/S VGND VGND VPWR VPWR _29028_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26239_ _26350_/S VGND VGND VPWR VPWR _26258_/S sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_137_CLK clkbuf_6_23__f_CLK/X VGND VGND VPWR VPWR _35800_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_139_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18992_ _18747_/X _18990_/X _18991_/X _18750_/X VGND VGND VPWR VPWR _18992_/X sky130_fd_sc_hd__a22o_1
XFILLER_3_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17943_ _33675_/Q _33611_/Q _33547_/Q _33483_/Q _17906_/X _17907_/X VGND VGND VPWR
+ VPWR _17943_/X sky130_fd_sc_hd__mux4_1
X_29929_ _29929_/A VGND VGND VPWR VPWR _35220_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32940_ _36141_/CLK _32940_/D VGND VGND VPWR VPWR _32940_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17874_ _17874_/A VGND VGND VPWR VPWR _32008_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_78_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19613_ _32121_/Q _32313_/Q _32377_/Q _35897_/Q _19580_/X _19368_/X VGND VGND VPWR
+ VPWR _19613_/X sky130_fd_sc_hd__mux4_1
XFILLER_226_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16825_ _16706_/X _16823_/X _16824_/X _16712_/X VGND VGND VPWR VPWR _16825_/X sky130_fd_sc_hd__a22o_1
X_32871_ _32871_/CLK _32871_/D VGND VGND VPWR VPWR _32871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34610_ _35377_/CLK _34610_/D VGND VGND VPWR VPWR _34610_/Q sky130_fd_sc_hd__dfxtp_1
X_31822_ _31822_/A VGND VGND VPWR VPWR _36117_/D sky130_fd_sc_hd__clkbuf_1
X_19544_ _32631_/Q _32567_/Q _32503_/Q _35959_/Q _19223_/X _19360_/X VGND VGND VPWR
+ VPWR _19544_/X sky130_fd_sc_hd__mux4_1
XFILLER_93_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35590_ _35721_/CLK _35590_/D VGND VGND VPWR VPWR _35590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16756_ _35625_/Q _34985_/Q _34345_/Q _33705_/Q _16438_/X _16439_/X VGND VGND VPWR
+ VPWR _16756_/X sky130_fd_sc_hd__mux4_1
XFILLER_111_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34541_ _36140_/CLK _34541_/D VGND VGND VPWR VPWR _34541_/Q sky130_fd_sc_hd__dfxtp_1
X_19475_ _19471_/X _19474_/X _19432_/X VGND VGND VPWR VPWR _19497_/A sky130_fd_sc_hd__o21ba_1
X_31753_ _36084_/Q input24/X _31771_/S VGND VGND VPWR VPWR _31754_/A sky130_fd_sc_hd__mux2_1
XFILLER_222_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16687_ _33063_/Q _32039_/Q _35815_/Q _35751_/Q _16372_/X _16373_/X VGND VGND VPWR
+ VPWR _16687_/X sky130_fd_sc_hd__mux4_1
XFILLER_185_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18426_ _18348_/X _18424_/X _18425_/X _18358_/X VGND VGND VPWR VPWR _18426_/X sky130_fd_sc_hd__a22o_1
X_30704_ _30704_/A VGND VGND VPWR VPWR _35587_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34472_ _36137_/CLK _34472_/D VGND VGND VPWR VPWR _34472_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31684_ _27834_/X _36052_/Q _31686_/S VGND VGND VPWR VPWR _31685_/A sky130_fd_sc_hd__mux2_1
X_36211_ _36211_/CLK _36211_/D VGND VGND VPWR VPWR _36211_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33423_ _33425_/CLK _33423_/D VGND VGND VPWR VPWR _33423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18357_ _20071_/A VGND VGND VPWR VPWR _20162_/A sky130_fd_sc_hd__buf_12
X_30635_ _30635_/A VGND VGND VPWR VPWR _35554_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_376_CLK clkbuf_6_42__f_CLK/X VGND VGND VPWR VPWR _35449_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_124_1445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17308_ _17206_/X _17306_/X _17307_/X _17209_/X VGND VGND VPWR VPWR _17308_/X sky130_fd_sc_hd__a22o_1
X_36142_ _36142_/CLK _36142_/D VGND VGND VPWR VPWR _36142_/Q sky130_fd_sc_hd__dfxtp_1
X_33354_ _33673_/CLK _33354_/D VGND VGND VPWR VPWR _33354_/Q sky130_fd_sc_hd__dfxtp_1
X_18288_ _33622_/Q _33558_/Q _33494_/Q _33430_/Q _18284_/X _18287_/X VGND VGND VPWR
+ VPWR _18288_/X sky130_fd_sc_hd__mux4_1
X_30566_ _35522_/Q _29466_/X _30576_/S VGND VGND VPWR VPWR _30567_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_6_8__f_CLK clkbuf_5_4_0_CLK/X VGND VGND VPWR VPWR _35560_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_119_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32305_ _35953_/CLK _32305_/D VGND VGND VPWR VPWR _32305_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_128_CLK clkbuf_6_21__f_CLK/X VGND VGND VPWR VPWR _36121_/CLK sky130_fd_sc_hd__clkbuf_16
X_17239_ _17199_/X _17237_/X _17238_/X _17204_/X VGND VGND VPWR VPWR _17239_/X sky130_fd_sc_hd__a22o_1
X_36073_ _36073_/CLK _36073_/D VGND VGND VPWR VPWR _36073_/Q sky130_fd_sc_hd__dfxtp_1
X_33285_ _33415_/CLK _33285_/D VGND VGND VPWR VPWR _33285_/Q sky130_fd_sc_hd__dfxtp_1
X_30497_ _35489_/Q _29364_/X _30513_/S VGND VGND VPWR VPWR _30498_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35024_ _35731_/CLK _35024_/D VGND VGND VPWR VPWR _35024_/Q sky130_fd_sc_hd__dfxtp_1
X_32236_ _35661_/CLK _32236_/D VGND VGND VPWR VPWR _32236_/Q sky130_fd_sc_hd__dfxtp_1
X_20250_ _32651_/Q _32587_/Q _32523_/Q _35979_/Q _19929_/X _20066_/X VGND VGND VPWR
+ VPWR _20250_/X sky130_fd_sc_hd__mux4_1
XFILLER_143_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20181_ _20177_/X _20180_/X _20138_/X VGND VGND VPWR VPWR _20203_/A sky130_fd_sc_hd__o21ba_2
XFILLER_118_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32167_ _35367_/CLK _32167_/D VGND VGND VPWR VPWR _32167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31118_ _31145_/S VGND VGND VPWR VPWR _31137_/S sky130_fd_sc_hd__buf_4
XFILLER_157_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32098_ _32356_/CLK _32098_/D VGND VGND VPWR VPWR _32098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_233_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23940_ _23027_/X _32515_/Q _23948_/S VGND VGND VPWR VPWR _23941_/A sky130_fd_sc_hd__mux2_1
X_35926_ _35990_/CLK _35926_/D VGND VGND VPWR VPWR _35926_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_300_CLK clkbuf_6_57__f_CLK/X VGND VGND VPWR VPWR _35843_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31049_ _35751_/Q input9/X _31053_/S VGND VGND VPWR VPWR _31050_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35857_ _35857_/CLK _35857_/D VGND VGND VPWR VPWR _35857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23871_ _22925_/X _32482_/Q _23885_/S VGND VGND VPWR VPWR _23872_/A sky130_fd_sc_hd__mux2_1
X_25610_ _25610_/A VGND VGND VPWR VPWR _33269_/D sky130_fd_sc_hd__clkbuf_1
X_22822_ _33428_/Q _33364_/Q _33300_/Q _33236_/Q _20637_/X _20639_/X VGND VGND VPWR
+ VPWR _22822_/X sky130_fd_sc_hd__mux4_1
XFILLER_211_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34808_ _35833_/CLK _34808_/D VGND VGND VPWR VPWR _34808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26590_ _26590_/A VGND VGND VPWR VPWR _33733_/D sky130_fd_sc_hd__clkbuf_1
X_35788_ _35852_/CLK _35788_/D VGND VGND VPWR VPWR _35788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25541_ _25541_/A VGND VGND VPWR VPWR _33237_/D sky130_fd_sc_hd__clkbuf_1
X_22753_ _34449_/Q _36177_/Q _34321_/Q _34257_/Q _22535_/X _22536_/X VGND VGND VPWR
+ VPWR _22753_/X sky130_fd_sc_hd__mux4_1
XFILLER_164_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34739_ _34927_/CLK _34739_/D VGND VGND VPWR VPWR _34739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28260_ _28260_/A VGND VGND VPWR VPWR _34460_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21704_ _32115_/Q _32307_/Q _32371_/Q _35891_/Q _21527_/X _21668_/X VGND VGND VPWR
+ VPWR _21704_/X sky130_fd_sc_hd__mux4_1
XFILLER_241_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25472_ _24892_/X _33204_/Q _25490_/S VGND VGND VPWR VPWR _25473_/A sky130_fd_sc_hd__mux2_1
XFILLER_198_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22684_ _35663_/Q _35023_/Q _34383_/Q _33743_/Q _22450_/X _22451_/X VGND VGND VPWR
+ VPWR _22684_/X sky130_fd_sc_hd__mux4_1
XFILLER_53_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27211_ input53/X VGND VGND VPWR VPWR _27211_/X sky130_fd_sc_hd__buf_4
XFILLER_209_1380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24423_ _24423_/A VGND VGND VPWR VPWR _32740_/D sky130_fd_sc_hd__clkbuf_1
X_28191_ _27760_/X _34428_/Q _28193_/S VGND VGND VPWR VPWR _28192_/A sky130_fd_sc_hd__mux2_1
X_21635_ _21631_/X _21634_/X _21387_/X _21388_/X VGND VGND VPWR VPWR _21650_/B sky130_fd_sc_hd__o211a_1
XFILLER_233_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_367_CLK clkbuf_6_43__f_CLK/X VGND VGND VPWR VPWR _36152_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_90_1466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27142_ _27142_/A VGND VGND VPWR VPWR _33976_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_205_1266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24354_ _23030_/X _32708_/Q _24360_/S VGND VGND VPWR VPWR _24355_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21566_ _35695_/Q _32203_/Q _35567_/Q _35503_/Q _21564_/X _21565_/X VGND VGND VPWR
+ VPWR _21566_/X sky130_fd_sc_hd__mux4_1
X_23305_ input17/X VGND VGND VPWR VPWR _23305_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_119_CLK clkbuf_6_21__f_CLK/X VGND VGND VPWR VPWR _34654_/CLK sky130_fd_sc_hd__clkbuf_16
X_20517_ _20517_/A _20517_/B _20517_/C _20517_/D VGND VGND VPWR VPWR _20518_/A sky130_fd_sc_hd__or4_1
X_27073_ _33954_/Q _27072_/X _27094_/S VGND VGND VPWR VPWR _27074_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24285_ _22928_/X _32675_/Q _24297_/S VGND VGND VPWR VPWR _24286_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21497_ _21493_/X _21496_/X _21387_/X _21388_/X VGND VGND VPWR VPWR _21514_/B sky130_fd_sc_hd__o211a_1
XFILLER_14_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26024_ _24911_/X _33466_/Q _26030_/S VGND VGND VPWR VPWR _26025_/A sky130_fd_sc_hd__mux2_1
X_23236_ _23236_/A VGND VGND VPWR VPWR _32151_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_238_1020 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20448_ _18301_/X _20446_/X _20447_/X _18307_/X VGND VGND VPWR VPWR _20448_/X sky130_fd_sc_hd__a22o_1
XFILLER_153_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1053 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23167_ _22999_/X _32122_/Q _23173_/S VGND VGND VPWR VPWR _23168_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20379_ _32143_/Q _32335_/Q _32399_/Q _35919_/Q _20286_/X _20074_/X VGND VGND VPWR
+ VPWR _20379_/X sky130_fd_sc_hd__mux4_1
XFILLER_106_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22118_ _22471_/A VGND VGND VPWR VPWR _22118_/X sky130_fd_sc_hd__buf_2
XFILLER_171_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23098_ _22897_/X _32089_/Q _23110_/S VGND VGND VPWR VPWR _23099_/A sky130_fd_sc_hd__mux2_1
X_27975_ _31147_/A _30607_/B VGND VGND VPWR VPWR _28108_/S sky130_fd_sc_hd__nor2_8
XFILLER_122_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29714_ _35118_/Q _29404_/X _29724_/S VGND VGND VPWR VPWR _29715_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26926_ _26926_/A VGND VGND VPWR VPWR _33890_/D sky130_fd_sc_hd__clkbuf_1
X_22049_ _21799_/X _22045_/X _22048_/X _21804_/X VGND VGND VPWR VPWR _22049_/X sky130_fd_sc_hd__a22o_1
XFILLER_85_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_929 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29645_ _29645_/A VGND VGND VPWR VPWR _35085_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26857_ _33858_/Q _23435_/X _26867_/S VGND VGND VPWR VPWR _26858_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16610_ _16606_/X _16609_/X _16434_/X _16435_/X VGND VGND VPWR VPWR _16627_/B sky130_fd_sc_hd__o211a_1
X_25808_ _24991_/X _33364_/Q _25810_/S VGND VGND VPWR VPWR _25809_/A sky130_fd_sc_hd__mux2_1
X_17590_ _33665_/Q _33601_/Q _33537_/Q _33473_/Q _17553_/X _17554_/X VGND VGND VPWR
+ VPWR _17590_/X sky130_fd_sc_hd__mux4_1
X_29576_ _29576_/A VGND VGND VPWR VPWR _35052_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26788_ _33825_/Q _23265_/X _26804_/S VGND VGND VPWR VPWR _26789_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28527_ _27658_/X _34587_/Q _28535_/S VGND VGND VPWR VPWR _28528_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16541_ _32099_/Q _32291_/Q _32355_/Q _35875_/Q _16221_/X _16362_/X VGND VGND VPWR
+ VPWR _16541_/X sky130_fd_sc_hd__mux4_1
XFILLER_141_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25739_ _24889_/X _33331_/Q _25739_/S VGND VGND VPWR VPWR _25740_/A sky130_fd_sc_hd__mux2_1
XFILLER_203_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_1388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19260_ _32111_/Q _32303_/Q _32367_/Q _35887_/Q _19227_/X _19015_/X VGND VGND VPWR
+ VPWR _19260_/X sky130_fd_sc_hd__mux4_1
XFILLER_232_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16472_ _16353_/X _16470_/X _16471_/X _16359_/X VGND VGND VPWR VPWR _16472_/X sky130_fd_sc_hd__a22o_1
X_28458_ _28458_/A VGND VGND VPWR VPWR _34554_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18211_ _35219_/Q _35155_/Q _35091_/Q _32275_/Q _16092_/X _16094_/X VGND VGND VPWR
+ VPWR _18211_/X sky130_fd_sc_hd__mux4_1
XFILLER_70_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27409_ _27409_/A VGND VGND VPWR VPWR _34088_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_358_CLK clkbuf_6_46__f_CLK/X VGND VGND VPWR VPWR _35197_/CLK sky130_fd_sc_hd__clkbuf_16
X_19191_ _32621_/Q _32557_/Q _32493_/Q _35949_/Q _18870_/X _19007_/X VGND VGND VPWR
+ VPWR _19191_/X sky130_fd_sc_hd__mux4_1
X_28389_ _28389_/A VGND VGND VPWR VPWR _34521_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18142_ _18138_/X _18141_/X _17846_/X _17847_/X VGND VGND VPWR VPWR _18157_/B sky130_fd_sc_hd__o211a_1
XFILLER_12_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30420_ _35453_/Q _29450_/X _30420_/S VGND VGND VPWR VPWR _30421_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18073_ _33935_/Q _33871_/Q _33807_/Q _36111_/Q _16062_/X _16064_/X VGND VGND VPWR
+ VPWR _18073_/X sky130_fd_sc_hd__mux4_1
X_30351_ _35420_/Q _29348_/X _30357_/S VGND VGND VPWR VPWR _30352_/A sky130_fd_sc_hd__mux2_1
X_17024_ _17850_/A VGND VGND VPWR VPWR _17024_/X sky130_fd_sc_hd__buf_4
X_33070_ _35822_/CLK _33070_/D VGND VGND VPWR VPWR _33070_/Q sky130_fd_sc_hd__dfxtp_1
X_30282_ _30282_/A VGND VGND VPWR VPWR _35387_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32021_ _36191_/CLK _32021_/D VGND VGND VPWR VPWR _32021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18975_ _18969_/X _18974_/X _18726_/X VGND VGND VPWR VPWR _18997_/A sky130_fd_sc_hd__o21ba_1
XFILLER_234_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17926_ _35658_/Q _35018_/Q _34378_/Q _33738_/Q _17850_/X _17851_/X VGND VGND VPWR
+ VPWR _17926_/X sky130_fd_sc_hd__mux4_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33972_ _34101_/CLK _33972_/D VGND VGND VPWR VPWR _33972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35711_ _35711_/CLK _35711_/D VGND VGND VPWR VPWR _35711_/Q sky130_fd_sc_hd__dfxtp_1
X_32923_ _35997_/CLK _32923_/D VGND VGND VPWR VPWR _32923_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17857_ _17857_/A VGND VGND VPWR VPWR _17857_/X sky130_fd_sc_hd__buf_2
XFILLER_226_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16808_ _17161_/A VGND VGND VPWR VPWR _16808_/X sky130_fd_sc_hd__clkbuf_4
X_35642_ _35645_/CLK _35642_/D VGND VGND VPWR VPWR _35642_/Q sky130_fd_sc_hd__dfxtp_1
X_32854_ _36117_/CLK _32854_/D VGND VGND VPWR VPWR _32854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17788_ _17782_/X _17787_/X _17504_/X VGND VGND VPWR VPWR _17796_/C sky130_fd_sc_hd__o21ba_1
XFILLER_226_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31805_ _36109_/Q input51/X _31813_/S VGND VGND VPWR VPWR _31806_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19527_ _35190_/Q _35126_/Q _35062_/Q _32246_/Q _19310_/X _19311_/X VGND VGND VPWR
+ VPWR _19527_/X sky130_fd_sc_hd__mux4_1
X_35573_ _35701_/CLK _35573_/D VGND VGND VPWR VPWR _35573_/Q sky130_fd_sc_hd__dfxtp_1
X_16739_ _33641_/Q _33577_/Q _33513_/Q _33449_/Q _16494_/X _16495_/X VGND VGND VPWR
+ VPWR _16739_/X sky130_fd_sc_hd__mux4_1
XFILLER_53_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32785_ _32913_/CLK _32785_/D VGND VGND VPWR VPWR _32785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34524_ _36229_/CLK _34524_/D VGND VGND VPWR VPWR _34524_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31736_ _36076_/Q input15/X _31750_/S VGND VGND VPWR VPWR _31737_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19458_ _19458_/A VGND VGND VPWR VPWR _19458_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_224_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18409_ _34135_/Q _34071_/Q _34007_/Q _33943_/Q _18309_/X _18311_/X VGND VGND VPWR
+ VPWR _18409_/X sky130_fd_sc_hd__mux4_1
X_34455_ _34647_/CLK _34455_/D VGND VGND VPWR VPWR _34455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_349_CLK clkbuf_6_47__f_CLK/X VGND VGND VPWR VPWR _34174_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_50_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31667_ _31667_/A VGND VGND VPWR VPWR _36043_/D sky130_fd_sc_hd__clkbuf_1
X_19389_ _19385_/X _19388_/X _19112_/X VGND VGND VPWR VPWR _19390_/D sky130_fd_sc_hd__o21ba_1
X_33406_ _35648_/CLK _33406_/D VGND VGND VPWR VPWR _33406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21420_ _33899_/Q _33835_/Q _33771_/Q _36075_/Q _21271_/X _21272_/X VGND VGND VPWR
+ VPWR _21420_/X sky130_fd_sc_hd__mux4_1
X_30618_ _30618_/A VGND VGND VPWR VPWR _35546_/D sky130_fd_sc_hd__clkbuf_1
X_34386_ _35730_/CLK _34386_/D VGND VGND VPWR VPWR _34386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31598_ _31598_/A VGND VGND VPWR VPWR _36010_/D sky130_fd_sc_hd__clkbuf_1
X_36125_ _36125_/CLK _36125_/D VGND VGND VPWR VPWR _36125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33337_ _33914_/CLK _33337_/D VGND VGND VPWR VPWR _33337_/Q sky130_fd_sc_hd__dfxtp_1
X_21351_ _32105_/Q _32297_/Q _32361_/Q _35881_/Q _21174_/X _21315_/X VGND VGND VPWR
+ VPWR _21351_/X sky130_fd_sc_hd__mux4_1
XFILLER_108_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30549_ _35514_/Q _29441_/X _30555_/S VGND VGND VPWR VPWR _30550_/A sky130_fd_sc_hd__mux2_1
X_20302_ _20159_/X _20300_/X _20301_/X _20162_/X VGND VGND VPWR VPWR _20302_/X sky130_fd_sc_hd__a22o_1
XFILLER_198_1387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36056_ _36057_/CLK _36056_/D VGND VGND VPWR VPWR _36056_/Q sky130_fd_sc_hd__dfxtp_1
X_24070_ _23018_/X _32576_/Q _24084_/S VGND VGND VPWR VPWR _24071_/A sky130_fd_sc_hd__mux2_1
XFILLER_239_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33268_ _34100_/CLK _33268_/D VGND VGND VPWR VPWR _33268_/Q sky130_fd_sc_hd__dfxtp_1
X_21282_ _21278_/X _21281_/X _21034_/X _21035_/X VGND VGND VPWR VPWR _21297_/B sky130_fd_sc_hd__o211a_1
XFILLER_190_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35007_ _36096_/CLK _35007_/D VGND VGND VPWR VPWR _35007_/Q sky130_fd_sc_hd__dfxtp_1
X_23021_ input38/X VGND VGND VPWR VPWR _23021_/X sky130_fd_sc_hd__buf_2
X_20233_ _35210_/Q _35146_/Q _35082_/Q _32266_/Q _20016_/X _20017_/X VGND VGND VPWR
+ VPWR _20233_/X sky130_fd_sc_hd__mux4_1
X_32219_ _35713_/CLK _32219_/D VGND VGND VPWR VPWR _32219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33199_ _36079_/CLK _33199_/D VGND VGND VPWR VPWR _33199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20164_ _20164_/A VGND VGND VPWR VPWR _20164_/X sky130_fd_sc_hd__clkbuf_4
XTAP_5007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27760_ input32/X VGND VGND VPWR VPWR _27760_/X sky130_fd_sc_hd__clkbuf_4
X_20095_ _20091_/X _20094_/X _19818_/X VGND VGND VPWR VPWR _20096_/D sky130_fd_sc_hd__o21ba_1
XFILLER_170_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24972_ _24972_/A VGND VGND VPWR VPWR _32973_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26711_ _33789_/Q _23417_/X _26711_/S VGND VGND VPWR VPWR _26712_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35909_ _35973_/CLK _35909_/D VGND VGND VPWR VPWR _35909_/Q sky130_fd_sc_hd__dfxtp_1
X_23923_ _23002_/X _32507_/Q _23927_/S VGND VGND VPWR VPWR _23924_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27691_ _27691_/A VGND VGND VPWR VPWR _34213_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29430_ _34998_/Q _29429_/X _29451_/S VGND VGND VPWR VPWR _29431_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23854_ _22900_/X _32474_/Q _23864_/S VGND VGND VPWR VPWR _23855_/A sky130_fd_sc_hd__mux2_1
X_26642_ _33756_/Q _23249_/X _26648_/S VGND VGND VPWR VPWR _26643_/A sky130_fd_sc_hd__mux2_1
XFILLER_57_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22805_ _20581_/X _22803_/X _22804_/X _20591_/X VGND VGND VPWR VPWR _22805_/X sky130_fd_sc_hd__a22o_1
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29361_ _29525_/S VGND VGND VPWR VPWR _29389_/S sky130_fd_sc_hd__buf_4
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26573_ _26573_/A VGND VGND VPWR VPWR _33725_/D sky130_fd_sc_hd__clkbuf_1
X_23785_ _23785_/A VGND VGND VPWR VPWR _32378_/D sky130_fd_sc_hd__clkbuf_1
X_20997_ _20953_/X _20995_/X _20996_/X _20959_/X VGND VGND VPWR VPWR _20997_/X sky130_fd_sc_hd__a22o_1
XFILLER_26_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28312_ _27739_/X _34485_/Q _28328_/S VGND VGND VPWR VPWR _28313_/A sky130_fd_sc_hd__mux2_1
X_25524_ _24970_/X _33229_/Q _25532_/S VGND VGND VPWR VPWR _25525_/A sky130_fd_sc_hd__mux2_1
X_22736_ _32657_/Q _32593_/Q _32529_/Q _35985_/Q _22582_/X _21477_/A VGND VGND VPWR
+ VPWR _22736_/X sky130_fd_sc_hd__mux4_1
XFILLER_129_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29292_ _29292_/A VGND VGND VPWR VPWR _34948_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28243_ _27837_/X _34453_/Q _28243_/S VGND VGND VPWR VPWR _28244_/A sky130_fd_sc_hd__mux2_1
X_25455_ _24868_/X _33196_/Q _25469_/S VGND VGND VPWR VPWR _25456_/A sky130_fd_sc_hd__mux2_1
X_22667_ _22667_/A _22667_/B _22667_/C _22667_/D VGND VGND VPWR VPWR _22668_/A sky130_fd_sc_hd__or4_4
XFILLER_16_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24406_ _24406_/A VGND VGND VPWR VPWR _32732_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21618_ _21618_/A _21618_/B _21618_/C _21618_/D VGND VGND VPWR VPWR _21619_/A sky130_fd_sc_hd__or4_4
X_25386_ _25386_/A VGND VGND VPWR VPWR _33164_/D sky130_fd_sc_hd__clkbuf_1
X_28174_ _28243_/S VGND VGND VPWR VPWR _28193_/S sky130_fd_sc_hd__buf_4
XFILLER_90_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22598_ _22598_/A VGND VGND VPWR VPWR _22598_/X sky130_fd_sc_hd__buf_6
XFILLER_166_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24337_ _23005_/X _32700_/Q _24339_/S VGND VGND VPWR VPWR _24338_/A sky130_fd_sc_hd__mux2_1
X_27125_ _33971_/Q _27124_/X _27125_/S VGND VGND VPWR VPWR _27126_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_1389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21549_ _21549_/A VGND VGND VPWR VPWR _36206_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27056_ input62/X VGND VGND VPWR VPWR _27056_/X sky130_fd_sc_hd__buf_4
X_24268_ _22903_/X _32667_/Q _24276_/S VGND VGND VPWR VPWR _24269_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26007_ _24886_/X _33458_/Q _26009_/S VGND VGND VPWR VPWR _26008_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23219_ _23076_/X _32147_/Q _23223_/S VGND VGND VPWR VPWR _23220_/A sky130_fd_sc_hd__mux2_1
XFILLER_135_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24199_ _32636_/Q _23414_/X _24201_/S VGND VGND VPWR VPWR _24200_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1048 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18760_ _18751_/X _18758_/X _18759_/X VGND VGND VPWR VPWR _18761_/D sky130_fd_sc_hd__o21ba_1
X_27958_ _27958_/A VGND VGND VPWR VPWR _34317_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_923 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17711_ _33092_/Q _32068_/Q _35844_/Q _35780_/Q _17431_/X _17432_/X VGND VGND VPWR
+ VPWR _17711_/X sky130_fd_sc_hd__mux4_1
XFILLER_209_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26909_ _26909_/A VGND VGND VPWR VPWR _33882_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18691_ _33375_/Q _33311_/Q _33247_/Q _33183_/Q _18302_/X _18303_/X VGND VGND VPWR
+ VPWR _18691_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_5_18_0_CLK clkbuf_2_2_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_18_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_222_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27889_ _27889_/A VGND VGND VPWR VPWR _34284_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29628_ _29628_/A VGND VGND VPWR VPWR _35077_/D sky130_fd_sc_hd__clkbuf_1
X_17642_ _33090_/Q _32066_/Q _35842_/Q _35778_/Q _17431_/X _17432_/X VGND VGND VPWR
+ VPWR _17642_/X sky130_fd_sc_hd__mux4_1
XTAP_4873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17573_ _35648_/Q _35008_/Q _34368_/Q _33728_/Q _17497_/X _17498_/X VGND VGND VPWR
+ VPWR _17573_/X sky130_fd_sc_hd__mux4_1
X_29559_ _29559_/A VGND VGND VPWR VPWR _35044_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19312_ _35184_/Q _35120_/Q _35056_/Q _32187_/Q _19310_/X _19311_/X VGND VGND VPWR
+ VPWR _19312_/X sky130_fd_sc_hd__mux4_1
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16524_ _16877_/A VGND VGND VPWR VPWR _16524_/X sky130_fd_sc_hd__buf_4
XFILLER_16_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32570_ _35962_/CLK _32570_/D VGND VGND VPWR VPWR _32570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31521_ _31521_/A VGND VGND VPWR VPWR _35974_/D sky130_fd_sc_hd__clkbuf_1
X_19243_ _19100_/X _19241_/X _19242_/X _19103_/X VGND VGND VPWR VPWR _19243_/X sky130_fd_sc_hd__a22o_1
X_16455_ _17161_/A VGND VGND VPWR VPWR _16455_/X sky130_fd_sc_hd__clkbuf_4
X_34240_ _34815_/CLK _34240_/D VGND VGND VPWR VPWR _34240_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19174_ _35180_/Q _35116_/Q _35052_/Q _32172_/Q _18957_/X _18958_/X VGND VGND VPWR
+ VPWR _19174_/X sky130_fd_sc_hd__mux4_1
X_31452_ _31452_/A VGND VGND VPWR VPWR _35941_/D sky130_fd_sc_hd__clkbuf_1
XPHY_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16386_ _33631_/Q _33567_/Q _33503_/Q _33439_/Q _16141_/X _16142_/X VGND VGND VPWR
+ VPWR _16386_/X sky130_fd_sc_hd__mux4_1
XFILLER_185_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18125_ _17864_/X _18123_/X _18124_/X _17869_/X VGND VGND VPWR VPWR _18125_/X sky130_fd_sc_hd__a22o_1
X_30403_ _30403_/A VGND VGND VPWR VPWR _35444_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34171_ _34877_/CLK _34171_/D VGND VGND VPWR VPWR _34171_/Q sky130_fd_sc_hd__dfxtp_1
X_31383_ _27788_/X _35909_/Q _31387_/S VGND VGND VPWR VPWR _31384_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33122_ _36002_/CLK _33122_/D VGND VGND VPWR VPWR _33122_/Q sky130_fd_sc_hd__dfxtp_1
X_30334_ _30334_/A VGND VGND VPWR VPWR _35412_/D sky130_fd_sc_hd__clkbuf_1
X_18056_ _35470_/Q _35406_/Q _35342_/Q _35278_/Q _17960_/X _17961_/X VGND VGND VPWR
+ VPWR _18056_/X sky130_fd_sc_hd__mux4_1
XFILLER_144_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17007_ _17003_/X _17004_/X _17005_/X _17006_/X VGND VGND VPWR VPWR _17007_/X sky130_fd_sc_hd__a22o_1
X_33053_ _35805_/CLK _33053_/D VGND VGND VPWR VPWR _33053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_503_CLK clkbuf_6_2__f_CLK/X VGND VGND VPWR VPWR _36070_/CLK sky130_fd_sc_hd__clkbuf_16
X_30265_ _30265_/A VGND VGND VPWR VPWR _35379_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32004_ _36202_/CLK _32004_/D VGND VGND VPWR VPWR _32004_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30196_ _35347_/Q _29518_/X _30200_/S VGND VGND VPWR VPWR _30197_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18958_ _19311_/A VGND VGND VPWR VPWR _18958_/X sky130_fd_sc_hd__buf_4
XFILLER_234_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17909_ _34186_/Q _34122_/Q _34058_/Q _33994_/Q _17799_/X _17800_/X VGND VGND VPWR
+ VPWR _17909_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33955_ _34148_/CLK _33955_/D VGND VGND VPWR VPWR _33955_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18889_ _35172_/Q _35108_/Q _35044_/Q _32164_/Q _18604_/X _18605_/X VGND VGND VPWR
+ VPWR _18889_/X sky130_fd_sc_hd__mux4_1
XFILLER_230_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20920_ _33885_/Q _33821_/Q _33757_/Q _36061_/Q _20918_/X _20919_/X VGND VGND VPWR
+ VPWR _20920_/X sky130_fd_sc_hd__mux4_1
X_32906_ _32906_/CLK _32906_/D VGND VGND VPWR VPWR _32906_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33886_ _36128_/CLK _33886_/D VGND VGND VPWR VPWR _33886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20851_ _32603_/Q _32539_/Q _32475_/Q _35931_/Q _20817_/X _22317_/A VGND VGND VPWR
+ VPWR _20851_/X sky130_fd_sc_hd__mux4_1
X_32837_ _32901_/CLK _32837_/D VGND VGND VPWR VPWR _32837_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35625_ _35625_/CLK _35625_/D VGND VGND VPWR VPWR _35625_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23570_ _23702_/S VGND VGND VPWR VPWR _23589_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_39_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35556_ _35747_/CLK _35556_/D VGND VGND VPWR VPWR _35556_/Q sky130_fd_sc_hd__dfxtp_1
X_20782_ _33881_/Q _33817_/Q _33753_/Q _36057_/Q _20712_/X _20713_/X VGND VGND VPWR
+ VPWR _20782_/X sky130_fd_sc_hd__mux4_1
X_32768_ _32896_/CLK _32768_/D VGND VGND VPWR VPWR _32768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34507_ _35208_/CLK _34507_/D VGND VGND VPWR VPWR _34507_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22521_ _32138_/Q _32330_/Q _32394_/Q _35914_/Q _22233_/X _22374_/X VGND VGND VPWR
+ VPWR _22521_/X sky130_fd_sc_hd__mux4_1
XFILLER_22_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31719_ _36068_/Q input6/X _31729_/S VGND VGND VPWR VPWR _31720_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35487_ _35551_/CLK _35487_/D VGND VGND VPWR VPWR _35487_/Q sky130_fd_sc_hd__dfxtp_1
X_32699_ _32891_/CLK _32699_/D VGND VGND VPWR VPWR _32699_/Q sky130_fd_sc_hd__dfxtp_1
X_25240_ _25267_/S VGND VGND VPWR VPWR _25259_/S sky130_fd_sc_hd__buf_4
X_34438_ _36165_/CLK _34438_/D VGND VGND VPWR VPWR _34438_/Q sky130_fd_sc_hd__dfxtp_1
X_22452_ _35656_/Q _35016_/Q _34376_/Q _33736_/Q _22450_/X _22451_/X VGND VGND VPWR
+ VPWR _22452_/X sky130_fd_sc_hd__mux4_1
XFILLER_176_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21403_ _21756_/A VGND VGND VPWR VPWR _21403_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_109_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25171_ _33063_/Q _23283_/X _25175_/S VGND VGND VPWR VPWR _25172_/A sky130_fd_sc_hd__mux2_1
X_22383_ _35462_/Q _35398_/Q _35334_/Q _35270_/Q _22207_/X _22208_/X VGND VGND VPWR
+ VPWR _22383_/X sky130_fd_sc_hd__mux4_1
X_34369_ _35777_/CLK _34369_/D VGND VGND VPWR VPWR _34369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36108_ _36109_/CLK _36108_/D VGND VGND VPWR VPWR _36108_/Q sky130_fd_sc_hd__dfxtp_1
X_24122_ _32599_/Q _23234_/X _24138_/S VGND VGND VPWR VPWR _24123_/A sky130_fd_sc_hd__mux2_1
XFILLER_175_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21334_ _34920_/Q _34856_/Q _34792_/Q _34728_/Q _21054_/X _21055_/X VGND VGND VPWR
+ VPWR _21334_/X sky130_fd_sc_hd__mux4_1
XFILLER_108_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28930_ _28930_/A VGND VGND VPWR VPWR _34776_/D sky130_fd_sc_hd__clkbuf_1
X_36039_ _36039_/CLK _36039_/D VGND VGND VPWR VPWR _36039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24053_ _22993_/X _32568_/Q _24063_/S VGND VGND VPWR VPWR _24054_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21265_ _21265_/A _21265_/B _21265_/C _21265_/D VGND VGND VPWR VPWR _21266_/A sky130_fd_sc_hd__or4_4
Xclkbuf_leaf_50_CLK clkbuf_leaf_57_CLK/A VGND VGND VPWR VPWR _35947_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_173_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23004_ _23004_/A VGND VGND VPWR VPWR _32059_/D sky130_fd_sc_hd__clkbuf_1
X_20216_ _20212_/X _20213_/X _20214_/X _20215_/X VGND VGND VPWR VPWR _20216_/X sky130_fd_sc_hd__a22o_1
X_28861_ _34744_/Q _27140_/X _28871_/S VGND VGND VPWR VPWR _28862_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_1338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21196_ _21196_/A VGND VGND VPWR VPWR _36196_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27812_ _27812_/A VGND VGND VPWR VPWR _34252_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_235_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20147_ _20147_/A VGND VGND VPWR VPWR _20147_/X sky130_fd_sc_hd__buf_2
XFILLER_132_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28792_ _34711_/Q _27038_/X _28808_/S VGND VGND VPWR VPWR _28793_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27743_ _27742_/X _34230_/Q _27764_/S VGND VGND VPWR VPWR _27744_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24955_ _24995_/S VGND VGND VPWR VPWR _24983_/S sky130_fd_sc_hd__buf_4
XTAP_4136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20078_ _20073_/X _20075_/X _20076_/X _20077_/X VGND VGND VPWR VPWR _20078_/X sky130_fd_sc_hd__a22o_1
XTAP_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_218_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23906_ _22977_/X _32499_/Q _23906_/S VGND VGND VPWR VPWR _23907_/A sky130_fd_sc_hd__mux2_1
XTAP_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27674_ _27838_/S VGND VGND VPWR VPWR _27702_/S sky130_fd_sc_hd__buf_4
XFILLER_18_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24886_ input21/X VGND VGND VPWR VPWR _24886_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29413_ input20/X VGND VGND VPWR VPWR _29413_/X sky130_fd_sc_hd__buf_2
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26625_ _26625_/A VGND VGND VPWR VPWR _31147_/B sky130_fd_sc_hd__buf_4
XTAP_3468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23837_ _23837_/A VGND VGND VPWR VPWR _32403_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29344_ _29344_/A VGND VGND VPWR VPWR _34970_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26556_ _24896_/X _33717_/Q _26572_/S VGND VGND VPWR VPWR _26557_/A sky130_fd_sc_hd__mux2_1
X_23768_ _23768_/A VGND VGND VPWR VPWR _32370_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25507_ _24945_/X _33221_/Q _25511_/S VGND VGND VPWR VPWR _25508_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22719_ _22715_/X _22718_/X _22457_/X VGND VGND VPWR VPWR _22727_/C sky130_fd_sc_hd__o21ba_1
XFILLER_158_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29275_ _29275_/A VGND VGND VPWR VPWR _34940_/D sky130_fd_sc_hd__clkbuf_1
X_26487_ _26487_/A VGND VGND VPWR VPWR _33685_/D sky130_fd_sc_hd__clkbuf_1
X_23699_ _23699_/A VGND VGND VPWR VPWR _32339_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16240_ _16091_/X _16238_/X _16239_/X _16101_/X VGND VGND VPWR VPWR _16240_/X sky130_fd_sc_hd__a22o_1
X_28226_ _28226_/A VGND VGND VPWR VPWR _34444_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25438_ _24843_/X _33188_/Q _25448_/S VGND VGND VPWR VPWR _25439_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25369_ _25369_/A VGND VGND VPWR VPWR _33156_/D sky130_fd_sc_hd__clkbuf_1
X_16171_ _16877_/A VGND VGND VPWR VPWR _16171_/X sky130_fd_sc_hd__buf_6
X_28157_ _28157_/A VGND VGND VPWR VPWR _34411_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27108_ _27108_/A VGND VGND VPWR VPWR _33965_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28088_ _34379_/Q _27199_/X _28100_/S VGND VGND VPWR VPWR _28089_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19930_ _32642_/Q _32578_/Q _32514_/Q _35970_/Q _19929_/X _19713_/X VGND VGND VPWR
+ VPWR _19930_/X sky130_fd_sc_hd__mux4_1
X_27039_ _33943_/Q _27038_/X _27063_/S VGND VGND VPWR VPWR _27040_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_41_CLK clkbuf_6_7__f_CLK/X VGND VGND VPWR VPWR _36007_/CLK sky130_fd_sc_hd__clkbuf_16
X_30050_ _30050_/A VGND VGND VPWR VPWR _35277_/D sky130_fd_sc_hd__clkbuf_1
X_19861_ _33920_/Q _33856_/Q _33792_/Q _36096_/Q _19677_/X _19678_/X VGND VGND VPWR
+ VPWR _19861_/X sky130_fd_sc_hd__mux4_1
XFILLER_123_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_5_1_0_CLK clkbuf_5_7_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_1_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_190_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18812_ _18808_/X _18811_/X _18734_/X _18735_/X VGND VGND VPWR VPWR _18829_/B sky130_fd_sc_hd__o211a_1
XTAP_6050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput93 _31970_/Q VGND VGND VPWR VPWR D1[12] sky130_fd_sc_hd__buf_2
XFILLER_7_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19792_ _19720_/X _19790_/X _19791_/X _19724_/X VGND VGND VPWR VPWR _19792_/X sky130_fd_sc_hd__a22o_1
XFILLER_228_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18743_ _33056_/Q _32032_/Q _35808_/Q _35744_/Q _18672_/X _18673_/X VGND VGND VPWR
+ VPWR _18743_/X sky130_fd_sc_hd__mux4_1
XFILLER_231_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_926 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33740_ _35661_/CLK _33740_/D VGND VGND VPWR VPWR _33740_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18674_ _33054_/Q _32030_/Q _35806_/Q _35742_/Q _18672_/X _18673_/X VGND VGND VPWR
+ VPWR _18674_/X sky130_fd_sc_hd__mux4_1
X_30952_ _35705_/Q input29/X _30960_/S VGND VGND VPWR VPWR _30953_/A sky130_fd_sc_hd__mux2_1
XTAP_4670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17625_ _33410_/Q _33346_/Q _33282_/Q _33218_/Q _17480_/X _17481_/X VGND VGND VPWR
+ VPWR _17625_/X sky130_fd_sc_hd__mux4_1
XTAP_4692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33671_ _34179_/CLK _33671_/D VGND VGND VPWR VPWR _33671_/Q sky130_fd_sc_hd__dfxtp_1
X_30883_ _35672_/Q input23/X _30897_/S VGND VGND VPWR VPWR _30884_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35410_ _35666_/CLK _35410_/D VGND VGND VPWR VPWR _35410_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32622_ _36015_/CLK _32622_/D VGND VGND VPWR VPWR _32622_/Q sky130_fd_sc_hd__dfxtp_1
X_17556_ _34176_/Q _34112_/Q _34048_/Q _33984_/Q _17446_/X _17447_/X VGND VGND VPWR
+ VPWR _17556_/X sky130_fd_sc_hd__mux4_1
XFILLER_17_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35341_ _35853_/CLK _35341_/D VGND VGND VPWR VPWR _35341_/Q sky130_fd_sc_hd__dfxtp_1
X_16507_ _33122_/Q _36002_/Q _32994_/Q _32930_/Q _16356_/X _16357_/X VGND VGND VPWR
+ VPWR _16507_/X sky130_fd_sc_hd__mux4_1
XFILLER_60_962 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32553_ _35947_/CLK _32553_/D VGND VGND VPWR VPWR _32553_/Q sky130_fd_sc_hd__dfxtp_1
X_17487_ _32638_/Q _32574_/Q _32510_/Q _35966_/Q _17276_/X _17413_/X VGND VGND VPWR
+ VPWR _17487_/X sky130_fd_sc_hd__mux4_1
XFILLER_31_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31504_ _27766_/X _35966_/Q _31522_/S VGND VGND VPWR VPWR _31505_/A sky130_fd_sc_hd__mux2_1
X_19226_ _19006_/X _19224_/X _19225_/X _19012_/X VGND VGND VPWR VPWR _19226_/X sky130_fd_sc_hd__a22o_1
X_35272_ _35466_/CLK _35272_/D VGND VGND VPWR VPWR _35272_/Q sky130_fd_sc_hd__dfxtp_1
X_16438_ _17998_/A VGND VGND VPWR VPWR _16438_/X sky130_fd_sc_hd__buf_6
XFILLER_165_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32484_ _36007_/CLK _32484_/D VGND VGND VPWR VPWR _32484_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34223_ _35822_/CLK _34223_/D VGND VGND VPWR VPWR _34223_/Q sky130_fd_sc_hd__dfxtp_1
X_31435_ _31435_/A VGND VGND VPWR VPWR _35933_/D sky130_fd_sc_hd__clkbuf_1
X_19157_ _19153_/X _19154_/X _19155_/X _19156_/X VGND VGND VPWR VPWR _19157_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_1275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16369_ _35614_/Q _34974_/Q _34334_/Q _33694_/Q _16053_/X _16055_/X VGND VGND VPWR
+ VPWR _16369_/X sky130_fd_sc_hd__mux4_1
XFILLER_157_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18108_ _17153_/A _18106_/X _18107_/X _17156_/A VGND VGND VPWR VPWR _18108_/X sky130_fd_sc_hd__a22o_1
XFILLER_11_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34154_ _35627_/CLK _34154_/D VGND VGND VPWR VPWR _34154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_864 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19088_ _20147_/A VGND VGND VPWR VPWR _19088_/X sky130_fd_sc_hd__clkbuf_4
X_31366_ _27763_/X _35901_/Q _31366_/S VGND VGND VPWR VPWR _31367_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33105_ _35855_/CLK _33105_/D VGND VGND VPWR VPWR _33105_/Q sky130_fd_sc_hd__dfxtp_1
X_18039_ _33678_/Q _33614_/Q _33550_/Q _33486_/Q _17906_/X _17907_/X VGND VGND VPWR
+ VPWR _18039_/X sky130_fd_sc_hd__mux4_1
X_30317_ _35404_/Q _29497_/X _30327_/S VGND VGND VPWR VPWR _30318_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34085_ _34085_/CLK _34085_/D VGND VGND VPWR VPWR _34085_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_236_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31297_ _27661_/X _35868_/Q _31303_/S VGND VGND VPWR VPWR _31298_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_32_CLK clkbuf_6_5__f_CLK/X VGND VGND VPWR VPWR _36129_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_114_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33036_ _35852_/CLK _33036_/D VGND VGND VPWR VPWR _33036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21050_ _21756_/A VGND VGND VPWR VPWR _21050_/X sky130_fd_sc_hd__buf_4
XFILLER_236_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30248_ _35371_/Q _29395_/X _30264_/S VGND VGND VPWR VPWR _30249_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20001_ _32900_/Q _32836_/Q _32772_/Q _32708_/Q _19999_/X _20000_/X VGND VGND VPWR
+ VPWR _20001_/X sky130_fd_sc_hd__mux4_1
XFILLER_232_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30179_ _30179_/A VGND VGND VPWR VPWR _35338_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_246_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34987_ _34987_/CLK _34987_/D VGND VGND VPWR VPWR _34987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21952_ _35706_/Q _32215_/Q _35578_/Q _35514_/Q _21917_/X _21918_/X VGND VGND VPWR
+ VPWR _21952_/X sky130_fd_sc_hd__mux4_1
X_24740_ _23002_/X _32891_/Q _24744_/S VGND VGND VPWR VPWR _24741_/A sky130_fd_sc_hd__mux2_1
X_33938_ _36115_/CLK _33938_/D VGND VGND VPWR VPWR _33938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20903_ _34652_/Q _34588_/Q _34524_/Q _34460_/Q _20833_/X _20834_/X VGND VGND VPWR
+ VPWR _20903_/X sky130_fd_sc_hd__mux4_1
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24671_ _22900_/X _32858_/Q _24681_/S VGND VGND VPWR VPWR _24672_/A sky130_fd_sc_hd__mux2_1
X_33869_ _33869_/CLK _33869_/D VGND VGND VPWR VPWR _33869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21883_ _21667_/X _21881_/X _21882_/X _21671_/X VGND VGND VPWR VPWR _21883_/X sky130_fd_sc_hd__a22o_1
XFILLER_243_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_99_CLK clkbuf_leaf_99_CLK/A VGND VGND VPWR VPWR _36211_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26410_ _26410_/A VGND VGND VPWR VPWR _33648_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23622_ _23622_/A VGND VGND VPWR VPWR _32302_/D sky130_fd_sc_hd__clkbuf_1
X_35608_ _35609_/CLK _35608_/D VGND VGND VPWR VPWR _35608_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20834_ _22599_/A VGND VGND VPWR VPWR _20834_/X sky130_fd_sc_hd__buf_6
X_27390_ _27390_/A VGND VGND VPWR VPWR _34079_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26341_ _26341_/A VGND VGND VPWR VPWR _33616_/D sky130_fd_sc_hd__clkbuf_1
X_23553_ _32271_/Q _23478_/X _23557_/S VGND VGND VPWR VPWR _23554_/A sky130_fd_sc_hd__mux2_1
XFILLER_223_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20765_ _20660_/X _20763_/X _20764_/X _20672_/X VGND VGND VPWR VPWR _20765_/X sky130_fd_sc_hd__a22o_1
X_35539_ _35730_/CLK _35539_/D VGND VGND VPWR VPWR _35539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_945 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22504_ _22504_/A VGND VGND VPWR VPWR _36233_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_995 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29060_ _34838_/Q _27033_/X _29078_/S VGND VGND VPWR VPWR _29061_/A sky130_fd_sc_hd__mux2_1
X_26272_ _26272_/A VGND VGND VPWR VPWR _33583_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23484_ input55/X VGND VGND VPWR VPWR _23484_/X sky130_fd_sc_hd__buf_4
X_20696_ _22466_/A VGND VGND VPWR VPWR _20696_/X sky130_fd_sc_hd__buf_4
XFILLER_126_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25223_ _25223_/A VGND VGND VPWR VPWR _33087_/D sky130_fd_sc_hd__clkbuf_1
X_28011_ _28011_/A VGND VGND VPWR VPWR _34342_/D sky130_fd_sc_hd__clkbuf_1
X_22435_ _33416_/Q _33352_/Q _33288_/Q _33224_/Q _22433_/X _22434_/X VGND VGND VPWR
+ VPWR _22435_/X sky130_fd_sc_hd__mux4_1
XFILLER_155_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25154_ _33055_/Q _23258_/X _25154_/S VGND VGND VPWR VPWR _25155_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22366_ _22366_/A VGND VGND VPWR VPWR _22366_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_151_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24105_ _23070_/X _32593_/Q _24105_/S VGND VGND VPWR VPWR _24106_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21317_ _32872_/Q _32808_/Q _32744_/Q _32680_/Q _21240_/X _21241_/X VGND VGND VPWR
+ VPWR _21317_/X sky130_fd_sc_hd__mux4_1
XFILLER_163_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25085_ _24927_/X _33023_/Q _25101_/S VGND VGND VPWR VPWR _25086_/A sky130_fd_sc_hd__mux2_1
X_29962_ _29962_/A VGND VGND VPWR VPWR _35235_/D sky130_fd_sc_hd__clkbuf_1
X_22297_ _22012_/X _22295_/X _22296_/X _22018_/X VGND VGND VPWR VPWR _22297_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_23_CLK clkbuf_6_4__f_CLK/X VGND VGND VPWR VPWR _36210_/CLK sky130_fd_sc_hd__clkbuf_16
X_28913_ _34769_/Q _27217_/X _28913_/S VGND VGND VPWR VPWR _28914_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24036_ _22968_/X _32560_/Q _24042_/S VGND VGND VPWR VPWR _24037_/A sky130_fd_sc_hd__mux2_1
X_21248_ _22462_/A VGND VGND VPWR VPWR _21248_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_105_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29893_ _35203_/Q _29469_/X _29901_/S VGND VGND VPWR VPWR _29894_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28844_ _34736_/Q _27115_/X _28850_/S VGND VGND VPWR VPWR _28845_/A sky130_fd_sc_hd__mux2_1
X_21179_ _35684_/Q _32191_/Q _35556_/Q _35492_/Q _20858_/X _20859_/X VGND VGND VPWR
+ VPWR _21179_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28775_ _28775_/A VGND VGND VPWR VPWR _34704_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25987_ _25987_/A VGND VGND VPWR VPWR _33448_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27726_ input20/X VGND VGND VPWR VPWR _27726_/X sky130_fd_sc_hd__buf_2
XTAP_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24938_ _24938_/A VGND VGND VPWR VPWR _32962_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_1214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27657_ _27657_/A VGND VGND VPWR VPWR _34202_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24869_ _24868_/X _32940_/Q _24890_/S VGND VGND VPWR VPWR _24870_/A sky130_fd_sc_hd__mux2_1
XTAP_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17410_ _17206_/X _17408_/X _17409_/X _17209_/X VGND VGND VPWR VPWR _17410_/X sky130_fd_sc_hd__a22o_1
XTAP_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26608_ _24973_/X _33742_/Q _26614_/S VGND VGND VPWR VPWR _26609_/A sky130_fd_sc_hd__mux2_1
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18390_ _20073_/A VGND VGND VPWR VPWR _19458_/A sky130_fd_sc_hd__buf_12
XFILLER_57_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27588_ _27588_/A VGND VGND VPWR VPWR _34173_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29327_ _29327_/A VGND VGND VPWR VPWR _34965_/D sky130_fd_sc_hd__clkbuf_1
X_17341_ _17337_/X _17340_/X _17132_/X VGND VGND VPWR VPWR _17371_/A sky130_fd_sc_hd__o21ba_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26539_ _24871_/X _33709_/Q _26551_/S VGND VGND VPWR VPWR _26540_/A sky130_fd_sc_hd__mux2_1
XFILLER_199_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17272_ _33400_/Q _33336_/Q _33272_/Q _33208_/Q _17127_/X _17128_/X VGND VGND VPWR
+ VPWR _17272_/X sky130_fd_sc_hd__mux4_1
X_29258_ _34932_/Q _27127_/X _29276_/S VGND VGND VPWR VPWR _29259_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19011_ _33128_/Q _36008_/Q _33000_/Q _32936_/Q _19009_/X _19010_/X VGND VGND VPWR
+ VPWR _19011_/X sky130_fd_sc_hd__mux4_1
XFILLER_224_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28209_ _28209_/A VGND VGND VPWR VPWR _34436_/D sky130_fd_sc_hd__clkbuf_1
X_16223_ _32858_/Q _32794_/Q _32730_/Q _32666_/Q _16037_/X _16039_/X VGND VGND VPWR
+ VPWR _16223_/X sky130_fd_sc_hd__mux4_1
X_29189_ _34900_/Q _27226_/X _29191_/S VGND VGND VPWR VPWR _29190_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31220_ _31220_/A VGND VGND VPWR VPWR _35831_/D sky130_fd_sc_hd__clkbuf_1
X_16154_ _33112_/Q _35992_/Q _32984_/Q _32920_/Q _16024_/X _16025_/X VGND VGND VPWR
+ VPWR _16154_/X sky130_fd_sc_hd__mux4_1
XFILLER_155_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31151_ _31151_/A VGND VGND VPWR VPWR _35798_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16085_ _17011_/A VGND VGND VPWR VPWR _16085_/X sky130_fd_sc_hd__buf_4
XFILLER_114_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_14_CLK clkbuf_6_3__f_CLK/X VGND VGND VPWR VPWR _35365_/CLK sky130_fd_sc_hd__clkbuf_16
X_30102_ _35302_/Q _29379_/X _30108_/S VGND VGND VPWR VPWR _30103_/A sky130_fd_sc_hd__mux2_1
X_19913_ _34689_/Q _34625_/Q _34561_/Q _34497_/Q _19592_/X _19593_/X VGND VGND VPWR
+ VPWR _19913_/X sky130_fd_sc_hd__mux4_1
XFILLER_177_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31082_ _31082_/A VGND VGND VPWR VPWR _35766_/D sky130_fd_sc_hd__clkbuf_1
X_34910_ _34911_/CLK _34910_/D VGND VGND VPWR VPWR _34910_/Q sky130_fd_sc_hd__dfxtp_1
X_19844_ _35199_/Q _35135_/Q _35071_/Q _32255_/Q _19663_/X _19664_/X VGND VGND VPWR
+ VPWR _19844_/X sky130_fd_sc_hd__mux4_1
X_30033_ _30033_/A VGND VGND VPWR VPWR _35269_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_934 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35890_ _35955_/CLK _35890_/D VGND VGND VPWR VPWR _35890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34841_ _34907_/CLK _34841_/D VGND VGND VPWR VPWR _34841_/Q sky130_fd_sc_hd__dfxtp_1
X_19775_ _19775_/A _19775_/B _19775_/C _19775_/D VGND VGND VPWR VPWR _19776_/A sky130_fd_sc_hd__or4_2
X_16987_ _16853_/X _16985_/X _16986_/X _16856_/X VGND VGND VPWR VPWR _16987_/X sky130_fd_sc_hd__a22o_1
XFILLER_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18726_ _20138_/A VGND VGND VPWR VPWR _18726_/X sky130_fd_sc_hd__clkbuf_4
X_34772_ _34964_/CLK _34772_/D VGND VGND VPWR VPWR _34772_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31984_ _34918_/CLK _31984_/D VGND VGND VPWR VPWR _31984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33723_ _35644_/CLK _33723_/D VGND VGND VPWR VPWR _33723_/Q sky130_fd_sc_hd__dfxtp_1
X_18657_ _20207_/A VGND VGND VPWR VPWR _18657_/X sky130_fd_sc_hd__clkbuf_4
X_30935_ _35697_/Q input20/X _30939_/S VGND VGND VPWR VPWR _30936_/A sky130_fd_sc_hd__mux2_1
XFILLER_236_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17608_ _17961_/A VGND VGND VPWR VPWR _17608_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_18_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33654_ _34166_/CLK _33654_/D VGND VGND VPWR VPWR _33654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30866_ _30866_/A VGND VGND VPWR VPWR _35664_/D sky130_fd_sc_hd__clkbuf_1
X_18588_ _20134_/A VGND VGND VPWR VPWR _18588_/X sky130_fd_sc_hd__buf_4
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32605_ _32797_/CLK _32605_/D VGND VGND VPWR VPWR _32605_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17539_ _35455_/Q _35391_/Q _35327_/Q _35263_/Q _17254_/X _17255_/X VGND VGND VPWR
+ VPWR _17539_/X sky130_fd_sc_hd__mux4_1
X_33585_ _33904_/CLK _33585_/D VGND VGND VPWR VPWR _33585_/Q sky130_fd_sc_hd__dfxtp_1
X_30797_ _30797_/A VGND VGND VPWR VPWR _35631_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35324_ _35708_/CLK _35324_/D VGND VGND VPWR VPWR _35324_/Q sky130_fd_sc_hd__dfxtp_1
X_20550_ _34197_/Q _34133_/Q _34069_/Q _34005_/Q _18349_/X _18350_/X VGND VGND VPWR
+ VPWR _20550_/X sky130_fd_sc_hd__mux4_1
X_32536_ _35992_/CLK _32536_/D VGND VGND VPWR VPWR _32536_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19209_ _19100_/X _19207_/X _19208_/X _19103_/X VGND VGND VPWR VPWR _19209_/X sky130_fd_sc_hd__a22o_1
XFILLER_242_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35255_ _35320_/CLK _35255_/D VGND VGND VPWR VPWR _35255_/Q sky130_fd_sc_hd__dfxtp_1
X_20481_ _35218_/Q _35154_/Q _35090_/Q _32274_/Q _18392_/X _18394_/X VGND VGND VPWR
+ VPWR _20481_/X sky130_fd_sc_hd__mux4_1
X_32467_ _36079_/CLK _32467_/D VGND VGND VPWR VPWR _32467_/Q sky130_fd_sc_hd__dfxtp_1
X_34206_ _36235_/CLK _34206_/D VGND VGND VPWR VPWR _34206_/Q sky130_fd_sc_hd__dfxtp_1
X_22220_ _22220_/A _22220_/B _22220_/C _22220_/D VGND VGND VPWR VPWR _22221_/A sky130_fd_sc_hd__or4_4
XFILLER_118_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31418_ _31418_/A _31418_/B VGND VGND VPWR VPWR _31551_/S sky130_fd_sc_hd__nand2_8
XFILLER_118_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35186_ _35828_/CLK _35186_/D VGND VGND VPWR VPWR _35186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32398_ _35921_/CLK _32398_/D VGND VGND VPWR VPWR _32398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_1438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22151_ _22151_/A VGND VGND VPWR VPWR _36223_/D sky130_fd_sc_hd__clkbuf_1
X_34137_ _36219_/CLK _34137_/D VGND VGND VPWR VPWR _34137_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31349_ _31349_/A VGND VGND VPWR VPWR _35892_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21102_ _33890_/Q _33826_/Q _33762_/Q _36066_/Q _20918_/X _20919_/X VGND VGND VPWR
+ VPWR _21102_/X sky130_fd_sc_hd__mux4_1
XFILLER_156_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34068_ _34773_/CLK _34068_/D VGND VGND VPWR VPWR _34068_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22082_ _33406_/Q _33342_/Q _33278_/Q _33214_/Q _22080_/X _22081_/X VGND VGND VPWR
+ VPWR _22082_/X sky130_fd_sc_hd__mux4_1
XTAP_6819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25910_ _24942_/X _33412_/Q _25916_/S VGND VGND VPWR VPWR _25911_/A sky130_fd_sc_hd__mux2_1
X_21033_ _20961_/X _21031_/X _21032_/X _20965_/X VGND VGND VPWR VPWR _21033_/X sky130_fd_sc_hd__a22o_1
X_33019_ _35191_/CLK _33019_/D VGND VGND VPWR VPWR _33019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_232_1015 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26890_ _33874_/Q _23487_/X _26896_/S VGND VGND VPWR VPWR _26891_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25841_ _24840_/X _33379_/Q _25853_/S VGND VGND VPWR VPWR _25842_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28560_ _28560_/A VGND VGND VPWR VPWR _34602_/D sky130_fd_sc_hd__clkbuf_1
X_25772_ _25772_/A VGND VGND VPWR VPWR _33346_/D sky130_fd_sc_hd__clkbuf_1
X_22984_ input25/X VGND VGND VPWR VPWR _22984_/X sky130_fd_sc_hd__buf_2
XFILLER_227_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27511_ _27511_/A VGND VGND VPWR VPWR _34136_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24723_ _22977_/X _32883_/Q _24723_/S VGND VGND VPWR VPWR _24724_/A sky130_fd_sc_hd__mux2_1
X_28491_ _27804_/X _34570_/Q _28505_/S VGND VGND VPWR VPWR _28492_/A sky130_fd_sc_hd__mux2_1
X_21935_ _33658_/Q _33594_/Q _33530_/Q _33466_/Q _21800_/X _21801_/X VGND VGND VPWR
+ VPWR _21935_/X sky130_fd_sc_hd__mux4_1
XFILLER_43_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27442_ _34104_/Q _27140_/X _27452_/S VGND VGND VPWR VPWR _27443_/A sky130_fd_sc_hd__mux2_1
XFILLER_231_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24654_ _24654_/A VGND VGND VPWR VPWR _32850_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21866_ _21862_/X _21865_/X _21765_/X VGND VGND VPWR VPWR _21867_/D sky130_fd_sc_hd__o21ba_1
XFILLER_128_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20817_ _22582_/A VGND VGND VPWR VPWR _20817_/X sky130_fd_sc_hd__buf_6
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23605_ _23605_/A VGND VGND VPWR VPWR _32294_/D sky130_fd_sc_hd__clkbuf_1
X_27373_ _34071_/Q _27038_/X _27389_/S VGND VGND VPWR VPWR _27374_/A sky130_fd_sc_hd__mux2_1
X_21797_ _21797_/A _21797_/B _21797_/C _21797_/D VGND VGND VPWR VPWR _21798_/A sky130_fd_sc_hd__or4_1
X_24585_ _24585_/A VGND VGND VPWR VPWR _32817_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29112_ _34863_/Q _27112_/X _29120_/S VGND VGND VPWR VPWR _29113_/A sky130_fd_sc_hd__mux2_1
X_26324_ _24954_/X _33608_/Q _26342_/S VGND VGND VPWR VPWR _26325_/A sky130_fd_sc_hd__mux2_1
XFILLER_243_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23536_ _32263_/Q _23450_/X _23536_/S VGND VGND VPWR VPWR _23537_/A sky130_fd_sc_hd__mux2_1
X_20748_ _33368_/Q _33304_/Q _33240_/Q _33176_/Q _20602_/X _20603_/X VGND VGND VPWR
+ VPWR _20748_/X sky130_fd_sc_hd__mux4_1
XFILLER_211_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29043_ _29043_/A VGND VGND VPWR VPWR _34830_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_1442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23467_ _32234_/Q _23466_/X _23485_/S VGND VGND VPWR VPWR _23468_/A sky130_fd_sc_hd__mux2_1
X_26255_ _26255_/A VGND VGND VPWR VPWR _33575_/D sky130_fd_sc_hd__clkbuf_1
X_20679_ _22535_/A VGND VGND VPWR VPWR _20679_/X sky130_fd_sc_hd__buf_6
XFILLER_11_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22418_ _33095_/Q _32071_/Q _35847_/Q _35783_/Q _22384_/X _22385_/X VGND VGND VPWR
+ VPWR _22418_/X sky130_fd_sc_hd__mux4_1
X_25206_ _25206_/A VGND VGND VPWR VPWR _33079_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26186_ _24951_/X _33543_/Q _26186_/S VGND VGND VPWR VPWR _26187_/A sky130_fd_sc_hd__mux2_1
X_23398_ _23398_/A VGND VGND VPWR VPWR _32211_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25137_ _25137_/A VGND VGND VPWR VPWR _33046_/D sky130_fd_sc_hd__clkbuf_1
X_22349_ _34693_/Q _34629_/Q _34565_/Q _34501_/Q _22245_/X _22246_/X VGND VGND VPWR
+ VPWR _22349_/X sky130_fd_sc_hd__mux4_1
XFILLER_88_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29945_ _29945_/A VGND VGND VPWR VPWR _35227_/D sky130_fd_sc_hd__clkbuf_1
X_25068_ _24902_/X _33015_/Q _25080_/S VGND VGND VPWR VPWR _25069_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_878 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16910_ _34413_/Q _36141_/Q _34285_/Q _34221_/Q _16876_/X _16877_/X VGND VGND VPWR
+ VPWR _16910_/X sky130_fd_sc_hd__mux4_1
X_24019_ _22943_/X _32552_/Q _24021_/S VGND VGND VPWR VPWR _24020_/A sky130_fd_sc_hd__mux2_1
XFILLER_219_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17890_ _35657_/Q _35017_/Q _34377_/Q _33737_/Q _17850_/X _17851_/X VGND VGND VPWR
+ VPWR _17890_/X sky130_fd_sc_hd__mux4_1
X_29876_ _35195_/Q _29444_/X _29880_/S VGND VGND VPWR VPWR _29877_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28827_ _34728_/Q _27090_/X _28829_/S VGND VGND VPWR VPWR _28828_/A sky130_fd_sc_hd__mux2_1
X_16841_ _34923_/Q _34859_/Q _34795_/Q _34731_/Q _16807_/X _16808_/X VGND VGND VPWR
+ VPWR _16841_/X sky130_fd_sc_hd__mux4_1
XFILLER_144_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19560_ _34679_/Q _34615_/Q _34551_/Q _34487_/Q _19239_/X _19240_/X VGND VGND VPWR
+ VPWR _19560_/X sky130_fd_sc_hd__mux4_1
X_28758_ _34696_/Q _27189_/X _28776_/S VGND VGND VPWR VPWR _28759_/A sky130_fd_sc_hd__mux2_1
X_16772_ _34154_/Q _34090_/Q _34026_/Q _33962_/Q _16740_/X _16741_/X VGND VGND VPWR
+ VPWR _16772_/X sky130_fd_sc_hd__mux4_1
XFILLER_18_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18511_ _34138_/Q _34074_/Q _34010_/Q _33946_/Q _18309_/X _18311_/X VGND VGND VPWR
+ VPWR _18511_/X sky130_fd_sc_hd__mux4_1
X_27709_ _27708_/X _34219_/Q _27733_/S VGND VGND VPWR VPWR _27710_/A sky130_fd_sc_hd__mux2_1
XTAP_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19491_ _35189_/Q _35125_/Q _35061_/Q _32242_/Q _19310_/X _19311_/X VGND VGND VPWR
+ VPWR _19491_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28689_ _28689_/A VGND VGND VPWR VPWR _34663_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30720_ _35595_/Q _29494_/X _30732_/S VGND VGND VPWR VPWR _30721_/A sky130_fd_sc_hd__mux2_1
X_18442_ _20207_/A VGND VGND VPWR VPWR _18442_/X sky130_fd_sc_hd__buf_4
XFILLER_94_1239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_3_CLK clkbuf_leaf_9_CLK/A VGND VGND VPWR VPWR _34920_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18373_ _18360_/X _18365_/X _18370_/X _18372_/X VGND VGND VPWR VPWR _18373_/X sky130_fd_sc_hd__a22o_1
X_30651_ _35562_/Q _29391_/X _30669_/S VGND VGND VPWR VPWR _30652_/A sky130_fd_sc_hd__mux2_1
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17324_ _17003_/X _17322_/X _17323_/X _17006_/X VGND VGND VPWR VPWR _17324_/X sky130_fd_sc_hd__a22o_1
X_33370_ _33818_/CLK _33370_/D VGND VGND VPWR VPWR _33370_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30582_ _30582_/A VGND VGND VPWR VPWR _35529_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32321_ _35970_/CLK _32321_/D VGND VGND VPWR VPWR _32321_/Q sky130_fd_sc_hd__dfxtp_1
X_17255_ _17961_/A VGND VGND VPWR VPWR _17255_/X sky130_fd_sc_hd__buf_4
XFILLER_179_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16206_ _16091_/X _16204_/X _16205_/X _16101_/X VGND VGND VPWR VPWR _16206_/X sky130_fd_sc_hd__a22o_1
X_35040_ _36197_/CLK _35040_/D VGND VGND VPWR VPWR _35040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32252_ _35577_/CLK _32252_/D VGND VGND VPWR VPWR _32252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17186_ _35445_/Q _35381_/Q _35317_/Q _35253_/Q _16901_/X _16902_/X VGND VGND VPWR
+ VPWR _17186_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_6_50__f_CLK clkbuf_5_25_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_50__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_127_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31203_ _31203_/A VGND VGND VPWR VPWR _35823_/D sky130_fd_sc_hd__clkbuf_1
X_16137_ _16133_/X _16136_/X _16104_/X VGND VGND VPWR VPWR _16138_/D sky130_fd_sc_hd__o21ba_1
XFILLER_155_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32183_ _35677_/CLK _32183_/D VGND VGND VPWR VPWR _32183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31134_ _31134_/A VGND VGND VPWR VPWR _35791_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16068_ _17766_/A VGND VGND VPWR VPWR _17936_/A sky130_fd_sc_hd__buf_12
XFILLER_233_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31065_ _31065_/A VGND VGND VPWR VPWR _35758_/D sky130_fd_sc_hd__clkbuf_1
X_35942_ _35944_/CLK _35942_/D VGND VGND VPWR VPWR _35942_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30016_ _30016_/A VGND VGND VPWR VPWR _35261_/D sky130_fd_sc_hd__clkbuf_1
X_19827_ _19506_/X _19825_/X _19826_/X _19509_/X VGND VGND VPWR VPWR _19827_/X sky130_fd_sc_hd__a22o_1
XFILLER_29_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35873_ _35939_/CLK _35873_/D VGND VGND VPWR VPWR _35873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34824_ _34954_/CLK _34824_/D VGND VGND VPWR VPWR _34824_/Q sky130_fd_sc_hd__dfxtp_1
X_19758_ _32893_/Q _32829_/Q _32765_/Q _32701_/Q _19646_/X _19647_/X VGND VGND VPWR
+ VPWR _19758_/X sky130_fd_sc_hd__mux4_1
XFILLER_42_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18709_ _34655_/Q _34591_/Q _34527_/Q _34463_/Q _18533_/X _18534_/X VGND VGND VPWR
+ VPWR _18709_/X sky130_fd_sc_hd__mux4_1
X_34755_ _34949_/CLK _34755_/D VGND VGND VPWR VPWR _34755_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31967_ _34148_/CLK _31967_/D VGND VGND VPWR VPWR _31967_/Q sky130_fd_sc_hd__dfxtp_1
X_19689_ _35707_/Q _32216_/Q _35579_/Q _35515_/Q _19617_/X _19618_/X VGND VGND VPWR
+ VPWR _19689_/X sky130_fd_sc_hd__mux4_1
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21720_ _21405_/X _21718_/X _21719_/X _21410_/X VGND VGND VPWR VPWR _21720_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33706_ _34987_/CLK _33706_/D VGND VGND VPWR VPWR _33706_/Q sky130_fd_sc_hd__dfxtp_1
X_30918_ _35689_/Q input11/X _30918_/S VGND VGND VPWR VPWR _30919_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34686_ _35071_/CLK _34686_/D VGND VGND VPWR VPWR _34686_/Q sky130_fd_sc_hd__dfxtp_1
X_31898_ _23405_/X _36153_/Q _31906_/S VGND VGND VPWR VPWR _31899_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33637_ _34146_/CLK _33637_/D VGND VGND VPWR VPWR _33637_/Q sky130_fd_sc_hd__dfxtp_1
X_21651_ _21651_/A VGND VGND VPWR VPWR _36209_/D sky130_fd_sc_hd__clkbuf_1
X_30849_ _35656_/Q input46/X _30867_/S VGND VGND VPWR VPWR _30850_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20602_ _22399_/A VGND VGND VPWR VPWR _20602_/X sky130_fd_sc_hd__buf_4
X_24370_ _24370_/A VGND VGND VPWR VPWR _32715_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_240_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21582_ _33648_/Q _33584_/Q _33520_/Q _33456_/Q _21447_/X _21448_/X VGND VGND VPWR
+ VPWR _21582_/X sky130_fd_sc_hd__mux4_1
X_33568_ _36202_/CLK _33568_/D VGND VGND VPWR VPWR _33568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23321_ _32178_/Q _23237_/X _23335_/S VGND VGND VPWR VPWR _23322_/A sky130_fd_sc_hd__mux2_1
X_20533_ _35732_/Q _32244_/Q _35604_/Q _35540_/Q _18293_/X _18295_/X VGND VGND VPWR
+ VPWR _20533_/X sky130_fd_sc_hd__mux4_1
XFILLER_177_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32519_ _35975_/CLK _32519_/D VGND VGND VPWR VPWR _32519_/Q sky130_fd_sc_hd__dfxtp_1
X_35307_ _35433_/CLK _35307_/D VGND VGND VPWR VPWR _35307_/Q sky130_fd_sc_hd__dfxtp_1
X_33499_ _33753_/CLK _33499_/D VGND VGND VPWR VPWR _33499_/Q sky130_fd_sc_hd__dfxtp_1
X_26040_ _26040_/A VGND VGND VPWR VPWR _33473_/D sky130_fd_sc_hd__clkbuf_1
X_23252_ input62/X VGND VGND VPWR VPWR _23252_/X sky130_fd_sc_hd__buf_4
X_20464_ _20212_/X _20462_/X _20463_/X _20215_/X VGND VGND VPWR VPWR _20464_/X sky130_fd_sc_hd__a22o_1
X_35238_ _35367_/CLK _35238_/D VGND VGND VPWR VPWR _35238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22203_ _22199_/X _22202_/X _22093_/X _22094_/X VGND VGND VPWR VPWR _22220_/B sky130_fd_sc_hd__o211a_1
XFILLER_10_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23183_ _23183_/A VGND VGND VPWR VPWR _32129_/D sky130_fd_sc_hd__clkbuf_1
X_35169_ _35297_/CLK _35169_/D VGND VGND VPWR VPWR _35169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20395_ _20164_/X _20393_/X _20394_/X _20169_/X VGND VGND VPWR VPWR _20395_/X sky130_fd_sc_hd__a22o_1
XFILLER_238_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22134_ _22020_/X _22132_/X _22133_/X _22024_/X VGND VGND VPWR VPWR _22134_/X sky130_fd_sc_hd__a22o_1
XFILLER_134_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27991_ _34333_/Q _27056_/X _27995_/S VGND VGND VPWR VPWR _27992_/A sky130_fd_sc_hd__mux2_1
XTAP_6616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput250 _32445_/Q VGND VGND VPWR VPWR D3[39] sky130_fd_sc_hd__buf_2
Xoutput261 _32455_/Q VGND VGND VPWR VPWR D3[49] sky130_fd_sc_hd__buf_2
XFILLER_47_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput272 _32465_/Q VGND VGND VPWR VPWR D3[59] sky130_fd_sc_hd__buf_2
X_29730_ _29730_/A VGND VGND VPWR VPWR _35125_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26942_ _33898_/Q _23292_/X _26960_/S VGND VGND VPWR VPWR _26943_/A sky130_fd_sc_hd__mux2_1
X_22065_ _33085_/Q _32061_/Q _35837_/Q _35773_/Q _22031_/X _22032_/X VGND VGND VPWR
+ VPWR _22065_/X sky130_fd_sc_hd__mux4_1
XTAP_6649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21016_ _21016_/A _21016_/B _21016_/C _21016_/D VGND VGND VPWR VPWR _21017_/A sky130_fd_sc_hd__or4_1
XTAP_5937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29661_ _29661_/A VGND VGND VPWR VPWR _35093_/D sky130_fd_sc_hd__clkbuf_1
X_26873_ _26873_/A VGND VGND VPWR VPWR _33865_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28612_ _28612_/A VGND VGND VPWR VPWR _34627_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25824_ _24815_/X _33371_/Q _25832_/S VGND VGND VPWR VPWR _25825_/A sky130_fd_sc_hd__mux2_1
XFILLER_134_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29592_ _35060_/Q _29422_/X _29610_/S VGND VGND VPWR VPWR _29593_/A sky130_fd_sc_hd__mux2_1
XFILLER_229_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28543_ _28543_/A VGND VGND VPWR VPWR _34594_/D sky130_fd_sc_hd__clkbuf_1
X_25755_ _25755_/A VGND VGND VPWR VPWR _33338_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22967_ _22967_/A VGND VGND VPWR VPWR _32047_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_963 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24706_ _24706_/A VGND VGND VPWR VPWR _32874_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28474_ _27779_/X _34562_/Q _28484_/S VGND VGND VPWR VPWR _28475_/A sky130_fd_sc_hd__mux2_1
X_21918_ _22400_/A VGND VGND VPWR VPWR _21918_/X sky130_fd_sc_hd__buf_4
XFILLER_231_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25686_ _25686_/A VGND VGND VPWR VPWR _33305_/D sky130_fd_sc_hd__clkbuf_1
X_22898_ _22897_/X _32025_/Q _22916_/S VGND VGND VPWR VPWR _22899_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27425_ _34096_/Q _27115_/X _27431_/S VGND VGND VPWR VPWR _27426_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24637_ _23049_/X _32842_/Q _24651_/S VGND VGND VPWR VPWR _24638_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21849_ _21667_/X _21847_/X _21848_/X _21671_/X VGND VGND VPWR VPWR _21849_/X sky130_fd_sc_hd__a22o_1
XFILLER_203_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27356_ _27356_/A VGND VGND VPWR VPWR _34063_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_208_1072 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24568_ _24568_/A VGND VGND VPWR VPWR _32809_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26307_ _24930_/X _33600_/Q _26321_/S VGND VGND VPWR VPWR _26308_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23519_ _23519_/A VGND VGND VPWR VPWR _32254_/D sky130_fd_sc_hd__clkbuf_1
X_27287_ _27287_/A VGND VGND VPWR VPWR _34030_/D sky130_fd_sc_hd__clkbuf_1
X_24499_ _24499_/A VGND VGND VPWR VPWR _32776_/D sky130_fd_sc_hd__clkbuf_1
X_29026_ _29026_/A VGND VGND VPWR VPWR _34822_/D sky130_fd_sc_hd__clkbuf_1
X_17040_ _33073_/Q _32049_/Q _35825_/Q _35761_/Q _16725_/X _16726_/X VGND VGND VPWR
+ VPWR _17040_/X sky130_fd_sc_hd__mux4_1
X_26238_ _26238_/A VGND VGND VPWR VPWR _33567_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26169_ _26169_/A VGND VGND VPWR VPWR _33534_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18991_ _35175_/Q _35111_/Q _35047_/Q _32167_/Q _18957_/X _18958_/X VGND VGND VPWR
+ VPWR _18991_/X sky130_fd_sc_hd__mux4_1
XFILLER_139_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17942_ _17942_/A VGND VGND VPWR VPWR _32010_/D sky130_fd_sc_hd__clkbuf_4
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_219_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29928_ _35220_/Q _29521_/X _29930_/S VGND VGND VPWR VPWR _29929_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17873_ _17873_/A _17873_/B _17873_/C _17873_/D VGND VGND VPWR VPWR _17874_/A sky130_fd_sc_hd__or4_2
X_29859_ _35187_/Q _29419_/X _29859_/S VGND VGND VPWR VPWR _29860_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16824_ _33131_/Q _36011_/Q _33003_/Q _32939_/Q _16709_/X _16710_/X VGND VGND VPWR
+ VPWR _16824_/X sky130_fd_sc_hd__mux4_1
X_19612_ _19359_/X _19610_/X _19611_/X _19365_/X VGND VGND VPWR VPWR _19612_/X sky130_fd_sc_hd__a22o_1
X_32870_ _32873_/CLK _32870_/D VGND VGND VPWR VPWR _32870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31821_ _36117_/Q input60/X _31821_/S VGND VGND VPWR VPWR _31822_/A sky130_fd_sc_hd__mux2_1
XFILLER_207_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19543_ _19539_/X _19542_/X _19432_/X VGND VGND VPWR VPWR _19567_/A sky130_fd_sc_hd__o21ba_1
XFILLER_111_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16755_ _35689_/Q _32196_/Q _35561_/Q _35497_/Q _16611_/X _16612_/X VGND VGND VPWR
+ VPWR _16755_/X sky130_fd_sc_hd__mux4_1
XFILLER_47_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34540_ _35754_/CLK _34540_/D VGND VGND VPWR VPWR _34540_/Q sky130_fd_sc_hd__dfxtp_1
X_31752_ _31821_/S VGND VGND VPWR VPWR _31771_/S sky130_fd_sc_hd__buf_4
X_19474_ _19153_/X _19472_/X _19473_/X _19156_/X VGND VGND VPWR VPWR _19474_/X sky130_fd_sc_hd__a22o_1
XFILLER_59_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16686_ _35431_/Q _35367_/Q _35303_/Q _35239_/Q _16548_/X _16549_/X VGND VGND VPWR
+ VPWR _16686_/X sky130_fd_sc_hd__mux4_1
XFILLER_61_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_222_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18425_ _35607_/Q _34967_/Q _34327_/Q _33687_/Q _18353_/X _18355_/X VGND VGND VPWR
+ VPWR _18425_/X sky130_fd_sc_hd__mux4_1
X_30703_ _35587_/Q _29469_/X _30711_/S VGND VGND VPWR VPWR _30704_/A sky130_fd_sc_hd__mux2_1
XFILLER_206_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34471_ _35365_/CLK _34471_/D VGND VGND VPWR VPWR _34471_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31683_ _31683_/A VGND VGND VPWR VPWR _36051_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33422_ _33425_/CLK _33422_/D VGND VGND VPWR VPWR _33422_/Q sky130_fd_sc_hd__dfxtp_1
X_36210_ _36210_/CLK _36210_/D VGND VGND VPWR VPWR _36210_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_222_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18356_ _35606_/Q _34966_/Q _34326_/Q _33686_/Q _18353_/X _18355_/X VGND VGND VPWR
+ VPWR _18356_/X sky130_fd_sc_hd__mux4_1
X_30634_ _35554_/Q _29367_/X _30648_/S VGND VGND VPWR VPWR _30635_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17307_ _33913_/Q _33849_/Q _33785_/Q _36089_/Q _17024_/X _17025_/X VGND VGND VPWR
+ VPWR _17307_/X sky130_fd_sc_hd__mux4_1
X_36141_ _36141_/CLK _36141_/D VGND VGND VPWR VPWR _36141_/Q sky130_fd_sc_hd__dfxtp_1
X_33353_ _34121_/CLK _33353_/D VGND VGND VPWR VPWR _33353_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30565_ _30565_/A VGND VGND VPWR VPWR _35521_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18287_ _20207_/A VGND VGND VPWR VPWR _18287_/X sky130_fd_sc_hd__buf_4
XFILLER_147_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32304_ _32879_/CLK _32304_/D VGND VGND VPWR VPWR _32304_/Q sky130_fd_sc_hd__dfxtp_1
X_17238_ _34167_/Q _34103_/Q _34039_/Q _33975_/Q _17093_/X _17094_/X VGND VGND VPWR
+ VPWR _17238_/X sky130_fd_sc_hd__mux4_1
X_36072_ _36072_/CLK _36072_/D VGND VGND VPWR VPWR _36072_/Q sky130_fd_sc_hd__dfxtp_1
X_33284_ _33415_/CLK _33284_/D VGND VGND VPWR VPWR _33284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30496_ _30496_/A VGND VGND VPWR VPWR _35488_/D sky130_fd_sc_hd__clkbuf_1
X_35023_ _35663_/CLK _35023_/D VGND VGND VPWR VPWR _35023_/Q sky130_fd_sc_hd__dfxtp_1
X_32235_ _35724_/CLK _32235_/D VGND VGND VPWR VPWR _32235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17169_ _33653_/Q _33589_/Q _33525_/Q _33461_/Q _16847_/X _16848_/X VGND VGND VPWR
+ VPWR _17169_/X sky130_fd_sc_hd__mux4_1
XFILLER_116_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20180_ _19859_/X _20178_/X _20179_/X _19862_/X VGND VGND VPWR VPWR _20180_/X sky130_fd_sc_hd__a22o_1
X_32166_ _35176_/CLK _32166_/D VGND VGND VPWR VPWR _32166_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_1266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31117_ _31117_/A VGND VGND VPWR VPWR _35783_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_131_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32097_ _32356_/CLK _32097_/D VGND VGND VPWR VPWR _32097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35925_ _35988_/CLK _35925_/D VGND VGND VPWR VPWR _35925_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31048_ _31048_/A VGND VGND VPWR VPWR _35750_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_762 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35856_ _35857_/CLK _35856_/D VGND VGND VPWR VPWR _35856_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23870_ _23870_/A VGND VGND VPWR VPWR _32481_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22821_ _20618_/X _22819_/X _22820_/X _20627_/X VGND VGND VPWR VPWR _22821_/X sky130_fd_sc_hd__a22o_1
X_34807_ _36151_/CLK _34807_/D VGND VGND VPWR VPWR _34807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35787_ _35852_/CLK _35787_/D VGND VGND VPWR VPWR _35787_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32999_ _36007_/CLK _32999_/D VGND VGND VPWR VPWR _32999_/Q sky130_fd_sc_hd__dfxtp_1
X_25540_ _24994_/X _33237_/Q _25540_/S VGND VGND VPWR VPWR _25541_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22752_ _22459_/X _22750_/X _22751_/X _22462_/X VGND VGND VPWR VPWR _22752_/X sky130_fd_sc_hd__a22o_1
XFILLER_25_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34738_ _34927_/CLK _34738_/D VGND VGND VPWR VPWR _34738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21703_ _21659_/X _21701_/X _21702_/X _21665_/X VGND VGND VPWR VPWR _21703_/X sky130_fd_sc_hd__a22o_1
X_22683_ _35727_/Q _32238_/Q _35599_/Q _35535_/Q _20593_/X _20595_/X VGND VGND VPWR
+ VPWR _22683_/X sky130_fd_sc_hd__mux4_1
X_25471_ _25540_/S VGND VGND VPWR VPWR _25490_/S sky130_fd_sc_hd__buf_4
XFILLER_77_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34669_ _35692_/CLK _34669_/D VGND VGND VPWR VPWR _34669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27210_ _27210_/A VGND VGND VPWR VPWR _33998_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_244_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24422_ _22931_/X _32740_/Q _24432_/S VGND VGND VPWR VPWR _24423_/A sky130_fd_sc_hd__mux2_1
X_21634_ _21314_/X _21632_/X _21633_/X _21318_/X VGND VGND VPWR VPWR _21634_/X sky130_fd_sc_hd__a22o_1
XFILLER_40_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28190_ _28190_/A VGND VGND VPWR VPWR _34427_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_762 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27141_ _33976_/Q _27140_/X _27156_/S VGND VGND VPWR VPWR _27142_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24353_ _24353_/A VGND VGND VPWR VPWR _32707_/D sky130_fd_sc_hd__clkbuf_1
X_21565_ _22400_/A VGND VGND VPWR VPWR _21565_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_205_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20516_ _20512_/X _20515_/X _20171_/A VGND VGND VPWR VPWR _20517_/D sky130_fd_sc_hd__o21ba_1
XFILLER_154_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23304_ _23304_/A VGND VGND VPWR VPWR _32173_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24284_ _24284_/A VGND VGND VPWR VPWR _32674_/D sky130_fd_sc_hd__clkbuf_1
X_27072_ input4/X VGND VGND VPWR VPWR _27072_/X sky130_fd_sc_hd__buf_4
X_21496_ _21314_/X _21494_/X _21495_/X _21318_/X VGND VGND VPWR VPWR _21496_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23235_ _32151_/Q _23234_/X _23259_/S VGND VGND VPWR VPWR _23236_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26023_ _26023_/A VGND VGND VPWR VPWR _33465_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20447_ _33105_/Q _32081_/Q _35857_/Q _35793_/Q _18379_/X _18380_/X VGND VGND VPWR
+ VPWR _20447_/X sky130_fd_sc_hd__mux4_1
XFILLER_88_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23166_ _23166_/A VGND VGND VPWR VPWR _32121_/D sky130_fd_sc_hd__clkbuf_1
XTAP_7125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20378_ _20065_/X _20376_/X _20377_/X _20071_/X VGND VGND VPWR VPWR _20378_/X sky130_fd_sc_hd__a22o_1
XFILLER_107_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22117_ _22111_/X _22112_/X _22115_/X _22116_/X VGND VGND VPWR VPWR _22117_/X sky130_fd_sc_hd__a22o_1
XTAP_6424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27974_ _27974_/A VGND VGND VPWR VPWR _34325_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23097_ _23097_/A VGND VGND VPWR VPWR _32088_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29713_ _29713_/A VGND VGND VPWR VPWR _35117_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26925_ _33890_/Q _23268_/X _26939_/S VGND VGND VPWR VPWR _26926_/A sky130_fd_sc_hd__mux2_1
X_22048_ _34173_/Q _34109_/Q _34045_/Q _33981_/Q _22046_/X _22047_/X VGND VGND VPWR
+ VPWR _22048_/X sky130_fd_sc_hd__mux4_1
XTAP_6479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29644_ _35085_/Q _29500_/X _29652_/S VGND VGND VPWR VPWR _29645_/A sky130_fd_sc_hd__mux2_1
XTAP_5767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26856_ _26856_/A VGND VGND VPWR VPWR _33857_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25807_ _25807_/A VGND VGND VPWR VPWR _33363_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29575_ _35052_/Q _29398_/X _29589_/S VGND VGND VPWR VPWR _29576_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26787_ _26787_/A VGND VGND VPWR VPWR _33824_/D sky130_fd_sc_hd__clkbuf_1
X_23999_ _23999_/A VGND VGND VPWR VPWR _32542_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28526_ _28526_/A VGND VGND VPWR VPWR _34586_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16540_ _16353_/X _16538_/X _16539_/X _16359_/X VGND VGND VPWR VPWR _16540_/X sky130_fd_sc_hd__a22o_1
XFILLER_244_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25738_ _25738_/A VGND VGND VPWR VPWR _33330_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16471_ _33121_/Q _36001_/Q _32993_/Q _32929_/Q _16356_/X _16357_/X VGND VGND VPWR
+ VPWR _16471_/X sky130_fd_sc_hd__mux4_1
X_28457_ _27754_/X _34554_/Q _28463_/S VGND VGND VPWR VPWR _28458_/A sky130_fd_sc_hd__mux2_1
X_25669_ _24985_/X _33298_/Q _25675_/S VGND VGND VPWR VPWR _25670_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18210_ _34707_/Q _34643_/Q _34579_/Q _34515_/Q _17998_/X _17999_/X VGND VGND VPWR
+ VPWR _18210_/X sky130_fd_sc_hd__mux4_1
X_27408_ _34088_/Q _27090_/X _27410_/S VGND VGND VPWR VPWR _27409_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19190_ _19186_/X _19189_/X _19079_/X VGND VGND VPWR VPWR _19214_/A sky130_fd_sc_hd__o21ba_1
X_28388_ _27652_/X _34521_/Q _28400_/S VGND VGND VPWR VPWR _28389_/A sky130_fd_sc_hd__mux2_1
XFILLER_227_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18141_ _17158_/A _18139_/X _18140_/X _17163_/A VGND VGND VPWR VPWR _18141_/X sky130_fd_sc_hd__a22o_1
X_27339_ _27339_/A VGND VGND VPWR VPWR _34055_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18072_ _33423_/Q _33359_/Q _33295_/Q _33231_/Q _17833_/X _17834_/X VGND VGND VPWR
+ VPWR _18072_/X sky130_fd_sc_hd__mux4_1
X_30350_ _30350_/A VGND VGND VPWR VPWR _35419_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29009_ _34814_/Q _27158_/X _29027_/S VGND VGND VPWR VPWR _29010_/A sky130_fd_sc_hd__mux2_1
X_17023_ _33393_/Q _33329_/Q _33265_/Q _33201_/Q _16774_/X _16775_/X VGND VGND VPWR
+ VPWR _17023_/X sky130_fd_sc_hd__mux4_1
XFILLER_125_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30281_ _35387_/Q _29444_/X _30285_/S VGND VGND VPWR VPWR _30282_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32020_ _36207_/CLK _32020_/D VGND VGND VPWR VPWR _32020_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_994 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18974_ _18800_/X _18970_/X _18973_/X _18803_/X VGND VGND VPWR VPWR _18974_/X sky130_fd_sc_hd__a22o_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17925_ _35722_/Q _32233_/Q _35594_/Q _35530_/Q _17670_/X _17671_/X VGND VGND VPWR
+ VPWR _17925_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33971_ _34099_/CLK _33971_/D VGND VGND VPWR VPWR _33971_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_294_CLK clkbuf_6_56__f_CLK/X VGND VGND VPWR VPWR _35907_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_117_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35710_ _35711_/CLK _35710_/D VGND VGND VPWR VPWR _35710_/Q sky130_fd_sc_hd__dfxtp_1
X_32922_ _34007_/CLK _32922_/D VGND VGND VPWR VPWR _32922_/Q sky130_fd_sc_hd__dfxtp_1
X_17856_ _17709_/X _17854_/X _17855_/X _17712_/X VGND VGND VPWR VPWR _17856_/X sky130_fd_sc_hd__a22o_1
XFILLER_26_1188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16807_ _17866_/A VGND VGND VPWR VPWR _16807_/X sky130_fd_sc_hd__buf_4
XFILLER_26_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35641_ _35641_/CLK _35641_/D VGND VGND VPWR VPWR _35641_/Q sky130_fd_sc_hd__dfxtp_1
X_17787_ _17709_/X _17783_/X _17786_/X _17712_/X VGND VGND VPWR VPWR _17787_/X sky130_fd_sc_hd__a22o_1
X_32853_ _35989_/CLK _32853_/D VGND VGND VPWR VPWR _32853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31804_ _31804_/A VGND VGND VPWR VPWR _36108_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_207_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16738_ _16738_/A VGND VGND VPWR VPWR _31976_/D sky130_fd_sc_hd__clkbuf_1
X_19526_ _34678_/Q _34614_/Q _34550_/Q _34486_/Q _19239_/X _19240_/X VGND VGND VPWR
+ VPWR _19526_/X sky130_fd_sc_hd__mux4_1
X_32784_ _32914_/CLK _32784_/D VGND VGND VPWR VPWR _32784_/Q sky130_fd_sc_hd__dfxtp_1
X_35572_ _35699_/CLK _35572_/D VGND VGND VPWR VPWR _35572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34523_ _35544_/CLK _34523_/D VGND VGND VPWR VPWR _34523_/Q sky130_fd_sc_hd__dfxtp_1
X_31735_ _31735_/A VGND VGND VPWR VPWR _36075_/D sky130_fd_sc_hd__clkbuf_1
X_19457_ _19453_/X _19454_/X _19455_/X _19456_/X VGND VGND VPWR VPWR _19457_/X sky130_fd_sc_hd__a22o_1
X_16669_ _16493_/X _16667_/X _16668_/X _16498_/X VGND VGND VPWR VPWR _16669_/X sky130_fd_sc_hd__a22o_1
X_18408_ _33623_/Q _33559_/Q _33495_/Q _33431_/Q _18284_/X _18287_/X VGND VGND VPWR
+ VPWR _18408_/X sky130_fd_sc_hd__mux4_1
X_34454_ _34647_/CLK _34454_/D VGND VGND VPWR VPWR _34454_/Q sky130_fd_sc_hd__dfxtp_1
X_31666_ _27807_/X _36043_/Q _31678_/S VGND VGND VPWR VPWR _31667_/A sky130_fd_sc_hd__mux2_1
X_19388_ _19105_/X _19386_/X _19387_/X _19110_/X VGND VGND VPWR VPWR _19388_/X sky130_fd_sc_hd__a22o_1
XFILLER_210_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18339_ _20134_/A VGND VGND VPWR VPWR _18339_/X sky130_fd_sc_hd__buf_4
X_30617_ _35546_/Q _29342_/X _30627_/S VGND VGND VPWR VPWR _30618_/A sky130_fd_sc_hd__mux2_1
X_33405_ _36092_/CLK _33405_/D VGND VGND VPWR VPWR _33405_/Q sky130_fd_sc_hd__dfxtp_1
X_34385_ _35664_/CLK _34385_/D VGND VGND VPWR VPWR _34385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31597_ _27704_/X _36010_/Q _31615_/S VGND VGND VPWR VPWR _31598_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_1107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36124_ _36235_/CLK _36124_/D VGND VGND VPWR VPWR _36124_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33336_ _36090_/CLK _33336_/D VGND VGND VPWR VPWR _33336_/Q sky130_fd_sc_hd__dfxtp_1
X_21350_ _21306_/X _21348_/X _21349_/X _21312_/X VGND VGND VPWR VPWR _21350_/X sky130_fd_sc_hd__a22o_1
X_30548_ _30548_/A VGND VGND VPWR VPWR _35513_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20301_ _35212_/Q _35148_/Q _35084_/Q _32268_/Q _20016_/X _20017_/X VGND VGND VPWR
+ VPWR _20301_/X sky130_fd_sc_hd__mux4_1
X_36055_ _36055_/CLK _36055_/D VGND VGND VPWR VPWR _36055_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33267_ _33393_/CLK _33267_/D VGND VGND VPWR VPWR _33267_/Q sky130_fd_sc_hd__dfxtp_1
X_21281_ _20961_/X _21279_/X _21280_/X _20965_/X VGND VGND VPWR VPWR _21281_/X sky130_fd_sc_hd__a22o_1
X_30479_ _30479_/A VGND VGND VPWR VPWR _35480_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_951 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23020_ _23020_/A VGND VGND VPWR VPWR _32064_/D sky130_fd_sc_hd__clkbuf_1
X_20232_ _34698_/Q _34634_/Q _34570_/Q _34506_/Q _19945_/X _19946_/X VGND VGND VPWR
+ VPWR _20232_/X sky130_fd_sc_hd__mux4_1
XFILLER_200_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35006_ _35777_/CLK _35006_/D VGND VGND VPWR VPWR _35006_/Q sky130_fd_sc_hd__dfxtp_1
X_32218_ _35709_/CLK _32218_/D VGND VGND VPWR VPWR _32218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33198_ _36079_/CLK _33198_/D VGND VGND VPWR VPWR _33198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20163_ _20159_/X _20160_/X _20161_/X _20162_/X VGND VGND VPWR VPWR _20163_/X sky130_fd_sc_hd__a22o_1
X_32149_ _35986_/CLK _32149_/D VGND VGND VPWR VPWR _32149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20094_ _19811_/X _20092_/X _20093_/X _19816_/X VGND VGND VPWR VPWR _20094_/X sky130_fd_sc_hd__a22o_1
X_24971_ _24970_/X _32973_/Q _24983_/S VGND VGND VPWR VPWR _24972_/A sky130_fd_sc_hd__mux2_1
XTAP_4307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_285_CLK clkbuf_6_58__f_CLK/X VGND VGND VPWR VPWR _36095_/CLK sky130_fd_sc_hd__clkbuf_16
X_26710_ _26710_/A VGND VGND VPWR VPWR _33788_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35908_ _35973_/CLK _35908_/D VGND VGND VPWR VPWR _35908_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23922_ _23922_/A VGND VGND VPWR VPWR _32506_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27690_ _27689_/X _34213_/Q _27702_/S VGND VGND VPWR VPWR _27691_/A sky130_fd_sc_hd__mux2_1
XTAP_3606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26641_ _26641_/A VGND VGND VPWR VPWR _33755_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23853_ _23853_/A VGND VGND VPWR VPWR _32473_/D sky130_fd_sc_hd__clkbuf_1
X_35839_ _35839_/CLK _35839_/D VGND VGND VPWR VPWR _35839_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22804_ _35667_/Q _35027_/Q _34387_/Q _33747_/Q _20712_/X _20713_/X VGND VGND VPWR
+ VPWR _22804_/X sky130_fd_sc_hd__mux4_1
X_29360_ input2/X VGND VGND VPWR VPWR _29360_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_232_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26572_ _24920_/X _33725_/Q _26572_/S VGND VGND VPWR VPWR _26573_/A sky130_fd_sc_hd__mux2_1
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20996_ _33119_/Q _35999_/Q _32991_/Q _32927_/Q _20956_/X _20957_/X VGND VGND VPWR
+ VPWR _20996_/X sky130_fd_sc_hd__mux4_1
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23784_ _22999_/X _32378_/Q _23790_/S VGND VGND VPWR VPWR _23785_/A sky130_fd_sc_hd__mux2_1
X_28311_ _28311_/A VGND VGND VPWR VPWR _34484_/D sky130_fd_sc_hd__clkbuf_1
X_25523_ _25523_/A VGND VGND VPWR VPWR _33228_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_225_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22735_ _22731_/X _22734_/X _22438_/X VGND VGND VPWR VPWR _22757_/A sky130_fd_sc_hd__o21ba_1
XFILLER_214_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29291_ _34948_/Q _27177_/X _29297_/S VGND VGND VPWR VPWR _29292_/A sky130_fd_sc_hd__mux2_1
XFILLER_197_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28242_ _28242_/A VGND VGND VPWR VPWR _34452_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1067 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25454_ _25454_/A VGND VGND VPWR VPWR _33195_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22666_ _22662_/X _22665_/X _22471_/X VGND VGND VPWR VPWR _22667_/D sky130_fd_sc_hd__o21ba_1
XFILLER_200_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24405_ _22906_/X _32732_/Q _24411_/S VGND VGND VPWR VPWR _24406_/A sky130_fd_sc_hd__mux2_1
XFILLER_205_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21617_ _21613_/X _21616_/X _21412_/X VGND VGND VPWR VPWR _21618_/D sky130_fd_sc_hd__o21ba_1
X_28173_ _28173_/A VGND VGND VPWR VPWR _34419_/D sky130_fd_sc_hd__clkbuf_1
X_25385_ _33164_/Q _23469_/X _25395_/S VGND VGND VPWR VPWR _25386_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22597_ _22593_/X _22596_/X _22457_/X VGND VGND VPWR VPWR _22607_/C sky130_fd_sc_hd__o21ba_1
XFILLER_90_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27124_ input22/X VGND VGND VPWR VPWR _27124_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_103_1327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24336_ _24336_/A VGND VGND VPWR VPWR _32699_/D sky130_fd_sc_hd__clkbuf_1
X_21548_ _21548_/A _21548_/B _21548_/C _21548_/D VGND VGND VPWR VPWR _21549_/A sky130_fd_sc_hd__or4_4
XFILLER_217_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27055_ _27055_/A VGND VGND VPWR VPWR _33948_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24267_ _24267_/A VGND VGND VPWR VPWR _32666_/D sky130_fd_sc_hd__clkbuf_1
X_21479_ _34924_/Q _34860_/Q _34796_/Q _34732_/Q _21407_/X _21408_/X VGND VGND VPWR
+ VPWR _21479_/X sky130_fd_sc_hd__mux4_1
XFILLER_101_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26006_ _26006_/A VGND VGND VPWR VPWR _33457_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23218_ _23218_/A VGND VGND VPWR VPWR _32146_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24198_ _24198_/A VGND VGND VPWR VPWR _32635_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23149_ _23149_/A VGND VGND VPWR VPWR _32113_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_1300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27957_ _27813_/X _34317_/Q _27965_/S VGND VGND VPWR VPWR _27958_/A sky130_fd_sc_hd__mux2_1
XTAP_5520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_276_CLK clkbuf_6_59__f_CLK/X VGND VGND VPWR VPWR _36100_/CLK sky130_fd_sc_hd__clkbuf_16
X_17710_ _35460_/Q _35396_/Q _35332_/Q _35268_/Q _17607_/X _17608_/X VGND VGND VPWR
+ VPWR _17710_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_721 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26908_ _33882_/Q _23243_/X _26918_/S VGND VGND VPWR VPWR _26909_/A sky130_fd_sc_hd__mux2_1
XTAP_5564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18690_ _18440_/X _18686_/X _18689_/X _18445_/X VGND VGND VPWR VPWR _18690_/X sky130_fd_sc_hd__a22o_1
XFILLER_29_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27888_ _27711_/X _34284_/Q _27902_/S VGND VGND VPWR VPWR _27889_/A sky130_fd_sc_hd__mux2_1
XTAP_5586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17641_ _35458_/Q _35394_/Q _35330_/Q _35266_/Q _17607_/X _17608_/X VGND VGND VPWR
+ VPWR _17641_/X sky130_fd_sc_hd__mux4_1
XTAP_4852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29627_ _35077_/Q _29475_/X _29631_/S VGND VGND VPWR VPWR _29628_/A sky130_fd_sc_hd__mux2_1
XTAP_4863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26839_ _26839_/A VGND VGND VPWR VPWR _33849_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17572_ _35712_/Q _32222_/Q _35584_/Q _35520_/Q _17317_/X _17318_/X VGND VGND VPWR
+ VPWR _17572_/X sky130_fd_sc_hd__mux4_1
X_29558_ _35044_/Q _29373_/X _29568_/S VGND VGND VPWR VPWR _29559_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19311_ _19311_/A VGND VGND VPWR VPWR _19311_/X sky130_fd_sc_hd__clkbuf_4
X_28509_ _27831_/X _34579_/Q _28513_/S VGND VGND VPWR VPWR _28510_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16523_ _17716_/A VGND VGND VPWR VPWR _16523_/X sky130_fd_sc_hd__buf_6
XFILLER_232_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29489_ _35017_/Q _29488_/X _29513_/S VGND VGND VPWR VPWR _29490_/A sky130_fd_sc_hd__mux2_1
XFILLER_225_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31520_ _27791_/X _35974_/Q _31522_/S VGND VGND VPWR VPWR _31521_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_846 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19242_ _35182_/Q _35118_/Q _35054_/Q _32174_/Q _18957_/X _18958_/X VGND VGND VPWR
+ VPWR _19242_/X sky130_fd_sc_hd__mux4_1
XFILLER_220_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16454_ _17866_/A VGND VGND VPWR VPWR _16454_/X sky130_fd_sc_hd__buf_4
XFILLER_232_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_936 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19173_ _34668_/Q _34604_/Q _34540_/Q _34476_/Q _18886_/X _18887_/X VGND VGND VPWR
+ VPWR _19173_/X sky130_fd_sc_hd__mux4_1
X_31451_ _27689_/X _35941_/Q _31459_/S VGND VGND VPWR VPWR _31452_/A sky130_fd_sc_hd__mux2_1
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16385_ _16385_/A VGND VGND VPWR VPWR _31966_/D sky130_fd_sc_hd__clkbuf_1
XPHY_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_200_CLK clkbuf_6_49__f_CLK/X VGND VGND VPWR VPWR _35849_/CLK sky130_fd_sc_hd__clkbuf_16
X_18124_ _34960_/Q _34896_/Q _34832_/Q _34768_/Q _17866_/X _17867_/X VGND VGND VPWR
+ VPWR _18124_/X sky130_fd_sc_hd__mux4_1
XFILLER_129_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30402_ _35444_/Q _29422_/X _30420_/S VGND VGND VPWR VPWR _30403_/A sky130_fd_sc_hd__mux2_1
X_34170_ _35320_/CLK _34170_/D VGND VGND VPWR VPWR _34170_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31382_ _31382_/A VGND VGND VPWR VPWR _35908_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33121_ _36002_/CLK _33121_/D VGND VGND VPWR VPWR _33121_/Q sky130_fd_sc_hd__dfxtp_1
X_18055_ _15981_/X _18053_/X _18054_/X _15991_/X VGND VGND VPWR VPWR _18055_/X sky130_fd_sc_hd__a22o_1
X_30333_ _35412_/Q _29521_/X _30335_/S VGND VGND VPWR VPWR _30334_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17006_ _17869_/A VGND VGND VPWR VPWR _17006_/X sky130_fd_sc_hd__clkbuf_4
X_33052_ _35804_/CLK _33052_/D VGND VGND VPWR VPWR _33052_/Q sky130_fd_sc_hd__dfxtp_1
X_30264_ _35379_/Q _29419_/X _30264_/S VGND VGND VPWR VPWR _30265_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32003_ _36207_/CLK _32003_/D VGND VGND VPWR VPWR _32003_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_634 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30195_ _30195_/A VGND VGND VPWR VPWR _35346_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18957_ _20016_/A VGND VGND VPWR VPWR _18957_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_86_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_267_CLK clkbuf_6_60__f_CLK/X VGND VGND VPWR VPWR _34690_/CLK sky130_fd_sc_hd__clkbuf_16
X_17908_ _33674_/Q _33610_/Q _33546_/Q _33482_/Q _17906_/X _17907_/X VGND VGND VPWR
+ VPWR _17908_/X sky130_fd_sc_hd__mux4_1
XFILLER_230_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33954_ _34085_/CLK _33954_/D VGND VGND VPWR VPWR _33954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18888_ _34660_/Q _34596_/Q _34532_/Q _34468_/Q _18886_/X _18887_/X VGND VGND VPWR
+ VPWR _18888_/X sky130_fd_sc_hd__mux4_1
XFILLER_55_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32905_ _32905_/CLK _32905_/D VGND VGND VPWR VPWR _32905_/Q sky130_fd_sc_hd__dfxtp_1
X_17839_ _17832_/X _17837_/X _17838_/X VGND VGND VPWR VPWR _17873_/A sky130_fd_sc_hd__o21ba_2
XFILLER_27_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33885_ _35551_/CLK _33885_/D VGND VGND VPWR VPWR _33885_/Q sky130_fd_sc_hd__dfxtp_1
X_20850_ _20846_/X _20849_/X _20615_/X VGND VGND VPWR VPWR _20874_/A sky130_fd_sc_hd__o21ba_1
X_35624_ _35624_/CLK _35624_/D VGND VGND VPWR VPWR _35624_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32836_ _32901_/CLK _32836_/D VGND VGND VPWR VPWR _32836_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19509_ _20215_/A VGND VGND VPWR VPWR _19509_/X sky130_fd_sc_hd__buf_6
XFILLER_179_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20781_ _33369_/Q _33305_/Q _33241_/Q _33177_/Q _20602_/X _20603_/X VGND VGND VPWR
+ VPWR _20781_/X sky130_fd_sc_hd__mux4_1
XFILLER_34_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35555_ _36135_/CLK _35555_/D VGND VGND VPWR VPWR _35555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32767_ _32896_/CLK _32767_/D VGND VGND VPWR VPWR _32767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34506_ _34698_/CLK _34506_/D VGND VGND VPWR VPWR _34506_/Q sky130_fd_sc_hd__dfxtp_1
X_22520_ _22365_/X _22518_/X _22519_/X _22371_/X VGND VGND VPWR VPWR _22520_/X sky130_fd_sc_hd__a22o_1
XFILLER_74_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31718_ _31718_/A VGND VGND VPWR VPWR _36067_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35486_ _35551_/CLK _35486_/D VGND VGND VPWR VPWR _35486_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32698_ _32890_/CLK _32698_/D VGND VGND VPWR VPWR _32698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_241_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34437_ _36164_/CLK _34437_/D VGND VGND VPWR VPWR _34437_/Q sky130_fd_sc_hd__dfxtp_1
X_22451_ _22451_/A VGND VGND VPWR VPWR _22451_/X sky130_fd_sc_hd__clkbuf_4
X_31649_ _27782_/X _36035_/Q _31657_/S VGND VGND VPWR VPWR _31650_/A sky130_fd_sc_hd__mux2_1
XFILLER_206_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21402_ _35178_/Q _35114_/Q _35050_/Q _32170_/Q _21257_/X _21258_/X VGND VGND VPWR
+ VPWR _21402_/X sky130_fd_sc_hd__mux4_1
XFILLER_182_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22382_ _22304_/X _22380_/X _22381_/X _22307_/X VGND VGND VPWR VPWR _22382_/X sky130_fd_sc_hd__a22o_1
X_25170_ _25170_/A VGND VGND VPWR VPWR _33062_/D sky130_fd_sc_hd__clkbuf_1
X_34368_ _35777_/CLK _34368_/D VGND VGND VPWR VPWR _34368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36107_ _36109_/CLK _36107_/D VGND VGND VPWR VPWR _36107_/Q sky130_fd_sc_hd__dfxtp_1
X_24121_ _24121_/A VGND VGND VPWR VPWR _32598_/D sky130_fd_sc_hd__clkbuf_1
X_21333_ _34408_/Q _36136_/Q _34280_/Q _34216_/Q _21123_/X _21124_/X VGND VGND VPWR
+ VPWR _21333_/X sky130_fd_sc_hd__mux4_1
XFILLER_159_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33319_ _36072_/CLK _33319_/D VGND VGND VPWR VPWR _33319_/Q sky130_fd_sc_hd__dfxtp_1
X_34299_ _36154_/CLK _34299_/D VGND VGND VPWR VPWR _34299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36038_ _36038_/CLK _36038_/D VGND VGND VPWR VPWR _36038_/Q sky130_fd_sc_hd__dfxtp_1
X_21264_ _21260_/X _21263_/X _21059_/X VGND VGND VPWR VPWR _21265_/D sky130_fd_sc_hd__o21ba_1
X_24052_ _24052_/A VGND VGND VPWR VPWR _32567_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_176_1450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20215_ _20215_/A VGND VGND VPWR VPWR _20215_/X sky130_fd_sc_hd__buf_4
X_23003_ _23002_/X _32059_/Q _23009_/S VGND VGND VPWR VPWR _23004_/A sky130_fd_sc_hd__mux2_1
X_28860_ _28860_/A VGND VGND VPWR VPWR _34743_/D sky130_fd_sc_hd__clkbuf_1
X_21195_ _21195_/A _21195_/B _21195_/C _21195_/D VGND VGND VPWR VPWR _21196_/A sky130_fd_sc_hd__or4_2
XFILLER_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27811_ _27810_/X _34252_/Q _27826_/S VGND VGND VPWR VPWR _27812_/A sky130_fd_sc_hd__mux2_1
X_20146_ _20146_/A VGND VGND VPWR VPWR _20146_/X sky130_fd_sc_hd__buf_2
X_28791_ _28791_/A VGND VGND VPWR VPWR _34710_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_258_CLK clkbuf_6_63__f_CLK/X VGND VGND VPWR VPWR _36161_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_83_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27742_ input26/X VGND VGND VPWR VPWR _27742_/X sky130_fd_sc_hd__buf_2
XFILLER_106_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24954_ input46/X VGND VGND VPWR VPWR _24954_/X sky130_fd_sc_hd__buf_4
X_20077_ _20077_/A VGND VGND VPWR VPWR _20077_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_170_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_6_27__f_CLK clkbuf_5_13_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_27__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XTAP_4148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_1388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23905_ _23905_/A VGND VGND VPWR VPWR _32498_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27673_ input2/X VGND VGND VPWR VPWR _27673_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24885_ _24885_/A VGND VGND VPWR VPWR _32945_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29412_ _29412_/A VGND VGND VPWR VPWR _34992_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26624_ _27232_/A _28786_/B VGND VGND VPWR VPWR _26625_/A sky130_fd_sc_hd__or2_1
XFILLER_17_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23836_ _23076_/X _32403_/Q _23840_/S VGND VGND VPWR VPWR _23837_/A sky130_fd_sc_hd__mux2_1
XTAP_3469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29343_ _34970_/Q _29342_/X _29358_/S VGND VGND VPWR VPWR _29344_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26555_ _26555_/A VGND VGND VPWR VPWR _33716_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23767_ _22974_/X _32370_/Q _23769_/S VGND VGND VPWR VPWR _23768_/A sky130_fd_sc_hd__mux2_1
XFILLER_214_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20979_ _20678_/X _20977_/X _20978_/X _20688_/X VGND VGND VPWR VPWR _20979_/X sky130_fd_sc_hd__a22o_1
XFILLER_202_903 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_430_CLK clkbuf_6_38__f_CLK/X VGND VGND VPWR VPWR _35187_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_82_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25506_ _25506_/A VGND VGND VPWR VPWR _33220_/D sky130_fd_sc_hd__clkbuf_1
X_22718_ _20601_/X _22716_/X _22717_/X _20607_/X VGND VGND VPWR VPWR _22718_/X sky130_fd_sc_hd__a22o_1
X_29274_ _34940_/Q _27152_/X _29276_/S VGND VGND VPWR VPWR _29275_/A sky130_fd_sc_hd__mux2_1
XFILLER_246_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26486_ _33685_/Q _23498_/X _26486_/S VGND VGND VPWR VPWR _26487_/A sky130_fd_sc_hd__mux2_1
X_23698_ _23076_/X _32339_/Q _23702_/S VGND VGND VPWR VPWR _23699_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28225_ _27810_/X _34444_/Q _28235_/S VGND VGND VPWR VPWR _28226_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25437_ _25437_/A VGND VGND VPWR VPWR _33187_/D sky130_fd_sc_hd__clkbuf_1
X_22649_ _32142_/Q _32334_/Q _32398_/Q _35918_/Q _22586_/X _22374_/X VGND VGND VPWR
+ VPWR _22649_/X sky130_fd_sc_hd__mux4_1
XFILLER_40_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16170_ _17716_/A VGND VGND VPWR VPWR _16170_/X sky130_fd_sc_hd__buf_6
X_28156_ _27708_/X _34411_/Q _28172_/S VGND VGND VPWR VPWR _28157_/A sky130_fd_sc_hd__mux2_1
X_25368_ _33156_/Q _23441_/X _25374_/S VGND VGND VPWR VPWR _25369_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_586 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27107_ _33965_/Q _27106_/X _27125_/S VGND VGND VPWR VPWR _27108_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24319_ _24319_/A VGND VGND VPWR VPWR _32691_/D sky130_fd_sc_hd__clkbuf_1
X_28087_ _28087_/A VGND VGND VPWR VPWR _34378_/D sky130_fd_sc_hd__clkbuf_1
X_25299_ _33123_/Q _23271_/X _25311_/S VGND VGND VPWR VPWR _25300_/A sky130_fd_sc_hd__mux2_1
X_27038_ input12/X VGND VGND VPWR VPWR _27038_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_99_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_1403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_497_CLK clkbuf_6_2__f_CLK/X VGND VGND VPWR VPWR _35622_/CLK sky130_fd_sc_hd__clkbuf_16
X_19860_ _33408_/Q _33344_/Q _33280_/Q _33216_/Q _19780_/X _19781_/X VGND VGND VPWR
+ VPWR _19860_/X sky130_fd_sc_hd__mux4_1
XFILLER_107_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18811_ _18661_/X _18809_/X _18810_/X _18665_/X VGND VGND VPWR VPWR _18811_/X sky130_fd_sc_hd__a22o_1
XTAP_6040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19791_ _32894_/Q _32830_/Q _32766_/Q _32702_/Q _19646_/X _19647_/X VGND VGND VPWR
+ VPWR _19791_/X sky130_fd_sc_hd__mux4_1
Xoutput94 _31971_/Q VGND VGND VPWR VPWR D1[13] sky130_fd_sc_hd__buf_2
XTAP_6062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28989_ _28989_/A VGND VGND VPWR VPWR _34804_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_249_CLK clkbuf_6_61__f_CLK/X VGND VGND VPWR VPWR _33673_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_6073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18742_ _35424_/Q _35360_/Q _35296_/Q _35232_/Q _18495_/X _18496_/X VGND VGND VPWR
+ VPWR _18742_/X sky130_fd_sc_hd__mux4_1
XTAP_6095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30951_ _30951_/A VGND VGND VPWR VPWR _35704_/D sky130_fd_sc_hd__clkbuf_1
X_18673_ _20236_/A VGND VGND VPWR VPWR _18673_/X sky130_fd_sc_hd__buf_4
XTAP_4660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17624_ _17552_/X _17622_/X _17623_/X _17557_/X VGND VGND VPWR VPWR _17624_/X sky130_fd_sc_hd__a22o_1
XTAP_4693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33670_ _34182_/CLK _33670_/D VGND VGND VPWR VPWR _33670_/Q sky130_fd_sc_hd__dfxtp_1
X_30882_ _30882_/A VGND VGND VPWR VPWR _35671_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17555_ _33664_/Q _33600_/Q _33536_/Q _33472_/Q _17553_/X _17554_/X VGND VGND VPWR
+ VPWR _17555_/X sky130_fd_sc_hd__mux4_1
XTAP_3992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32621_ _36013_/CLK _32621_/D VGND VGND VPWR VPWR _32621_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16506_ _32610_/Q _32546_/Q _32482_/Q _35938_/Q _16217_/X _16354_/X VGND VGND VPWR
+ VPWR _16506_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_421_CLK clkbuf_6_33__f_CLK/X VGND VGND VPWR VPWR _35056_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_232_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35340_ _35471_/CLK _35340_/D VGND VGND VPWR VPWR _35340_/Q sky130_fd_sc_hd__dfxtp_1
X_32552_ _32552_/CLK _32552_/D VGND VGND VPWR VPWR _32552_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17486_ _17479_/X _17484_/X _17485_/X VGND VGND VPWR VPWR _17520_/A sky130_fd_sc_hd__o21ba_1
XFILLER_108_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31503_ _31551_/S VGND VGND VPWR VPWR _31522_/S sky130_fd_sc_hd__buf_4
X_16437_ _35680_/Q _32186_/Q _35552_/Q _35488_/Q _16258_/X _16259_/X VGND VGND VPWR
+ VPWR _16437_/X sky130_fd_sc_hd__mux4_1
X_19225_ _33134_/Q _36014_/Q _33006_/Q _32942_/Q _19009_/X _19010_/X VGND VGND VPWR
+ VPWR _19225_/X sky130_fd_sc_hd__mux4_1
XFILLER_220_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35271_ _35845_/CLK _35271_/D VGND VGND VPWR VPWR _35271_/Q sky130_fd_sc_hd__dfxtp_1
X_32483_ _35938_/CLK _32483_/D VGND VGND VPWR VPWR _32483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31434_ _27664_/X _35933_/Q _31438_/S VGND VGND VPWR VPWR _31435_/A sky130_fd_sc_hd__mux2_1
X_19156_ _20215_/A VGND VGND VPWR VPWR _19156_/X sky130_fd_sc_hd__clkbuf_4
X_34222_ _36142_/CLK _34222_/D VGND VGND VPWR VPWR _34222_/Q sky130_fd_sc_hd__dfxtp_1
X_16368_ _35678_/Q _32184_/Q _35550_/Q _35486_/Q _16258_/X _16259_/X VGND VGND VPWR
+ VPWR _16368_/X sky130_fd_sc_hd__mux4_1
XFILLER_157_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_1287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18107_ _33168_/Q _36048_/Q _33040_/Q _32976_/Q _16032_/X _17161_/A VGND VGND VPWR
+ VPWR _18107_/X sky130_fd_sc_hd__mux4_1
XFILLER_157_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34153_ _34153_/CLK _34153_/D VGND VGND VPWR VPWR _34153_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19087_ _20146_/A VGND VGND VPWR VPWR _19087_/X sky130_fd_sc_hd__clkbuf_4
X_31365_ _31365_/A VGND VGND VPWR VPWR _35900_/D sky130_fd_sc_hd__clkbuf_1
X_16299_ _33052_/Q _32028_/Q _35804_/Q _35740_/Q _16067_/X _16069_/X VGND VGND VPWR
+ VPWR _16299_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30316_ _30316_/A VGND VGND VPWR VPWR _35403_/D sky130_fd_sc_hd__clkbuf_1
X_33104_ _35855_/CLK _33104_/D VGND VGND VPWR VPWR _33104_/Q sky130_fd_sc_hd__dfxtp_1
X_18038_ _18038_/A VGND VGND VPWR VPWR _32013_/D sky130_fd_sc_hd__buf_2
X_34084_ _34148_/CLK _34084_/D VGND VGND VPWR VPWR _34084_/Q sky130_fd_sc_hd__dfxtp_1
X_31296_ _31296_/A VGND VGND VPWR VPWR _35867_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_488_CLK _35560_/CLK VGND VGND VPWR VPWR _34987_/CLK sky130_fd_sc_hd__clkbuf_16
X_33035_ _36044_/CLK _33035_/D VGND VGND VPWR VPWR _33035_/Q sky130_fd_sc_hd__dfxtp_1
X_30247_ _30247_/A VGND VGND VPWR VPWR _35370_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_1191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20000_ _20134_/A VGND VGND VPWR VPWR _20000_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_119_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30178_ _35338_/Q _29491_/X _30192_/S VGND VGND VPWR VPWR _30179_/A sky130_fd_sc_hd__mux2_1
X_19989_ _34180_/Q _34116_/Q _34052_/Q _33988_/Q _19746_/X _19747_/X VGND VGND VPWR
+ VPWR _19989_/X sky130_fd_sc_hd__mux4_1
XFILLER_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34986_ _35690_/CLK _34986_/D VGND VGND VPWR VPWR _34986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_223_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33937_ _34440_/CLK _33937_/D VGND VGND VPWR VPWR _33937_/Q sky130_fd_sc_hd__dfxtp_1
X_21951_ _22459_/A VGND VGND VPWR VPWR _21951_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_55_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20902_ _20896_/X _20901_/X _20675_/X VGND VGND VPWR VPWR _20912_/C sky130_fd_sc_hd__o21ba_1
XFILLER_243_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24670_ _24670_/A VGND VGND VPWR VPWR _32857_/D sky130_fd_sc_hd__clkbuf_1
X_33868_ _33934_/CLK _33868_/D VGND VGND VPWR VPWR _33868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21882_ _32888_/Q _32824_/Q _32760_/Q _32696_/Q _21593_/X _21594_/X VGND VGND VPWR
+ VPWR _21882_/X sky130_fd_sc_hd__mux4_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35607_ _35801_/CLK _35607_/D VGND VGND VPWR VPWR _35607_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23621_ _22962_/X _32302_/Q _23631_/S VGND VGND VPWR VPWR _23622_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20833_ _22598_/A VGND VGND VPWR VPWR _20833_/X sky130_fd_sc_hd__buf_6
X_32819_ _32906_/CLK _32819_/D VGND VGND VPWR VPWR _32819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33799_ _36159_/CLK _33799_/D VGND VGND VPWR VPWR _33799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_412_CLK clkbuf_6_32__f_CLK/X VGND VGND VPWR VPWR _33904_/CLK sky130_fd_sc_hd__clkbuf_16
X_26340_ _24979_/X _33616_/Q _26342_/S VGND VGND VPWR VPWR _26341_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23552_ _23552_/A VGND VGND VPWR VPWR _32270_/D sky130_fd_sc_hd__clkbuf_1
X_35538_ _35730_/CLK _35538_/D VGND VGND VPWR VPWR _35538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20764_ _33048_/Q _32024_/Q _35800_/Q _35736_/Q _20667_/X _20669_/X VGND VGND VPWR
+ VPWR _20764_/X sky130_fd_sc_hd__mux4_1
XFILLER_208_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22503_ _22503_/A _22503_/B _22503_/C _22503_/D VGND VGND VPWR VPWR _22504_/A sky130_fd_sc_hd__or4_4
XFILLER_196_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26271_ _24877_/X _33583_/Q _26279_/S VGND VGND VPWR VPWR _26272_/A sky130_fd_sc_hd__mux2_1
X_20695_ _34390_/Q _36118_/Q _34262_/Q _34198_/Q _20692_/X _20694_/X VGND VGND VPWR
+ VPWR _20695_/X sky130_fd_sc_hd__mux4_1
XFILLER_210_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23483_ _23483_/A VGND VGND VPWR VPWR _32239_/D sky130_fd_sc_hd__clkbuf_1
X_35469_ _35471_/CLK _35469_/D VGND VGND VPWR VPWR _35469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28010_ _34342_/Q _27084_/X _28016_/S VGND VGND VPWR VPWR _28011_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25222_ _33087_/Q _23426_/X _25238_/S VGND VGND VPWR VPWR _25223_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22434_ _22434_/A VGND VGND VPWR VPWR _22434_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_10_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_5_17_0_CLK clkbuf_2_2_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_17_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_13_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25153_ _25153_/A VGND VGND VPWR VPWR _33054_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22365_ _22365_/A VGND VGND VPWR VPWR _22365_/X sky130_fd_sc_hd__clkbuf_4
X_24104_ _24104_/A VGND VGND VPWR VPWR _32592_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21316_ _32104_/Q _32296_/Q _32360_/Q _35880_/Q _21174_/X _21315_/X VGND VGND VPWR
+ VPWR _21316_/X sky130_fd_sc_hd__mux4_1
X_22296_ _33156_/Q _36036_/Q _33028_/Q _32964_/Q _22015_/X _22016_/X VGND VGND VPWR
+ VPWR _22296_/X sky130_fd_sc_hd__mux4_1
X_25084_ _25084_/A VGND VGND VPWR VPWR _33022_/D sky130_fd_sc_hd__clkbuf_1
X_29961_ _35235_/Q _29370_/X _29973_/S VGND VGND VPWR VPWR _29962_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_479_CLK clkbuf_6_10__f_CLK/X VGND VGND VPWR VPWR _34093_/CLK sky130_fd_sc_hd__clkbuf_16
X_28912_ _28912_/A VGND VGND VPWR VPWR _34768_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21247_ _35622_/Q _34982_/Q _34342_/Q _33702_/Q _21038_/X _21039_/X VGND VGND VPWR
+ VPWR _21247_/X sky130_fd_sc_hd__mux4_1
X_24035_ _24035_/A VGND VGND VPWR VPWR _32559_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_176_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29892_ _29892_/A VGND VGND VPWR VPWR _35202_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28843_ _28843_/A VGND VGND VPWR VPWR _34735_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21178_ _21173_/X _21177_/X _21034_/X _21035_/X VGND VGND VPWR VPWR _21195_/B sky130_fd_sc_hd__o211a_1
XFILLER_89_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20129_ _20129_/A VGND VGND VPWR VPWR _32455_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28774_ _34704_/Q _27214_/X _28776_/S VGND VGND VPWR VPWR _28775_/A sky130_fd_sc_hd__mux2_1
XFILLER_237_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25986_ _24855_/X _33448_/Q _25988_/S VGND VGND VPWR VPWR _25987_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27725_ _27725_/A VGND VGND VPWR VPWR _34224_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24937_ _24936_/X _32962_/Q _24952_/S VGND VGND VPWR VPWR _24938_/A sky130_fd_sc_hd__mux2_1
XTAP_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27656_ _27655_/X _34202_/Q _27671_/S VGND VGND VPWR VPWR _27657_/A sky130_fd_sc_hd__mux2_1
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24868_ input15/X VGND VGND VPWR VPWR _24868_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26607_ _26607_/A VGND VGND VPWR VPWR _33741_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23819_ _23819_/A VGND VGND VPWR VPWR _32394_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27587_ _34173_/Q _27155_/X _27587_/S VGND VGND VPWR VPWR _27588_/A sky130_fd_sc_hd__mux2_1
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24799_ _31418_/B _31553_/B VGND VGND VPWR VPWR _24995_/S sky130_fd_sc_hd__nand2_8
XFILLER_26_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_403_CLK clkbuf_6_34__f_CLK/X VGND VGND VPWR VPWR _35701_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29326_ _34965_/Q _27229_/X _29326_/S VGND VGND VPWR VPWR _29327_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17340_ _17206_/X _17338_/X _17339_/X _17209_/X VGND VGND VPWR VPWR _17340_/X sky130_fd_sc_hd__a22o_1
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26538_ _26538_/A VGND VGND VPWR VPWR _33708_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17271_ _17199_/X _17269_/X _17270_/X _17204_/X VGND VGND VPWR VPWR _17271_/X sky130_fd_sc_hd__a22o_1
X_29257_ _29326_/S VGND VGND VPWR VPWR _29276_/S sky130_fd_sc_hd__buf_4
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26469_ _26469_/A VGND VGND VPWR VPWR _33676_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19010_ _20207_/A VGND VGND VPWR VPWR _19010_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_109_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28208_ _27785_/X _34436_/Q _28214_/S VGND VGND VPWR VPWR _28209_/A sky130_fd_sc_hd__mux2_1
X_16222_ _32090_/Q _32282_/Q _32346_/Q _35866_/Q _16221_/X _17867_/A VGND VGND VPWR
+ VPWR _16222_/X sky130_fd_sc_hd__mux4_1
X_29188_ _29188_/A VGND VGND VPWR VPWR _34899_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_1134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16153_ _32600_/Q _32536_/Q _32472_/Q _35928_/Q _17866_/A _17717_/A VGND VGND VPWR
+ VPWR _16153_/X sky130_fd_sc_hd__mux4_1
X_28139_ _27683_/X _34403_/Q _28151_/S VGND VGND VPWR VPWR _28140_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31150_ _27639_/X _35798_/Q _31168_/S VGND VGND VPWR VPWR _31151_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16084_ _17766_/A VGND VGND VPWR VPWR _17011_/A sky130_fd_sc_hd__buf_12
XFILLER_115_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30101_ _30101_/A VGND VGND VPWR VPWR _35301_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19912_ _19906_/X _19911_/X _19804_/X VGND VGND VPWR VPWR _19920_/C sky130_fd_sc_hd__o21ba_1
XFILLER_190_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31081_ _35766_/Q input26/X _31095_/S VGND VGND VPWR VPWR _31082_/A sky130_fd_sc_hd__mux2_1
XFILLER_244_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30032_ _35269_/Q _29475_/X _30036_/S VGND VGND VPWR VPWR _30033_/A sky130_fd_sc_hd__mux2_1
X_19843_ _34687_/Q _34623_/Q _34559_/Q _34495_/Q _19592_/X _19593_/X VGND VGND VPWR
+ VPWR _19843_/X sky130_fd_sc_hd__mux4_1
XFILLER_116_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34840_ _34904_/CLK _34840_/D VGND VGND VPWR VPWR _34840_/Q sky130_fd_sc_hd__dfxtp_1
X_19774_ _19770_/X _19773_/X _19465_/X VGND VGND VPWR VPWR _19775_/D sky130_fd_sc_hd__o21ba_1
XFILLER_84_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16986_ _33904_/Q _33840_/Q _33776_/Q _36080_/Q _16671_/X _16672_/X VGND VGND VPWR
+ VPWR _16986_/X sky130_fd_sc_hd__mux4_1
XFILLER_49_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_871 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18725_ _18447_/X _18723_/X _18724_/X _18450_/X VGND VGND VPWR VPWR _18725_/X sky130_fd_sc_hd__a22o_1
X_34771_ _34964_/CLK _34771_/D VGND VGND VPWR VPWR _34771_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31983_ _34918_/CLK _31983_/D VGND VGND VPWR VPWR _31983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_6_10__f_CLK clkbuf_5_5_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_10__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_33722_ _35197_/CLK _33722_/D VGND VGND VPWR VPWR _33722_/Q sky130_fd_sc_hd__dfxtp_1
X_18656_ _20206_/A VGND VGND VPWR VPWR _18656_/X sky130_fd_sc_hd__buf_4
X_30934_ _30934_/A VGND VGND VPWR VPWR _35696_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17607_ _17960_/A VGND VGND VPWR VPWR _17607_/X sky130_fd_sc_hd__buf_4
XFILLER_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30865_ _35664_/Q input54/X _30867_/S VGND VGND VPWR VPWR _30866_/A sky130_fd_sc_hd__mux2_1
X_33653_ _34101_/CLK _33653_/D VGND VGND VPWR VPWR _33653_/Q sky130_fd_sc_hd__dfxtp_1
X_18587_ _20133_/A VGND VGND VPWR VPWR _18587_/X sky130_fd_sc_hd__buf_4
XFILLER_18_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32604_ _35998_/CLK _32604_/D VGND VGND VPWR VPWR _32604_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17538_ _17351_/X _17536_/X _17537_/X _17354_/X VGND VGND VPWR VPWR _17538_/X sky130_fd_sc_hd__a22o_1
X_33584_ _34035_/CLK _33584_/D VGND VGND VPWR VPWR _33584_/Q sky130_fd_sc_hd__dfxtp_1
X_30796_ _35631_/Q input18/X _30804_/S VGND VGND VPWR VPWR _30797_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35323_ _35451_/CLK _35323_/D VGND VGND VPWR VPWR _35323_/Q sky130_fd_sc_hd__dfxtp_1
X_32535_ _35929_/CLK _32535_/D VGND VGND VPWR VPWR _32535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_968 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17469_ _35197_/Q _35133_/Q _35069_/Q _32253_/Q _17363_/X _17364_/X VGND VGND VPWR
+ VPWR _17469_/X sky130_fd_sc_hd__mux4_1
XFILLER_20_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_242_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19208_ _35181_/Q _35117_/Q _35053_/Q _32173_/Q _18957_/X _18958_/X VGND VGND VPWR
+ VPWR _19208_/X sky130_fd_sc_hd__mux4_1
X_20480_ _34706_/Q _34642_/Q _34578_/Q _34514_/Q _20298_/X _20299_/X VGND VGND VPWR
+ VPWR _20480_/X sky130_fd_sc_hd__mux4_1
XFILLER_165_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35254_ _35765_/CLK _35254_/D VGND VGND VPWR VPWR _35254_/Q sky130_fd_sc_hd__dfxtp_1
X_32466_ _36079_/CLK _32466_/D VGND VGND VPWR VPWR _32466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34205_ _36235_/CLK _34205_/D VGND VGND VPWR VPWR _34205_/Q sky130_fd_sc_hd__dfxtp_1
X_31417_ _31417_/A VGND VGND VPWR VPWR _35925_/D sky130_fd_sc_hd__clkbuf_1
X_19139_ _19100_/X _19137_/X _19138_/X _19103_/X VGND VGND VPWR VPWR _19139_/X sky130_fd_sc_hd__a22o_1
X_32397_ _35916_/CLK _32397_/D VGND VGND VPWR VPWR _32397_/Q sky130_fd_sc_hd__dfxtp_1
X_35185_ _35828_/CLK _35185_/D VGND VGND VPWR VPWR _35185_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22150_ _22150_/A _22150_/B _22150_/C _22150_/D VGND VGND VPWR VPWR _22151_/A sky130_fd_sc_hd__or4_4
X_34136_ _35610_/CLK _34136_/D VGND VGND VPWR VPWR _34136_/Q sky130_fd_sc_hd__dfxtp_1
X_31348_ _27735_/X _35892_/Q _31366_/S VGND VGND VPWR VPWR _31349_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21101_ _33378_/Q _33314_/Q _33250_/Q _33186_/Q _21021_/X _21022_/X VGND VGND VPWR
+ VPWR _21101_/X sky130_fd_sc_hd__mux4_1
XFILLER_218_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22081_ _22434_/A VGND VGND VPWR VPWR _22081_/X sky130_fd_sc_hd__buf_4
X_34067_ _34963_/CLK _34067_/D VGND VGND VPWR VPWR _34067_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31279_ _27834_/X _35860_/Q _31281_/S VGND VGND VPWR VPWR _31280_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21032_ _32864_/Q _32800_/Q _32736_/Q _32672_/Q _20887_/X _20888_/X VGND VGND VPWR
+ VPWR _21032_/X sky130_fd_sc_hd__mux4_1
X_33018_ _36026_/CLK _33018_/D VGND VGND VPWR VPWR _33018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25840_ _25840_/A VGND VGND VPWR VPWR _33378_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25771_ _24936_/X _33346_/Q _25781_/S VGND VGND VPWR VPWR _25772_/A sky130_fd_sc_hd__mux2_1
X_34969_ _35609_/CLK _34969_/D VGND VGND VPWR VPWR _34969_/Q sky130_fd_sc_hd__dfxtp_1
X_22983_ _22983_/A VGND VGND VPWR VPWR _32052_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27510_ _34136_/Q _27041_/X _27524_/S VGND VGND VPWR VPWR _27511_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24722_ _24722_/A VGND VGND VPWR VPWR _32882_/D sky130_fd_sc_hd__clkbuf_1
X_28490_ _28490_/A VGND VGND VPWR VPWR _34569_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21934_ _21934_/A VGND VGND VPWR VPWR _36217_/D sky130_fd_sc_hd__buf_6
XFILLER_103_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27441_ _27441_/A VGND VGND VPWR VPWR _34103_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24653_ _23073_/X _32850_/Q _24659_/S VGND VGND VPWR VPWR _24654_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21865_ _21758_/X _21863_/X _21864_/X _21763_/X VGND VGND VPWR VPWR _21865_/X sky130_fd_sc_hd__a22o_1
XFILLER_93_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23604_ _22937_/X _32294_/Q _23610_/S VGND VGND VPWR VPWR _23605_/A sky130_fd_sc_hd__mux2_1
X_27372_ _27372_/A VGND VGND VPWR VPWR _34070_/D sky130_fd_sc_hd__clkbuf_1
X_20816_ _20812_/X _20815_/X _20615_/X VGND VGND VPWR VPWR _20842_/A sky130_fd_sc_hd__o21ba_1
XFILLER_169_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24584_ _22971_/X _32817_/Q _24588_/S VGND VGND VPWR VPWR _24585_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21796_ _21792_/X _21795_/X _21765_/X VGND VGND VPWR VPWR _21797_/D sky130_fd_sc_hd__o21ba_1
XFILLER_70_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_223_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29111_ _29111_/A VGND VGND VPWR VPWR _34862_/D sky130_fd_sc_hd__clkbuf_1
X_26323_ _26350_/S VGND VGND VPWR VPWR _26342_/S sky130_fd_sc_hd__buf_4
Xclkbuf_5_0_0_CLK clkbuf_5_7_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_0_0_CLK/X sky130_fd_sc_hd__clkbuf_8
X_23535_ _23535_/A VGND VGND VPWR VPWR _32262_/D sky130_fd_sc_hd__clkbuf_1
X_20747_ _22464_/A VGND VGND VPWR VPWR _20747_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_243_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29042_ _34830_/Q _27208_/X _29048_/S VGND VGND VPWR VPWR _29043_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26254_ _24852_/X _33575_/Q _26258_/S VGND VGND VPWR VPWR _26255_/A sky130_fd_sc_hd__mux2_1
X_23466_ input49/X VGND VGND VPWR VPWR _23466_/X sky130_fd_sc_hd__buf_4
XFILLER_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20678_ _21753_/A VGND VGND VPWR VPWR _20678_/X sky130_fd_sc_hd__buf_4
XFILLER_195_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25205_ _33079_/Q _23399_/X _25217_/S VGND VGND VPWR VPWR _25206_/A sky130_fd_sc_hd__mux2_1
X_22417_ _35463_/Q _35399_/Q _35335_/Q _35271_/Q _22207_/X _22208_/X VGND VGND VPWR
+ VPWR _22417_/X sky130_fd_sc_hd__mux4_1
X_26185_ _26185_/A VGND VGND VPWR VPWR _33542_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23397_ _32211_/Q _23396_/X _23418_/S VGND VGND VPWR VPWR _23398_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25136_ _33046_/Q _23225_/X _25154_/S VGND VGND VPWR VPWR _25137_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22348_ _22344_/X _22347_/X _22104_/X VGND VGND VPWR VPWR _22356_/C sky130_fd_sc_hd__o21ba_1
XFILLER_191_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29944_ _35227_/Q _29345_/X _29952_/S VGND VGND VPWR VPWR _29945_/A sky130_fd_sc_hd__mux2_1
X_25067_ _25067_/A VGND VGND VPWR VPWR _33014_/D sky130_fd_sc_hd__clkbuf_1
X_22279_ _34691_/Q _34627_/Q _34563_/Q _34499_/Q _22245_/X _22246_/X VGND VGND VPWR
+ VPWR _22279_/X sky130_fd_sc_hd__mux4_1
XFILLER_219_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24018_ _24018_/A VGND VGND VPWR VPWR _32551_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29875_ _29875_/A VGND VGND VPWR VPWR _35194_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28826_ _28826_/A VGND VGND VPWR VPWR _34727_/D sky130_fd_sc_hd__clkbuf_1
X_16840_ _34411_/Q _36139_/Q _34283_/Q _34219_/Q _16523_/X _16524_/X VGND VGND VPWR
+ VPWR _16840_/X sky130_fd_sc_hd__mux4_1
XFILLER_8_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16771_ _33642_/Q _33578_/Q _33514_/Q _33450_/Q _16494_/X _16495_/X VGND VGND VPWR
+ VPWR _16771_/X sky130_fd_sc_hd__mux4_1
X_28757_ _28784_/S VGND VGND VPWR VPWR _28776_/S sky130_fd_sc_hd__buf_4
XFILLER_150_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25969_ _26080_/S VGND VGND VPWR VPWR _25988_/S sky130_fd_sc_hd__buf_8
XFILLER_24_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18510_ _33626_/Q _33562_/Q _33498_/Q _33434_/Q _18441_/X _18442_/X VGND VGND VPWR
+ VPWR _18510_/X sky130_fd_sc_hd__mux4_1
XFILLER_4_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27708_ input14/X VGND VGND VPWR VPWR _27708_/X sky130_fd_sc_hd__buf_2
XTAP_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19490_ _34677_/Q _34613_/Q _34549_/Q _34485_/Q _19239_/X _19240_/X VGND VGND VPWR
+ VPWR _19490_/X sky130_fd_sc_hd__mux4_1
XTAP_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28688_ _34663_/Q _27087_/X _28692_/S VGND VGND VPWR VPWR _28689_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18441_ _20206_/A VGND VGND VPWR VPWR _18441_/X sky130_fd_sc_hd__buf_6
XFILLER_61_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27639_ input1/X VGND VGND VPWR VPWR _27639_/X sky130_fd_sc_hd__buf_2
XFILLER_46_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18372_ _20169_/A VGND VGND VPWR VPWR _18372_/X sky130_fd_sc_hd__buf_4
X_30650_ _30740_/S VGND VGND VPWR VPWR _30669_/S sky130_fd_sc_hd__buf_4
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_1354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17323_ _33081_/Q _32057_/Q _35833_/Q _35769_/Q _17078_/X _17079_/X VGND VGND VPWR
+ VPWR _17323_/X sky130_fd_sc_hd__mux4_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29309_ _29309_/A VGND VGND VPWR VPWR _34956_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30581_ _35529_/Q _29488_/X _30597_/S VGND VGND VPWR VPWR _30582_/A sky130_fd_sc_hd__mux2_1
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32320_ _35969_/CLK _32320_/D VGND VGND VPWR VPWR _32320_/Q sky130_fd_sc_hd__dfxtp_1
X_17254_ _17960_/A VGND VGND VPWR VPWR _17254_/X sky130_fd_sc_hd__buf_6
XFILLER_202_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16205_ _34905_/Q _34841_/Q _34777_/Q _34713_/Q _16096_/X _16098_/X VGND VGND VPWR
+ VPWR _16205_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32251_ _35194_/CLK _32251_/D VGND VGND VPWR VPWR _32251_/Q sky130_fd_sc_hd__dfxtp_1
X_17185_ _16998_/X _17183_/X _17184_/X _17001_/X VGND VGND VPWR VPWR _17185_/X sky130_fd_sc_hd__a22o_1
XFILLER_155_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31202_ _27720_/X _35823_/Q _31210_/S VGND VGND VPWR VPWR _31203_/A sky130_fd_sc_hd__mux2_1
X_16136_ _16091_/X _16134_/X _16135_/X _16101_/X VGND VGND VPWR VPWR _16136_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32182_ _35547_/CLK _32182_/D VGND VGND VPWR VPWR _32182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31133_ _35791_/Q input53/X _31137_/S VGND VGND VPWR VPWR _31134_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16067_ _17935_/A VGND VGND VPWR VPWR _16067_/X sky130_fd_sc_hd__buf_8
XFILLER_170_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31064_ _35758_/Q input17/X _31074_/S VGND VGND VPWR VPWR _31065_/A sky130_fd_sc_hd__mux2_1
X_35941_ _35941_/CLK _35941_/D VGND VGND VPWR VPWR _35941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30015_ _35261_/Q _29450_/X _30015_/S VGND VGND VPWR VPWR _30016_/A sky130_fd_sc_hd__mux2_1
X_19826_ _33919_/Q _33855_/Q _33791_/Q _36095_/Q _19677_/X _19678_/X VGND VGND VPWR
+ VPWR _19826_/X sky130_fd_sc_hd__mux4_1
X_35872_ _35875_/CLK _35872_/D VGND VGND VPWR VPWR _35872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_819 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34823_ _36113_/CLK _34823_/D VGND VGND VPWR VPWR _34823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19757_ _32125_/Q _32317_/Q _32381_/Q _35901_/Q _19580_/X _19721_/X VGND VGND VPWR
+ VPWR _19757_/X sky130_fd_sc_hd__mux4_1
XFILLER_68_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16969_ _35439_/Q _35375_/Q _35311_/Q _35247_/Q _16901_/X _16902_/X VGND VGND VPWR
+ VPWR _16969_/X sky130_fd_sc_hd__mux4_1
XFILLER_17_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18708_ _18704_/X _18707_/X _18375_/X VGND VGND VPWR VPWR _18716_/C sky130_fd_sc_hd__o21ba_1
X_34754_ _36163_/CLK _34754_/D VGND VGND VPWR VPWR _34754_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31966_ _34148_/CLK _31966_/D VGND VGND VPWR VPWR _31966_/Q sky130_fd_sc_hd__dfxtp_1
X_19688_ _19684_/X _19687_/X _19440_/X _19441_/X VGND VGND VPWR VPWR _19703_/B sky130_fd_sc_hd__o211a_1
XFILLER_25_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33705_ _35625_/CLK _33705_/D VGND VGND VPWR VPWR _33705_/Q sky130_fd_sc_hd__dfxtp_1
X_18639_ _18378_/X _18637_/X _18638_/X _18388_/X VGND VGND VPWR VPWR _18639_/X sky130_fd_sc_hd__a22o_1
X_30917_ _30917_/A VGND VGND VPWR VPWR _35688_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_225_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34685_ _34685_/CLK _34685_/D VGND VGND VPWR VPWR _34685_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31897_ _31897_/A VGND VGND VPWR VPWR _36152_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33636_ _34151_/CLK _33636_/D VGND VGND VPWR VPWR _33636_/Q sky130_fd_sc_hd__dfxtp_1
X_21650_ _21650_/A _21650_/B _21650_/C _21650_/D VGND VGND VPWR VPWR _21651_/A sky130_fd_sc_hd__or4_4
X_30848_ _30875_/S VGND VGND VPWR VPWR _30867_/S sky130_fd_sc_hd__buf_4
XFILLER_36_1102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20601_ _22464_/A VGND VGND VPWR VPWR _20601_/X sky130_fd_sc_hd__clkbuf_4
X_33567_ _36191_/CLK _33567_/D VGND VGND VPWR VPWR _33567_/Q sky130_fd_sc_hd__dfxtp_1
X_21581_ _21581_/A VGND VGND VPWR VPWR _36207_/D sky130_fd_sc_hd__clkbuf_1
X_30779_ _35623_/Q input9/X _30783_/S VGND VGND VPWR VPWR _30780_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23320_ _23320_/A VGND VGND VPWR VPWR _32177_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35306_ _35685_/CLK _35306_/D VGND VGND VPWR VPWR _35306_/Q sky130_fd_sc_hd__dfxtp_1
X_20532_ _20528_/X _20531_/X _20146_/A _20147_/A VGND VGND VPWR VPWR _20547_/B sky130_fd_sc_hd__o211a_1
X_32518_ _35974_/CLK _32518_/D VGND VGND VPWR VPWR _32518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33498_ _33753_/CLK _33498_/D VGND VGND VPWR VPWR _33498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20463_ _33938_/Q _33874_/Q _33810_/Q _36114_/Q _18362_/X _18364_/X VGND VGND VPWR
+ VPWR _20463_/X sky130_fd_sc_hd__mux4_1
X_23251_ _23251_/A VGND VGND VPWR VPWR _32156_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35237_ _35365_/CLK _35237_/D VGND VGND VPWR VPWR _35237_/Q sky130_fd_sc_hd__dfxtp_1
X_32449_ _36075_/CLK _32449_/D VGND VGND VPWR VPWR _32449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22202_ _22020_/X _22200_/X _22201_/X _22024_/X VGND VGND VPWR VPWR _22202_/X sky130_fd_sc_hd__a22o_1
XFILLER_134_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20394_ _34959_/Q _34895_/Q _34831_/Q _34767_/Q _20166_/X _20167_/X VGND VGND VPWR
+ VPWR _20394_/X sky130_fd_sc_hd__mux4_1
XFILLER_165_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23182_ _23021_/X _32129_/Q _23194_/S VGND VGND VPWR VPWR _23183_/A sky130_fd_sc_hd__mux2_1
X_35168_ _35168_/CLK _35168_/D VGND VGND VPWR VPWR _35168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34119_ _34185_/CLK _34119_/D VGND VGND VPWR VPWR _34119_/Q sky130_fd_sc_hd__dfxtp_1
X_22133_ _32895_/Q _32831_/Q _32767_/Q _32703_/Q _21946_/X _21947_/X VGND VGND VPWR
+ VPWR _22133_/X sky130_fd_sc_hd__mux4_1
X_27990_ _27990_/A VGND VGND VPWR VPWR _34332_/D sky130_fd_sc_hd__clkbuf_1
X_35099_ _35800_/CLK _35099_/D VGND VGND VPWR VPWR _35099_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput240 _32408_/Q VGND VGND VPWR VPWR D3[2] sky130_fd_sc_hd__buf_2
XTAP_6606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput251 _32409_/Q VGND VGND VPWR VPWR D3[3] sky130_fd_sc_hd__buf_2
XTAP_6617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput262 _32410_/Q VGND VGND VPWR VPWR D3[4] sky130_fd_sc_hd__buf_2
XTAP_6628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26941_ _27031_/S VGND VGND VPWR VPWR _26960_/S sky130_fd_sc_hd__buf_4
XFILLER_58_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput273 _32411_/Q VGND VGND VPWR VPWR D3[5] sky130_fd_sc_hd__buf_2
XFILLER_47_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22064_ _35453_/Q _35389_/Q _35325_/Q _35261_/Q _21854_/X _21855_/X VGND VGND VPWR
+ VPWR _22064_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21015_ _21011_/X _21014_/X _20704_/X VGND VGND VPWR VPWR _21016_/D sky130_fd_sc_hd__o21ba_1
XTAP_5927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26872_ _33865_/Q _23460_/X _26888_/S VGND VGND VPWR VPWR _26873_/A sky130_fd_sc_hd__mux2_1
XTAP_5938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29660_ _35093_/Q _29524_/X _29660_/S VGND VGND VPWR VPWR _29661_/A sky130_fd_sc_hd__mux2_1
XTAP_5949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28611_ _27782_/X _34627_/Q _28619_/S VGND VGND VPWR VPWR _28612_/A sky130_fd_sc_hd__mux2_1
X_25823_ _25823_/A VGND VGND VPWR VPWR _33370_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29591_ _29660_/S VGND VGND VPWR VPWR _29610_/S sky130_fd_sc_hd__buf_6
XFILLER_28_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25754_ _24911_/X _33338_/Q _25760_/S VGND VGND VPWR VPWR _25755_/A sky130_fd_sc_hd__mux2_1
X_28542_ _27680_/X _34594_/Q _28556_/S VGND VGND VPWR VPWR _28543_/A sky130_fd_sc_hd__mux2_1
X_22966_ _22965_/X _32047_/Q _22978_/S VGND VGND VPWR VPWR _22967_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24705_ _22949_/X _32874_/Q _24723_/S VGND VGND VPWR VPWR _24706_/A sky130_fd_sc_hd__mux2_1
XFILLER_244_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28473_ _28473_/A VGND VGND VPWR VPWR _34561_/D sky130_fd_sc_hd__clkbuf_1
X_21917_ _22399_/A VGND VGND VPWR VPWR _21917_/X sky130_fd_sc_hd__buf_6
X_25685_ _24809_/X _33305_/Q _25697_/S VGND VGND VPWR VPWR _25686_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22897_ input34/X VGND VGND VPWR VPWR _22897_/X sky130_fd_sc_hd__buf_2
XFILLER_216_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27424_ _27424_/A VGND VGND VPWR VPWR _34095_/D sky130_fd_sc_hd__clkbuf_1
X_24636_ _24636_/A VGND VGND VPWR VPWR _32841_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21848_ _32887_/Q _32823_/Q _32759_/Q _32695_/Q _21593_/X _21594_/X VGND VGND VPWR
+ VPWR _21848_/X sky130_fd_sc_hd__mux4_1
X_27355_ _34063_/Q _27211_/X _27359_/S VGND VGND VPWR VPWR _27356_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24567_ _22946_/X _32809_/Q _24567_/S VGND VGND VPWR VPWR _24568_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21779_ _32117_/Q _32309_/Q _32373_/Q _35893_/Q _21527_/X _21668_/X VGND VGND VPWR
+ VPWR _21779_/X sky130_fd_sc_hd__mux4_1
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26306_ _26306_/A VGND VGND VPWR VPWR _33599_/D sky130_fd_sc_hd__clkbuf_1
X_23518_ _32254_/Q _23420_/X _23536_/S VGND VGND VPWR VPWR _23519_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27286_ _34030_/Q _27109_/X _27296_/S VGND VGND VPWR VPWR _27287_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24498_ _23042_/X _32776_/Q _24516_/S VGND VGND VPWR VPWR _24499_/A sky130_fd_sc_hd__mux2_1
X_29025_ _34822_/Q _27183_/X _29027_/S VGND VGND VPWR VPWR _29026_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26237_ _24827_/X _33567_/Q _26237_/S VGND VGND VPWR VPWR _26238_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23449_ _23449_/A VGND VGND VPWR VPWR _32228_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26168_ _24923_/X _33534_/Q _26186_/S VGND VGND VPWR VPWR _26169_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25119_ _25119_/A VGND VGND VPWR VPWR _33039_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26099_ _26099_/A VGND VGND VPWR VPWR _33501_/D sky130_fd_sc_hd__clkbuf_1
X_18990_ _34663_/Q _34599_/Q _34535_/Q _34471_/Q _18886_/X _18887_/X VGND VGND VPWR
+ VPWR _18990_/X sky130_fd_sc_hd__mux4_1
XFILLER_215_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29927_ _29927_/A VGND VGND VPWR VPWR _35219_/D sky130_fd_sc_hd__clkbuf_1
X_17941_ _17941_/A _17941_/B _17941_/C _17941_/D VGND VGND VPWR VPWR _17942_/A sky130_fd_sc_hd__or4_2
XFILLER_112_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_922 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17872_ _17863_/X _17870_/X _17871_/X VGND VGND VPWR VPWR _17873_/D sky130_fd_sc_hd__o21ba_1
XFILLER_117_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29858_ _29858_/A VGND VGND VPWR VPWR _35186_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19611_ _33145_/Q _36025_/Q _33017_/Q _32953_/Q _19362_/X _19363_/X VGND VGND VPWR
+ VPWR _19611_/X sky130_fd_sc_hd__mux4_1
X_28809_ _28809_/A VGND VGND VPWR VPWR _34719_/D sky130_fd_sc_hd__clkbuf_1
X_16823_ _32619_/Q _32555_/Q _32491_/Q _35947_/Q _16570_/X _16707_/X VGND VGND VPWR
+ VPWR _16823_/X sky130_fd_sc_hd__mux4_1
X_29789_ _35154_/Q _29515_/X _29795_/S VGND VGND VPWR VPWR _29790_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31820_ _31820_/A VGND VGND VPWR VPWR _36116_/D sky130_fd_sc_hd__clkbuf_1
X_19542_ _19506_/X _19540_/X _19541_/X _19509_/X VGND VGND VPWR VPWR _19542_/X sky130_fd_sc_hd__a22o_1
XFILLER_65_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16754_ _16750_/X _16753_/X _16434_/X _16435_/X VGND VGND VPWR VPWR _16769_/B sky130_fd_sc_hd__o211a_1
XFILLER_98_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19473_ _33909_/Q _33845_/Q _33781_/Q _36085_/Q _19324_/X _19325_/X VGND VGND VPWR
+ VPWR _19473_/X sky130_fd_sc_hd__mux4_1
X_31751_ _31751_/A VGND VGND VPWR VPWR _36083_/D sky130_fd_sc_hd__clkbuf_1
X_16685_ _16645_/X _16683_/X _16684_/X _16648_/X VGND VGND VPWR VPWR _16685_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18424_ _35671_/Q _32177_/Q _35543_/Q _35479_/Q _18349_/X _18350_/X VGND VGND VPWR
+ VPWR _18424_/X sky130_fd_sc_hd__mux4_1
X_30702_ _30702_/A VGND VGND VPWR VPWR _35586_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34470_ _36135_/CLK _34470_/D VGND VGND VPWR VPWR _34470_/Q sky130_fd_sc_hd__dfxtp_1
X_31682_ _27831_/X _36051_/Q _31686_/S VGND VGND VPWR VPWR _31683_/A sky130_fd_sc_hd__mux2_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33421_ _34186_/CLK _33421_/D VGND VGND VPWR VPWR _33421_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18355_ _20299_/A VGND VGND VPWR VPWR _18355_/X sky130_fd_sc_hd__buf_4
X_30633_ _30633_/A VGND VGND VPWR VPWR _35553_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17306_ _33401_/Q _33337_/Q _33273_/Q _33209_/Q _17127_/X _17128_/X VGND VGND VPWR
+ VPWR _17306_/X sky130_fd_sc_hd__mux4_1
X_36140_ _36140_/CLK _36140_/D VGND VGND VPWR VPWR _36140_/Q sky130_fd_sc_hd__dfxtp_1
X_33352_ _33420_/CLK _33352_/D VGND VGND VPWR VPWR _33352_/Q sky130_fd_sc_hd__dfxtp_1
X_30564_ _35521_/Q _29463_/X _30576_/S VGND VGND VPWR VPWR _30565_/A sky130_fd_sc_hd__mux2_1
X_18286_ _18363_/A VGND VGND VPWR VPWR _20207_/A sky130_fd_sc_hd__buf_12
XFILLER_30_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32303_ _35952_/CLK _32303_/D VGND VGND VPWR VPWR _32303_/Q sky130_fd_sc_hd__dfxtp_1
X_17237_ _33655_/Q _33591_/Q _33527_/Q _33463_/Q _17200_/X _17201_/X VGND VGND VPWR
+ VPWR _17237_/X sky130_fd_sc_hd__mux4_1
X_36071_ _36072_/CLK _36071_/D VGND VGND VPWR VPWR _36071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33283_ _36097_/CLK _33283_/D VGND VGND VPWR VPWR _33283_/Q sky130_fd_sc_hd__dfxtp_1
X_30495_ _35488_/Q _29360_/X _30513_/S VGND VGND VPWR VPWR _30496_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35022_ _35664_/CLK _35022_/D VGND VGND VPWR VPWR _35022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32234_ _35723_/CLK _32234_/D VGND VGND VPWR VPWR _32234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17168_ _17168_/A VGND VGND VPWR VPWR _31988_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16119_ _16018_/X _16117_/X _16118_/X _16027_/X VGND VGND VPWR VPWR _16119_/X sky130_fd_sc_hd__a22o_1
X_32165_ _35168_/CLK _32165_/D VGND VGND VPWR VPWR _32165_/Q sky130_fd_sc_hd__dfxtp_1
X_17099_ _16853_/X _17097_/X _17098_/X _16856_/X VGND VGND VPWR VPWR _17099_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_805 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31116_ _35783_/Q input44/X _31116_/S VGND VGND VPWR VPWR _31117_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32096_ _32356_/CLK _32096_/D VGND VGND VPWR VPWR _32096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35924_ _35989_/CLK _35924_/D VGND VGND VPWR VPWR _35924_/Q sky130_fd_sc_hd__dfxtp_1
X_31047_ _35750_/Q input8/X _31053_/S VGND VGND VPWR VPWR _31048_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19809_ _20162_/A VGND VGND VPWR VPWR _19809_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_936 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35855_ _35855_/CLK _35855_/D VGND VGND VPWR VPWR _35855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22820_ _34196_/Q _34132_/Q _34068_/Q _34004_/Q _20649_/X _20650_/X VGND VGND VPWR
+ VPWR _22820_/X sky130_fd_sc_hd__mux4_1
X_34806_ _36151_/CLK _34806_/D VGND VGND VPWR VPWR _34806_/Q sky130_fd_sc_hd__dfxtp_1
X_35786_ _35849_/CLK _35786_/D VGND VGND VPWR VPWR _35786_/Q sky130_fd_sc_hd__dfxtp_1
X_32998_ _36005_/CLK _32998_/D VGND VGND VPWR VPWR _32998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_811 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22751_ _35217_/Q _35153_/Q _35089_/Q _32273_/Q _20692_/X _20694_/X VGND VGND VPWR
+ VPWR _22751_/X sky130_fd_sc_hd__mux4_1
X_34737_ _35439_/CLK _34737_/D VGND VGND VPWR VPWR _34737_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31949_ _31949_/A VGND VGND VPWR VPWR _36177_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21702_ _33139_/Q _36019_/Q _33011_/Q _32947_/Q _21662_/X _21663_/X VGND VGND VPWR
+ VPWR _21702_/X sky130_fd_sc_hd__mux4_1
X_25470_ _25470_/A VGND VGND VPWR VPWR _33203_/D sky130_fd_sc_hd__clkbuf_1
X_22682_ _22678_/X _22681_/X _22446_/X _22447_/X VGND VGND VPWR VPWR _22697_/B sky130_fd_sc_hd__o211a_2
X_34668_ _34924_/CLK _34668_/D VGND VGND VPWR VPWR _34668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24421_ _24421_/A VGND VGND VPWR VPWR _32739_/D sky130_fd_sc_hd__clkbuf_1
X_33619_ _34897_/CLK _33619_/D VGND VGND VPWR VPWR _33619_/Q sky130_fd_sc_hd__dfxtp_1
X_21633_ _32881_/Q _32817_/Q _32753_/Q _32689_/Q _21593_/X _21594_/X VGND VGND VPWR
+ VPWR _21633_/X sky130_fd_sc_hd__mux4_1
XFILLER_240_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_551 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34599_ _35365_/CLK _34599_/D VGND VGND VPWR VPWR _34599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27140_ input28/X VGND VGND VPWR VPWR _27140_/X sky130_fd_sc_hd__buf_2
X_24352_ _23027_/X _32707_/Q _24360_/S VGND VGND VPWR VPWR _24353_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21564_ _22399_/A VGND VGND VPWR VPWR _21564_/X sky130_fd_sc_hd__buf_4
XFILLER_21_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23303_ _32173_/Q _23302_/X _23424_/S VGND VGND VPWR VPWR _23304_/A sky130_fd_sc_hd__mux2_1
X_20515_ _18360_/X _20513_/X _20514_/X _18372_/X VGND VGND VPWR VPWR _20515_/X sky130_fd_sc_hd__a22o_1
XFILLER_14_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27071_ _27071_/A VGND VGND VPWR VPWR _33953_/D sky130_fd_sc_hd__clkbuf_1
X_24283_ _22925_/X _32674_/Q _24297_/S VGND VGND VPWR VPWR _24284_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21495_ _32877_/Q _32813_/Q _32749_/Q _32685_/Q _21240_/X _21241_/X VGND VGND VPWR
+ VPWR _21495_/X sky130_fd_sc_hd__mux4_1
XFILLER_219_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26022_ _24908_/X _33465_/Q _26030_/S VGND VGND VPWR VPWR _26023_/A sky130_fd_sc_hd__mux2_1
X_23234_ input12/X VGND VGND VPWR VPWR _23234_/X sky130_fd_sc_hd__buf_4
XFILLER_119_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20446_ _35473_/Q _35409_/Q _35345_/Q _35281_/Q _20260_/X _20261_/X VGND VGND VPWR
+ VPWR _20446_/X sky130_fd_sc_hd__mux4_1
XFILLER_88_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_1323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23165_ _22996_/X _32121_/Q _23173_/S VGND VGND VPWR VPWR _23166_/A sky130_fd_sc_hd__mux2_1
XTAP_7126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20377_ _33167_/Q _36047_/Q _33039_/Q _32975_/Q _20068_/X _20069_/X VGND VGND VPWR
+ VPWR _20377_/X sky130_fd_sc_hd__mux4_1
XFILLER_49_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22116_ _22469_/A VGND VGND VPWR VPWR _22116_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_192_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27973_ _27837_/X _34325_/Q _27973_/S VGND VGND VPWR VPWR _27974_/A sky130_fd_sc_hd__mux2_1
XTAP_6425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23096_ _22894_/X _32088_/Q _23110_/S VGND VGND VPWR VPWR _23097_/A sky130_fd_sc_hd__mux2_1
XTAP_6436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29712_ _35117_/Q _29401_/X _29724_/S VGND VGND VPWR VPWR _29713_/A sky130_fd_sc_hd__mux2_1
XTAP_5724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26924_ _26924_/A VGND VGND VPWR VPWR _33889_/D sky130_fd_sc_hd__clkbuf_1
X_22047_ _22561_/A VGND VGND VPWR VPWR _22047_/X sky130_fd_sc_hd__buf_8
XFILLER_248_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_774 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29643_ _29643_/A VGND VGND VPWR VPWR _35084_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26855_ _33857_/Q _23432_/X _26867_/S VGND VGND VPWR VPWR _26856_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25806_ _24988_/X _33363_/Q _25810_/S VGND VGND VPWR VPWR _25807_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26786_ _33824_/Q _23261_/X _26804_/S VGND VGND VPWR VPWR _26787_/A sky130_fd_sc_hd__mux2_1
X_29574_ _29574_/A VGND VGND VPWR VPWR _35051_/D sky130_fd_sc_hd__clkbuf_1
X_23998_ _22912_/X _32542_/Q _24000_/S VGND VGND VPWR VPWR _23999_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28525_ _27655_/X _34586_/Q _28535_/S VGND VGND VPWR VPWR _28526_/A sky130_fd_sc_hd__mux2_1
X_25737_ _24886_/X _33330_/Q _25739_/S VGND VGND VPWR VPWR _25738_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22949_ input13/X VGND VGND VPWR VPWR _22949_/X sky130_fd_sc_hd__buf_2
XFILLER_21_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16470_ _32609_/Q _32545_/Q _32481_/Q _35937_/Q _16217_/X _16354_/X VGND VGND VPWR
+ VPWR _16470_/X sky130_fd_sc_hd__mux4_1
X_25668_ _25668_/A VGND VGND VPWR VPWR _33297_/D sky130_fd_sc_hd__clkbuf_1
X_28456_ _28456_/A VGND VGND VPWR VPWR _34553_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24619_ _24619_/A VGND VGND VPWR VPWR _32833_/D sky130_fd_sc_hd__clkbuf_1
X_27407_ _27407_/A VGND VGND VPWR VPWR _34087_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28387_ _28387_/A VGND VGND VPWR VPWR _34520_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25599_ _25599_/A VGND VGND VPWR VPWR _33264_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27338_ _34055_/Q _27186_/X _27338_/S VGND VGND VPWR VPWR _27339_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18140_ _32913_/Q _32849_/Q _32785_/Q _32721_/Q _15984_/X _15987_/X VGND VGND VPWR
+ VPWR _18140_/X sky130_fd_sc_hd__mux4_1
XFILLER_223_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_746 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18071_ _17905_/X _18069_/X _18070_/X _17910_/X VGND VGND VPWR VPWR _18071_/X sky130_fd_sc_hd__a22o_1
X_27269_ _34022_/Q _27084_/X _27275_/S VGND VGND VPWR VPWR _27270_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17022_ _16846_/X _17020_/X _17021_/X _16851_/X VGND VGND VPWR VPWR _17022_/X sky130_fd_sc_hd__a22o_1
X_29008_ _29056_/S VGND VGND VPWR VPWR _29027_/S sky130_fd_sc_hd__buf_4
XFILLER_184_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30280_ _30280_/A VGND VGND VPWR VPWR _35386_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_940 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18973_ _33895_/Q _33831_/Q _33767_/Q _36071_/Q _18971_/X _18972_/X VGND VGND VPWR
+ VPWR _18973_/X sky130_fd_sc_hd__mux4_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17924_ _17920_/X _17923_/X _17846_/X _17847_/X VGND VGND VPWR VPWR _17941_/B sky130_fd_sc_hd__o211a_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33970_ _34035_/CLK _33970_/D VGND VGND VPWR VPWR _33970_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32921_ _34135_/CLK _32921_/D VGND VGND VPWR VPWR _32921_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_722 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17855_ _33096_/Q _32072_/Q _35848_/Q _35784_/Q _17784_/X _17785_/X VGND VGND VPWR
+ VPWR _17855_/X sky130_fd_sc_hd__mux4_1
XFILLER_61_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35640_ _35704_/CLK _35640_/D VGND VGND VPWR VPWR _35640_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16806_ _34410_/Q _36138_/Q _34282_/Q _34218_/Q _16523_/X _16524_/X VGND VGND VPWR
+ VPWR _16806_/X sky130_fd_sc_hd__mux4_1
XFILLER_187_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32852_ _32869_/CLK _32852_/D VGND VGND VPWR VPWR _32852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17786_ _33094_/Q _32070_/Q _35846_/Q _35782_/Q _17784_/X _17785_/X VGND VGND VPWR
+ VPWR _17786_/X sky130_fd_sc_hd__mux4_1
XFILLER_82_928 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31803_ _36108_/Q input50/X _31813_/S VGND VGND VPWR VPWR _31804_/A sky130_fd_sc_hd__mux2_1
X_19525_ _19521_/X _19524_/X _19451_/X VGND VGND VPWR VPWR _19535_/C sky130_fd_sc_hd__o21ba_1
X_35571_ _35699_/CLK _35571_/D VGND VGND VPWR VPWR _35571_/Q sky130_fd_sc_hd__dfxtp_1
X_16737_ _16737_/A _16737_/B _16737_/C _16737_/D VGND VGND VPWR VPWR _16738_/A sky130_fd_sc_hd__or4_2
X_32783_ _32911_/CLK _32783_/D VGND VGND VPWR VPWR _32783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_1224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34522_ _36229_/CLK _34522_/D VGND VGND VPWR VPWR _34522_/Q sky130_fd_sc_hd__dfxtp_1
X_31734_ _36075_/Q input14/X _31750_/S VGND VGND VPWR VPWR _31735_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19456_ _19456_/A VGND VGND VPWR VPWR _19456_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_223_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16668_ _34151_/Q _34087_/Q _34023_/Q _33959_/Q _16387_/X _16388_/X VGND VGND VPWR
+ VPWR _16668_/X sky130_fd_sc_hd__mux4_2
XFILLER_179_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18407_ _18407_/A VGND VGND VPWR VPWR _32406_/D sky130_fd_sc_hd__buf_4
X_34453_ _36181_/CLK _34453_/D VGND VGND VPWR VPWR _34453_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31665_ _31665_/A VGND VGND VPWR VPWR _36042_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19387_ _34930_/Q _34866_/Q _34802_/Q _34738_/Q _19107_/X _19108_/X VGND VGND VPWR
+ VPWR _19387_/X sky130_fd_sc_hd__mux4_1
X_16599_ _16493_/X _16597_/X _16598_/X _16498_/X VGND VGND VPWR VPWR _16599_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33404_ _36093_/CLK _33404_/D VGND VGND VPWR VPWR _33404_/Q sky130_fd_sc_hd__dfxtp_1
X_18338_ _18363_/A VGND VGND VPWR VPWR _20134_/A sky130_fd_sc_hd__buf_12
X_30616_ _30616_/A VGND VGND VPWR VPWR _35545_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34384_ _35664_/CLK _34384_/D VGND VGND VPWR VPWR _34384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31596_ _31686_/S VGND VGND VPWR VPWR _31615_/S sky130_fd_sc_hd__buf_4
XFILLER_30_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36123_ _36127_/CLK _36123_/D VGND VGND VPWR VPWR _36123_/Q sky130_fd_sc_hd__dfxtp_1
X_33335_ _36087_/CLK _33335_/D VGND VGND VPWR VPWR _33335_/Q sky130_fd_sc_hd__dfxtp_1
X_18269_ _18265_/X _18268_/X _17857_/A VGND VGND VPWR VPWR _18277_/C sky130_fd_sc_hd__o21ba_1
XFILLER_136_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30547_ _35513_/Q _29438_/X _30555_/S VGND VGND VPWR VPWR _30548_/A sky130_fd_sc_hd__mux2_1
X_20300_ _34700_/Q _34636_/Q _34572_/Q _34508_/Q _20298_/X _20299_/X VGND VGND VPWR
+ VPWR _20300_/X sky130_fd_sc_hd__mux4_1
XFILLER_163_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36054_ _36054_/CLK _36054_/D VGND VGND VPWR VPWR _36054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21280_ _32871_/Q _32807_/Q _32743_/Q _32679_/Q _21240_/X _21241_/X VGND VGND VPWR
+ VPWR _21280_/X sky130_fd_sc_hd__mux4_1
X_33266_ _33393_/CLK _33266_/D VGND VGND VPWR VPWR _33266_/Q sky130_fd_sc_hd__dfxtp_1
X_30478_ _35480_/Q _29336_/X _30492_/S VGND VGND VPWR VPWR _30479_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35005_ _35645_/CLK _35005_/D VGND VGND VPWR VPWR _35005_/Q sky130_fd_sc_hd__dfxtp_1
X_20231_ _20227_/X _20230_/X _20157_/X VGND VGND VPWR VPWR _20241_/C sky130_fd_sc_hd__o21ba_1
X_32217_ _35453_/CLK _32217_/D VGND VGND VPWR VPWR _32217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33197_ _36077_/CLK _33197_/D VGND VGND VPWR VPWR _33197_/Q sky130_fd_sc_hd__dfxtp_1
X_20162_ _20162_/A VGND VGND VPWR VPWR _20162_/X sky130_fd_sc_hd__clkbuf_4
X_32148_ _35922_/CLK _32148_/D VGND VGND VPWR VPWR _32148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20093_ _34950_/Q _34886_/Q _34822_/Q _34758_/Q _19813_/X _19814_/X VGND VGND VPWR
+ VPWR _20093_/X sky130_fd_sc_hd__mux4_1
X_24970_ input51/X VGND VGND VPWR VPWR _24970_/X sky130_fd_sc_hd__buf_6
X_32079_ _35853_/CLK _32079_/D VGND VGND VPWR VPWR _32079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23921_ _22999_/X _32506_/Q _23927_/S VGND VGND VPWR VPWR _23922_/A sky130_fd_sc_hd__mux2_1
XTAP_4319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35907_ _35907_/CLK _35907_/D VGND VGND VPWR VPWR _35907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_245_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26640_ _33755_/Q _23246_/X _26648_/S VGND VGND VPWR VPWR _26641_/A sky130_fd_sc_hd__mux2_1
XTAP_3618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23852_ _22897_/X _32473_/Q _23864_/S VGND VGND VPWR VPWR _23853_/A sky130_fd_sc_hd__mux2_1
X_35838_ _35903_/CLK _35838_/D VGND VGND VPWR VPWR _35838_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22803_ _35731_/Q _32243_/Q _35603_/Q _35539_/Q _20593_/X _20595_/X VGND VGND VPWR
+ VPWR _22803_/X sky130_fd_sc_hd__mux4_1
XFILLER_44_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26571_ _26571_/A VGND VGND VPWR VPWR _33724_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35769_ _35769_/CLK _35769_/D VGND VGND VPWR VPWR _35769_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23783_ _23783_/A VGND VGND VPWR VPWR _32377_/D sky130_fd_sc_hd__clkbuf_1
X_20995_ _32607_/Q _32543_/Q _32479_/Q _35935_/Q _20817_/X _20954_/X VGND VGND VPWR
+ VPWR _20995_/X sky130_fd_sc_hd__mux4_1
XFILLER_37_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25522_ _24967_/X _33228_/Q _25532_/S VGND VGND VPWR VPWR _25523_/A sky130_fd_sc_hd__mux2_1
XFILLER_198_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28310_ _27735_/X _34484_/Q _28328_/S VGND VGND VPWR VPWR _28311_/A sky130_fd_sc_hd__mux2_1
X_22734_ _22512_/X _22732_/X _22733_/X _22515_/X VGND VGND VPWR VPWR _22734_/X sky130_fd_sc_hd__a22o_1
X_29290_ _29290_/A VGND VGND VPWR VPWR _34947_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28241_ _27834_/X _34452_/Q _28243_/S VGND VGND VPWR VPWR _28242_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25453_ _24865_/X _33195_/Q _25469_/S VGND VGND VPWR VPWR _25454_/A sky130_fd_sc_hd__mux2_1
X_22665_ _22464_/X _22663_/X _22664_/X _22469_/X VGND VGND VPWR VPWR _22665_/X sky130_fd_sc_hd__a22o_1
XFILLER_111_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1079 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24404_ _24404_/A VGND VGND VPWR VPWR _32731_/D sky130_fd_sc_hd__clkbuf_1
X_21616_ _21405_/X _21614_/X _21615_/X _21410_/X VGND VGND VPWR VPWR _21616_/X sky130_fd_sc_hd__a22o_1
X_28172_ _27732_/X _34419_/Q _28172_/S VGND VGND VPWR VPWR _28173_/A sky130_fd_sc_hd__mux2_1
X_25384_ _25384_/A VGND VGND VPWR VPWR _33163_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22596_ _22309_/X _22594_/X _22595_/X _22312_/X VGND VGND VPWR VPWR _22596_/X sky130_fd_sc_hd__a22o_1
XFILLER_205_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27123_ _27123_/A VGND VGND VPWR VPWR _33970_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24335_ _23002_/X _32699_/Q _24339_/S VGND VGND VPWR VPWR _24336_/A sky130_fd_sc_hd__mux2_1
X_21547_ _21543_/X _21546_/X _21412_/X VGND VGND VPWR VPWR _21548_/D sky130_fd_sc_hd__o21ba_1
XFILLER_193_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27054_ _33948_/Q _27053_/X _27063_/S VGND VGND VPWR VPWR _27055_/A sky130_fd_sc_hd__mux2_1
X_24266_ _22900_/X _32666_/Q _24276_/S VGND VGND VPWR VPWR _24267_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21478_ _34412_/Q _36140_/Q _34284_/Q _34220_/Q _21476_/X _21477_/X VGND VGND VPWR
+ VPWR _21478_/X sky130_fd_sc_hd__mux4_1
XFILLER_153_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26005_ _24883_/X _33457_/Q _26009_/S VGND VGND VPWR VPWR _26006_/A sky130_fd_sc_hd__mux2_1
X_23217_ _23073_/X _32146_/Q _23223_/S VGND VGND VPWR VPWR _23218_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20429_ _33681_/Q _33617_/Q _33553_/Q _33489_/Q _20206_/X _20207_/X VGND VGND VPWR
+ VPWR _20429_/X sky130_fd_sc_hd__mux4_1
XFILLER_181_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24197_ _32635_/Q _23411_/X _24201_/S VGND VGND VPWR VPWR _24198_/A sky130_fd_sc_hd__mux2_1
XTAP_6200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23148_ _22971_/X _32113_/Q _23152_/S VGND VGND VPWR VPWR _23149_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27956_ _27956_/A VGND VGND VPWR VPWR _34316_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23079_ input59/X VGND VGND VPWR VPWR _23079_/X sky130_fd_sc_hd__buf_2
XFILLER_0_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26907_ _26907_/A VGND VGND VPWR VPWR _33881_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27887_ _27887_/A VGND VGND VPWR VPWR _34283_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29626_ _29626_/A VGND VGND VPWR VPWR _35076_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17640_ _17351_/X _17638_/X _17639_/X _17354_/X VGND VGND VPWR VPWR _17640_/X sky130_fd_sc_hd__a22o_1
XTAP_5598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26838_ _33849_/Q _23405_/X _26846_/S VGND VGND VPWR VPWR _26839_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17571_ _17567_/X _17570_/X _17493_/X _17494_/X VGND VGND VPWR VPWR _17588_/B sky130_fd_sc_hd__o211a_1
X_29557_ _29557_/A VGND VGND VPWR VPWR _35043_/D sky130_fd_sc_hd__clkbuf_1
X_26769_ _33816_/Q _23237_/X _26783_/S VGND VGND VPWR VPWR _26770_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_1192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19310_ _20016_/A VGND VGND VPWR VPWR _19310_/X sky130_fd_sc_hd__buf_4
XFILLER_232_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28508_ _28508_/A VGND VGND VPWR VPWR _34578_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16522_ _16447_/X _16520_/X _16521_/X _16450_/X VGND VGND VPWR VPWR _16522_/X sky130_fd_sc_hd__a22o_1
XFILLER_147_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29488_ input47/X VGND VGND VPWR VPWR _29488_/X sky130_fd_sc_hd__buf_2
XFILLER_45_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_808 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19241_ _34670_/Q _34606_/Q _34542_/Q _34478_/Q _19239_/X _19240_/X VGND VGND VPWR
+ VPWR _19241_/X sky130_fd_sc_hd__mux4_1
X_16453_ _34400_/Q _36128_/Q _34272_/Q _34208_/Q _16170_/X _16171_/X VGND VGND VPWR
+ VPWR _16453_/X sky130_fd_sc_hd__mux4_2
X_28439_ _28439_/A VGND VGND VPWR VPWR _34545_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16384_ _16384_/A _16384_/B _16384_/C _16384_/D VGND VGND VPWR VPWR _16385_/A sky130_fd_sc_hd__or4_4
X_19172_ _19168_/X _19171_/X _19098_/X VGND VGND VPWR VPWR _19182_/C sky130_fd_sc_hd__o21ba_1
X_31450_ _31450_/A VGND VGND VPWR VPWR _35940_/D sky130_fd_sc_hd__clkbuf_1
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18123_ _34448_/Q _36176_/Q _34320_/Q _34256_/Q _17935_/X _17936_/X VGND VGND VPWR
+ VPWR _18123_/X sky130_fd_sc_hd__mux4_1
X_30401_ _30470_/S VGND VGND VPWR VPWR _30420_/S sky130_fd_sc_hd__buf_6
XFILLER_200_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31381_ _27785_/X _35908_/Q _31387_/S VGND VGND VPWR VPWR _31382_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33120_ _36003_/CLK _33120_/D VGND VGND VPWR VPWR _33120_/Q sky130_fd_sc_hd__dfxtp_1
X_18054_ _35662_/Q _35022_/Q _34382_/Q _33742_/Q _17850_/X _17851_/X VGND VGND VPWR
+ VPWR _18054_/X sky130_fd_sc_hd__mux4_1
X_30332_ _30332_/A VGND VGND VPWR VPWR _35411_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17005_ _33072_/Q _32048_/Q _35824_/Q _35760_/Q _16725_/X _16726_/X VGND VGND VPWR
+ VPWR _17005_/X sky130_fd_sc_hd__mux4_1
X_33051_ _34007_/CLK _33051_/D VGND VGND VPWR VPWR _33051_/Q sky130_fd_sc_hd__dfxtp_1
X_30263_ _30263_/A VGND VGND VPWR VPWR _35378_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32002_ _36197_/CLK _32002_/D VGND VGND VPWR VPWR _32002_/Q sky130_fd_sc_hd__dfxtp_1
X_30194_ _35346_/Q _29515_/X _30200_/S VGND VGND VPWR VPWR _30195_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18956_ _34662_/Q _34598_/Q _34534_/Q _34470_/Q _18886_/X _18887_/X VGND VGND VPWR
+ VPWR _18956_/X sky130_fd_sc_hd__mux4_1
X_17907_ _17907_/A VGND VGND VPWR VPWR _17907_/X sky130_fd_sc_hd__buf_4
XFILLER_66_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33953_ _34594_/CLK _33953_/D VGND VGND VPWR VPWR _33953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18887_ _20299_/A VGND VGND VPWR VPWR _18887_/X sky130_fd_sc_hd__buf_4
X_32904_ _32904_/CLK _32904_/D VGND VGND VPWR VPWR _32904_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17838_ _17838_/A VGND VGND VPWR VPWR _17838_/X sky130_fd_sc_hd__buf_2
XFILLER_187_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33884_ _36058_/CLK _33884_/D VGND VGND VPWR VPWR _33884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35623_ _35624_/CLK _35623_/D VGND VGND VPWR VPWR _35623_/Q sky130_fd_sc_hd__dfxtp_1
X_32835_ _35907_/CLK _32835_/D VGND VGND VPWR VPWR _32835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17769_ _17774_/A VGND VGND VPWR VPWR _17769_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_242_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19508_ _33910_/Q _33846_/Q _33782_/Q _36086_/Q _19324_/X _19325_/X VGND VGND VPWR
+ VPWR _19508_/X sky130_fd_sc_hd__mux4_1
X_35554_ _35554_/CLK _35554_/D VGND VGND VPWR VPWR _35554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20780_ _20740_/X _20778_/X _20779_/X _20745_/X VGND VGND VPWR VPWR _20780_/X sky130_fd_sc_hd__a22o_1
X_32766_ _32891_/CLK _32766_/D VGND VGND VPWR VPWR _32766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34505_ _34633_/CLK _34505_/D VGND VGND VPWR VPWR _34505_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31717_ _36067_/Q input5/X _31729_/S VGND VGND VPWR VPWR _31718_/A sky130_fd_sc_hd__mux2_1
X_19439_ _19367_/X _19437_/X _19438_/X _19371_/X VGND VGND VPWR VPWR _19439_/X sky130_fd_sc_hd__a22o_1
X_35485_ _35613_/CLK _35485_/D VGND VGND VPWR VPWR _35485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_1339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32697_ _32887_/CLK _32697_/D VGND VGND VPWR VPWR _32697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34436_ _36164_/CLK _34436_/D VGND VGND VPWR VPWR _34436_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22450_ _22450_/A VGND VGND VPWR VPWR _22450_/X sky130_fd_sc_hd__buf_4
X_31648_ _31648_/A VGND VGND VPWR VPWR _36034_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21401_ _34666_/Q _34602_/Q _34538_/Q _34474_/Q _21186_/X _21187_/X VGND VGND VPWR
+ VPWR _21401_/X sky130_fd_sc_hd__mux4_1
X_22381_ _35654_/Q _35014_/Q _34374_/Q _33734_/Q _22097_/X _22098_/X VGND VGND VPWR
+ VPWR _22381_/X sky130_fd_sc_hd__mux4_1
X_34367_ _35777_/CLK _34367_/D VGND VGND VPWR VPWR _34367_/Q sky130_fd_sc_hd__dfxtp_1
X_31579_ _31579_/A VGND VGND VPWR VPWR _36001_/D sky130_fd_sc_hd__clkbuf_1
X_36106_ _36106_/CLK _36106_/D VGND VGND VPWR VPWR _36106_/Q sky130_fd_sc_hd__dfxtp_1
X_24120_ _32598_/Q _23225_/X _24138_/S VGND VGND VPWR VPWR _24121_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33318_ _35620_/CLK _33318_/D VGND VGND VPWR VPWR _33318_/Q sky130_fd_sc_hd__dfxtp_1
X_21332_ _21047_/X _21330_/X _21331_/X _21050_/X VGND VGND VPWR VPWR _21332_/X sky130_fd_sc_hd__a22o_1
XFILLER_15_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34298_ _36153_/CLK _34298_/D VGND VGND VPWR VPWR _34298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36037_ _36037_/CLK _36037_/D VGND VGND VPWR VPWR _36037_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24051_ _22990_/X _32567_/Q _24063_/S VGND VGND VPWR VPWR _24052_/A sky130_fd_sc_hd__mux2_1
X_33249_ _36065_/CLK _33249_/D VGND VGND VPWR VPWR _33249_/Q sky130_fd_sc_hd__dfxtp_1
X_21263_ _21052_/X _21261_/X _21262_/X _21057_/X VGND VGND VPWR VPWR _21263_/X sky130_fd_sc_hd__a22o_1
XFILLER_190_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_1462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23002_ input31/X VGND VGND VPWR VPWR _23002_/X sky130_fd_sc_hd__buf_2
X_20214_ _33930_/Q _33866_/Q _33802_/Q _36106_/Q _20030_/X _20031_/X VGND VGND VPWR
+ VPWR _20214_/X sky130_fd_sc_hd__mux4_1
XFILLER_150_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21194_ _21190_/X _21193_/X _21059_/X VGND VGND VPWR VPWR _21195_/D sky130_fd_sc_hd__o21ba_1
X_27810_ input50/X VGND VGND VPWR VPWR _27810_/X sky130_fd_sc_hd__clkbuf_4
X_20145_ _20073_/X _20143_/X _20144_/X _20077_/X VGND VGND VPWR VPWR _20145_/X sky130_fd_sc_hd__a22o_1
X_28790_ _34710_/Q _27033_/X _28808_/S VGND VGND VPWR VPWR _28791_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24953_ _24953_/A VGND VGND VPWR VPWR _32967_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27741_ _27741_/A VGND VGND VPWR VPWR _34229_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20076_ _32902_/Q _32838_/Q _32774_/Q _32710_/Q _19999_/X _20000_/X VGND VGND VPWR
+ VPWR _20076_/X sky130_fd_sc_hd__mux4_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23904_ _22974_/X _32498_/Q _23906_/S VGND VGND VPWR VPWR _23905_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27672_ _27672_/A VGND VGND VPWR VPWR _34207_/D sky130_fd_sc_hd__clkbuf_1
X_24884_ _24883_/X _32945_/Q _24890_/S VGND VGND VPWR VPWR _24885_/A sky130_fd_sc_hd__mux2_1
XTAP_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29411_ _34992_/Q _29410_/X _29420_/S VGND VGND VPWR VPWR _29412_/A sky130_fd_sc_hd__mux2_1
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26623_ _26623_/A VGND VGND VPWR VPWR _33749_/D sky130_fd_sc_hd__clkbuf_1
X_23835_ _23835_/A VGND VGND VPWR VPWR _32402_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29342_ input45/X VGND VGND VPWR VPWR _29342_/X sky130_fd_sc_hd__buf_2
X_26554_ _24892_/X _33716_/Q _26572_/S VGND VGND VPWR VPWR _26555_/A sky130_fd_sc_hd__mux2_1
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23766_ _23766_/A VGND VGND VPWR VPWR _32369_/D sky130_fd_sc_hd__clkbuf_1
X_20978_ _35166_/Q _35102_/Q _35038_/Q _32158_/Q _20904_/X _20905_/X VGND VGND VPWR
+ VPWR _20978_/X sky130_fd_sc_hd__mux4_1
XFILLER_198_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25505_ _24942_/X _33220_/Q _25511_/S VGND VGND VPWR VPWR _25506_/A sky130_fd_sc_hd__mux2_1
X_22717_ _33104_/Q _32080_/Q _35856_/Q _35792_/Q _20679_/X _20680_/X VGND VGND VPWR
+ VPWR _22717_/X sky130_fd_sc_hd__mux4_1
XFILLER_242_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26485_ _26485_/A VGND VGND VPWR VPWR _33684_/D sky130_fd_sc_hd__clkbuf_1
X_29273_ _29273_/A VGND VGND VPWR VPWR _34939_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23697_ _23697_/A VGND VGND VPWR VPWR _32338_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_207_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28224_ _28224_/A VGND VGND VPWR VPWR _34443_/D sky130_fd_sc_hd__clkbuf_1
X_25436_ _24840_/X _33187_/Q _25448_/S VGND VGND VPWR VPWR _25437_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22648_ _22365_/X _22646_/X _22647_/X _22371_/X VGND VGND VPWR VPWR _22648_/X sky130_fd_sc_hd__a22o_1
XFILLER_224_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_194_CLK clkbuf_6_49__f_CLK/X VGND VGND VPWR VPWR _35852_/CLK sky130_fd_sc_hd__clkbuf_16
X_25367_ _25367_/A VGND VGND VPWR VPWR _33155_/D sky130_fd_sc_hd__clkbuf_1
X_28155_ _28155_/A VGND VGND VPWR VPWR _34410_/D sky130_fd_sc_hd__clkbuf_1
X_22579_ _33932_/Q _33868_/Q _33804_/Q _36108_/Q _22330_/X _22331_/X VGND VGND VPWR
+ VPWR _22579_/X sky130_fd_sc_hd__mux4_1
XFILLER_210_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27106_ input16/X VGND VGND VPWR VPWR _27106_/X sky130_fd_sc_hd__buf_2
X_24318_ _22977_/X _32691_/Q _24318_/S VGND VGND VPWR VPWR _24319_/A sky130_fd_sc_hd__mux2_1
X_28086_ _34378_/Q _27196_/X _28100_/S VGND VGND VPWR VPWR _28087_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25298_ _25298_/A VGND VGND VPWR VPWR _33122_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_523 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27037_ _27037_/A VGND VGND VPWR VPWR _33942_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24249_ _32660_/Q _23495_/X _24251_/S VGND VGND VPWR VPWR _24250_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18810_ _32866_/Q _32802_/Q _32738_/Q _32674_/Q _18587_/X _18588_/X VGND VGND VPWR
+ VPWR _18810_/X sky130_fd_sc_hd__mux4_1
XTAP_6030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19790_ _32126_/Q _32318_/Q _32382_/Q _35902_/Q _19580_/X _19721_/X VGND VGND VPWR
+ VPWR _19790_/X sky130_fd_sc_hd__mux4_1
X_28988_ _34804_/Q _27127_/X _29006_/S VGND VGND VPWR VPWR _28989_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput95 _31972_/Q VGND VGND VPWR VPWR D1[14] sky130_fd_sc_hd__buf_2
XFILLER_1_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18741_ _18592_/X _18737_/X _18740_/X _18595_/X VGND VGND VPWR VPWR _18741_/X sky130_fd_sc_hd__a22o_1
XTAP_6085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27939_ _27939_/A VGND VGND VPWR VPWR _34308_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30950_ _35704_/Q input28/X _30960_/S VGND VGND VPWR VPWR _30951_/A sky130_fd_sc_hd__mux2_1
X_18672_ _20235_/A VGND VGND VPWR VPWR _18672_/X sky130_fd_sc_hd__buf_6
XFILLER_97_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17623_ _34178_/Q _34114_/Q _34050_/Q _33986_/Q _17446_/X _17447_/X VGND VGND VPWR
+ VPWR _17623_/X sky130_fd_sc_hd__mux4_1
XFILLER_149_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29609_ _29609_/A VGND VGND VPWR VPWR _35068_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_236_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30881_ _35671_/Q input12/X _30897_/S VGND VGND VPWR VPWR _30882_/A sky130_fd_sc_hd__mux2_1
XTAP_4694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32620_ _36141_/CLK _32620_/D VGND VGND VPWR VPWR _32620_/Q sky130_fd_sc_hd__dfxtp_1
X_17554_ _17907_/A VGND VGND VPWR VPWR _17554_/X sky130_fd_sc_hd__buf_4
XTAP_3993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16505_ _16499_/X _16504_/X _16426_/X VGND VGND VPWR VPWR _16529_/A sky130_fd_sc_hd__o21ba_1
X_32551_ _35941_/CLK _32551_/D VGND VGND VPWR VPWR _32551_/Q sky130_fd_sc_hd__dfxtp_1
X_17485_ _17838_/A VGND VGND VPWR VPWR _17485_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_177_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19224_ _32622_/Q _32558_/Q _32494_/Q _35950_/Q _19223_/X _19007_/X VGND VGND VPWR
+ VPWR _19224_/X sky130_fd_sc_hd__mux4_1
X_31502_ _31502_/A VGND VGND VPWR VPWR _35965_/D sky130_fd_sc_hd__clkbuf_1
X_35270_ _35847_/CLK _35270_/D VGND VGND VPWR VPWR _35270_/Q sky130_fd_sc_hd__dfxtp_1
X_16436_ _16430_/X _16433_/X _16434_/X _16435_/X VGND VGND VPWR VPWR _16461_/B sky130_fd_sc_hd__o211a_2
X_32482_ _35938_/CLK _32482_/D VGND VGND VPWR VPWR _32482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34221_ _36141_/CLK _34221_/D VGND VGND VPWR VPWR _34221_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31433_ _31433_/A VGND VGND VPWR VPWR _35932_/D sky130_fd_sc_hd__clkbuf_1
X_19155_ _33900_/Q _33836_/Q _33772_/Q _36076_/Q _18971_/X _18972_/X VGND VGND VPWR
+ VPWR _19155_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_185_CLK clkbuf_leaf_65_CLK/A VGND VGND VPWR VPWR _36051_/CLK sky130_fd_sc_hd__clkbuf_16
X_16367_ _16360_/X _16366_/X _16044_/X _16046_/X VGND VGND VPWR VPWR _16384_/B sky130_fd_sc_hd__o211a_1
XFILLER_191_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18106_ _32656_/Q _32592_/Q _32528_/Q _35984_/Q _17982_/X _16877_/A VGND VGND VPWR
+ VPWR _18106_/X sky130_fd_sc_hd__mux4_1
X_34152_ _36065_/CLK _34152_/D VGND VGND VPWR VPWR _34152_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16298_ _35420_/Q _35356_/Q _35292_/Q _35228_/Q _16195_/X _16196_/X VGND VGND VPWR
+ VPWR _16298_/X sky130_fd_sc_hd__mux4_1
X_31364_ _27760_/X _35900_/Q _31366_/S VGND VGND VPWR VPWR _31365_/A sky130_fd_sc_hd__mux2_1
X_19086_ _19014_/X _19084_/X _19085_/X _19018_/X VGND VGND VPWR VPWR _19086_/X sky130_fd_sc_hd__a22o_1
X_33103_ _35852_/CLK _33103_/D VGND VGND VPWR VPWR _33103_/Q sky130_fd_sc_hd__dfxtp_1
X_18037_ _18037_/A _18037_/B _18037_/C _18037_/D VGND VGND VPWR VPWR _18038_/A sky130_fd_sc_hd__or4_2
X_30315_ _35403_/Q _29494_/X _30327_/S VGND VGND VPWR VPWR _30316_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34083_ _34151_/CLK _34083_/D VGND VGND VPWR VPWR _34083_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_6_33__f_CLK clkbuf_5_16_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_33__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_31295_ _27658_/X _35867_/Q _31303_/S VGND VGND VPWR VPWR _31296_/A sky130_fd_sc_hd__mux2_1
X_33034_ _36042_/CLK _33034_/D VGND VGND VPWR VPWR _33034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30246_ _35370_/Q _29391_/X _30264_/S VGND VGND VPWR VPWR _30247_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30177_ _30177_/A VGND VGND VPWR VPWR _35337_/D sky130_fd_sc_hd__clkbuf_1
X_19988_ _33668_/Q _33604_/Q _33540_/Q _33476_/Q _19853_/X _19854_/X VGND VGND VPWR
+ VPWR _19988_/X sky130_fd_sc_hd__mux4_1
XFILLER_115_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18939_ _32102_/Q _32294_/Q _32358_/Q _35878_/Q _18874_/X _18662_/X VGND VGND VPWR
+ VPWR _18939_/X sky130_fd_sc_hd__mux4_1
XFILLER_246_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34985_ _35625_/CLK _34985_/D VGND VGND VPWR VPWR _34985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_834 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33936_ _36113_/CLK _33936_/D VGND VGND VPWR VPWR _33936_/Q sky130_fd_sc_hd__dfxtp_1
X_21950_ _21944_/X _21949_/X _21740_/X _21741_/X VGND VGND VPWR VPWR _21971_/B sky130_fd_sc_hd__o211a_1
XFILLER_243_804 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20901_ _20897_/X _20898_/X _20899_/X _20900_/X VGND VGND VPWR VPWR _20901_/X sky130_fd_sc_hd__a22o_1
XFILLER_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33867_ _36106_/CLK _33867_/D VGND VGND VPWR VPWR _33867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21881_ _32120_/Q _32312_/Q _32376_/Q _35896_/Q _21880_/X _21668_/X VGND VGND VPWR
+ VPWR _21881_/X sky130_fd_sc_hd__mux4_1
XFILLER_227_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35606_ _35993_/CLK _35606_/D VGND VGND VPWR VPWR _35606_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23620_ _23620_/A VGND VGND VPWR VPWR _32301_/D sky130_fd_sc_hd__clkbuf_1
X_20832_ _20828_/X _20831_/X _20675_/X VGND VGND VPWR VPWR _20842_/C sky130_fd_sc_hd__o21ba_1
X_32818_ _32818_/CLK _32818_/D VGND VGND VPWR VPWR _32818_/Q sky130_fd_sc_hd__dfxtp_1
X_33798_ _36159_/CLK _33798_/D VGND VGND VPWR VPWR _33798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23551_ _32270_/Q _23475_/X _23557_/S VGND VGND VPWR VPWR _23552_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35537_ _35729_/CLK _35537_/D VGND VGND VPWR VPWR _35537_/Q sky130_fd_sc_hd__dfxtp_1
X_20763_ _35416_/Q _35352_/Q _35288_/Q _35224_/Q _20662_/X _20664_/X VGND VGND VPWR
+ VPWR _20763_/X sky130_fd_sc_hd__mux4_1
XFILLER_51_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32749_ _32877_/CLK _32749_/D VGND VGND VPWR VPWR _32749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22502_ _22498_/X _22501_/X _22471_/X VGND VGND VPWR VPWR _22503_/D sky130_fd_sc_hd__o21ba_1
XFILLER_11_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26270_ _26270_/A VGND VGND VPWR VPWR _33582_/D sky130_fd_sc_hd__clkbuf_1
X_23482_ _32239_/Q _23481_/X _23485_/S VGND VGND VPWR VPWR _23483_/A sky130_fd_sc_hd__mux2_1
X_35468_ _35596_/CLK _35468_/D VGND VGND VPWR VPWR _35468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20694_ _21477_/A VGND VGND VPWR VPWR _20694_/X sky130_fd_sc_hd__buf_4
XFILLER_149_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25221_ _25221_/A VGND VGND VPWR VPWR _33086_/D sky130_fd_sc_hd__clkbuf_1
X_22433_ _22433_/A VGND VGND VPWR VPWR _22433_/X sky130_fd_sc_hd__buf_4
X_34419_ _34611_/CLK _34419_/D VGND VGND VPWR VPWR _34419_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_176_CLK clkbuf_leaf_77_CLK/A VGND VGND VPWR VPWR _35860_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_13_1306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35399_ _35463_/CLK _35399_/D VGND VGND VPWR VPWR _35399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25152_ _33054_/Q _23255_/X _25154_/S VGND VGND VPWR VPWR _25153_/A sky130_fd_sc_hd__mux2_1
X_22364_ _22360_/X _22363_/X _22085_/X VGND VGND VPWR VPWR _22396_/A sky130_fd_sc_hd__o21ba_1
XFILLER_176_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24103_ _23067_/X _32592_/Q _24105_/S VGND VGND VPWR VPWR _24104_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21315_ _22374_/A VGND VGND VPWR VPWR _21315_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_201_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25083_ _24923_/X _33022_/Q _25101_/S VGND VGND VPWR VPWR _25084_/A sky130_fd_sc_hd__mux2_1
X_29960_ _29960_/A VGND VGND VPWR VPWR _35234_/D sky130_fd_sc_hd__clkbuf_1
X_22295_ _32644_/Q _32580_/Q _32516_/Q _35972_/Q _22229_/X _22013_/X VGND VGND VPWR
+ VPWR _22295_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28911_ _34768_/Q _27214_/X _28913_/S VGND VGND VPWR VPWR _28912_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24034_ _22965_/X _32559_/Q _24042_/S VGND VGND VPWR VPWR _24035_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21246_ _35686_/Q _32193_/Q _35558_/Q _35494_/Q _21211_/X _21212_/X VGND VGND VPWR
+ VPWR _21246_/X sky130_fd_sc_hd__mux4_1
XFILLER_104_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29891_ _35202_/Q _29466_/X _29901_/S VGND VGND VPWR VPWR _29892_/A sky130_fd_sc_hd__mux2_1
XFILLER_176_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28842_ _34735_/Q _27112_/X _28850_/S VGND VGND VPWR VPWR _28843_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21177_ _20961_/X _21175_/X _21176_/X _20965_/X VGND VGND VPWR VPWR _21177_/X sky130_fd_sc_hd__a22o_1
XFILLER_120_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20128_ _20128_/A _20128_/B _20128_/C _20128_/D VGND VGND VPWR VPWR _20129_/A sky130_fd_sc_hd__or4_4
X_28773_ _28773_/A VGND VGND VPWR VPWR _34703_/D sky130_fd_sc_hd__clkbuf_1
X_25985_ _25985_/A VGND VGND VPWR VPWR _33447_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27724_ _27723_/X _34224_/Q _27733_/S VGND VGND VPWR VPWR _27725_/A sky130_fd_sc_hd__mux2_1
X_20059_ _34182_/Q _34118_/Q _34054_/Q _33990_/Q _19746_/X _19747_/X VGND VGND VPWR
+ VPWR _20059_/X sky130_fd_sc_hd__mux4_1
XFILLER_213_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_100_CLK clkbuf_leaf_99_CLK/A VGND VGND VPWR VPWR _33753_/CLK sky130_fd_sc_hd__clkbuf_16
X_24936_ input39/X VGND VGND VPWR VPWR _24936_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_150_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_218_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27655_ input45/X VGND VGND VPWR VPWR _27655_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24867_ _24867_/A VGND VGND VPWR VPWR _32939_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26606_ _24970_/X _33741_/Q _26614_/S VGND VGND VPWR VPWR _26607_/A sky130_fd_sc_hd__mux2_1
XTAP_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23818_ _23049_/X _32394_/Q _23832_/S VGND VGND VPWR VPWR _23819_/A sky130_fd_sc_hd__mux2_1
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24798_ _24798_/A VGND VGND VPWR VPWR _31418_/B sky130_fd_sc_hd__buf_6
X_27586_ _27586_/A VGND VGND VPWR VPWR _34172_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29325_ _29325_/A VGND VGND VPWR VPWR _34964_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26537_ _24868_/X _33708_/Q _26551_/S VGND VGND VPWR VPWR _26538_/A sky130_fd_sc_hd__mux2_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23749_ _23749_/A VGND VGND VPWR VPWR _32361_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17270_ _34168_/Q _34104_/Q _34040_/Q _33976_/Q _17093_/X _17094_/X VGND VGND VPWR
+ VPWR _17270_/X sky130_fd_sc_hd__mux4_1
XFILLER_13_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29256_ _29256_/A VGND VGND VPWR VPWR _34931_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26468_ _33676_/Q _23469_/X _26478_/S VGND VGND VPWR VPWR _26469_/A sky130_fd_sc_hd__mux2_1
XFILLER_202_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28207_ _28207_/A VGND VGND VPWR VPWR _34435_/D sky130_fd_sc_hd__clkbuf_1
X_16221_ _17986_/A VGND VGND VPWR VPWR _16221_/X sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_167_CLK clkbuf_6_30__f_CLK/X VGND VGND VPWR VPWR _35730_/CLK sky130_fd_sc_hd__clkbuf_16
X_25419_ _24815_/X _33179_/Q _25427_/S VGND VGND VPWR VPWR _25420_/A sky130_fd_sc_hd__mux2_1
X_29187_ _34899_/Q _27223_/X _29191_/S VGND VGND VPWR VPWR _29188_/A sky130_fd_sc_hd__mux2_1
X_26399_ _33643_/Q _23296_/X _26415_/S VGND VGND VPWR VPWR _26400_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16152_ _16146_/X _16151_/X _16015_/X VGND VGND VPWR VPWR _16176_/A sky130_fd_sc_hd__o21ba_1
XFILLER_31_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28138_ _28138_/A VGND VGND VPWR VPWR _34402_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16083_ _17716_/A VGND VGND VPWR VPWR _16083_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_154_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28069_ _34370_/Q _27171_/X _28079_/S VGND VGND VPWR VPWR _28070_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19911_ _19656_/X _19909_/X _19910_/X _19659_/X VGND VGND VPWR VPWR _19911_/X sky130_fd_sc_hd__a22o_1
X_30100_ _35301_/Q _29376_/X _30108_/S VGND VGND VPWR VPWR _30101_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31080_ _31080_/A VGND VGND VPWR VPWR _35765_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30031_ _30031_/A VGND VGND VPWR VPWR _35268_/D sky130_fd_sc_hd__clkbuf_1
X_19842_ _19838_/X _19841_/X _19804_/X VGND VGND VPWR VPWR _19850_/C sky130_fd_sc_hd__o21ba_1
XFILLER_3_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19773_ _19458_/X _19771_/X _19772_/X _19463_/X VGND VGND VPWR VPWR _19773_/X sky130_fd_sc_hd__a22o_1
X_16985_ _33392_/Q _33328_/Q _33264_/Q _33200_/Q _16774_/X _16775_/X VGND VGND VPWR
+ VPWR _16985_/X sky130_fd_sc_hd__mux4_1
X_18724_ _33888_/Q _33824_/Q _33760_/Q _36064_/Q _18618_/X _18619_/X VGND VGND VPWR
+ VPWR _18724_/X sky130_fd_sc_hd__mux4_1
X_34770_ _34964_/CLK _34770_/D VGND VGND VPWR VPWR _34770_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31982_ _34918_/CLK _31982_/D VGND VGND VPWR VPWR _31982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_883 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33721_ _35769_/CLK _33721_/D VGND VGND VPWR VPWR _33721_/Q sky130_fd_sc_hd__dfxtp_1
X_18655_ _32606_/Q _32542_/Q _32478_/Q _35934_/Q _18517_/X _18654_/X VGND VGND VPWR
+ VPWR _18655_/X sky130_fd_sc_hd__mux4_1
X_30933_ _35696_/Q input19/X _30939_/S VGND VGND VPWR VPWR _30934_/A sky130_fd_sc_hd__mux2_1
XTAP_4480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17606_ _17351_/X _17604_/X _17605_/X _17354_/X VGND VGND VPWR VPWR _17606_/X sky130_fd_sc_hd__a22o_1
X_33652_ _34101_/CLK _33652_/D VGND VGND VPWR VPWR _33652_/Q sky130_fd_sc_hd__dfxtp_1
X_30864_ _30864_/A VGND VGND VPWR VPWR _35663_/D sky130_fd_sc_hd__clkbuf_1
X_18586_ _32092_/Q _32284_/Q _32348_/Q _35868_/Q _18521_/X _20167_/A VGND VGND VPWR
+ VPWR _18586_/X sky130_fd_sc_hd__mux4_1
XTAP_3790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32603_ _35995_/CLK _32603_/D VGND VGND VPWR VPWR _32603_/Q sky130_fd_sc_hd__dfxtp_1
X_17537_ _35647_/Q _35007_/Q _34367_/Q _33727_/Q _17497_/X _17498_/X VGND VGND VPWR
+ VPWR _17537_/X sky130_fd_sc_hd__mux4_1
XFILLER_17_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33583_ _36080_/CLK _33583_/D VGND VGND VPWR VPWR _33583_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30795_ _30795_/A VGND VGND VPWR VPWR _35630_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35322_ _36026_/CLK _35322_/D VGND VGND VPWR VPWR _35322_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32534_ _36119_/CLK _32534_/D VGND VGND VPWR VPWR _32534_/Q sky130_fd_sc_hd__dfxtp_1
X_17468_ _34685_/Q _34621_/Q _34557_/Q _34493_/Q _17292_/X _17293_/X VGND VGND VPWR
+ VPWR _17468_/X sky130_fd_sc_hd__mux4_1
XFILLER_75_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19207_ _34669_/Q _34605_/Q _34541_/Q _34477_/Q _18886_/X _18887_/X VGND VGND VPWR
+ VPWR _19207_/X sky130_fd_sc_hd__mux4_1
X_35253_ _35446_/CLK _35253_/D VGND VGND VPWR VPWR _35253_/Q sky130_fd_sc_hd__dfxtp_1
X_16419_ _34144_/Q _34080_/Q _34016_/Q _33952_/Q _16387_/X _16388_/X VGND VGND VPWR
+ VPWR _16419_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_158_CLK clkbuf_6_31__f_CLK/X VGND VGND VPWR VPWR _36176_/CLK sky130_fd_sc_hd__clkbuf_16
X_32465_ _36079_/CLK _32465_/D VGND VGND VPWR VPWR _32465_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17399_ _34427_/Q _36155_/Q _34299_/Q _34235_/Q _17229_/X _17230_/X VGND VGND VPWR
+ VPWR _17399_/X sky130_fd_sc_hd__mux4_1
XFILLER_146_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34204_ _36235_/CLK _34204_/D VGND VGND VPWR VPWR _34204_/Q sky130_fd_sc_hd__dfxtp_1
X_31416_ _27837_/X _35925_/Q _31416_/S VGND VGND VPWR VPWR _31417_/A sky130_fd_sc_hd__mux2_1
X_19138_ _35179_/Q _35115_/Q _35051_/Q _32171_/Q _18957_/X _18958_/X VGND VGND VPWR
+ VPWR _19138_/X sky130_fd_sc_hd__mux4_1
XFILLER_160_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35184_ _35377_/CLK _35184_/D VGND VGND VPWR VPWR _35184_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32396_ _35916_/CLK _32396_/D VGND VGND VPWR VPWR _32396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34135_ _34135_/CLK _34135_/D VGND VGND VPWR VPWR _34135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19069_ _19069_/A _19069_/B _19069_/C _19069_/D VGND VGND VPWR VPWR _19070_/A sky130_fd_sc_hd__or4_2
X_31347_ _31416_/S VGND VGND VPWR VPWR _31366_/S sky130_fd_sc_hd__buf_4
XFILLER_133_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_1099 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21100_ _22512_/A VGND VGND VPWR VPWR _21100_/X sky130_fd_sc_hd__buf_4
X_34066_ _34963_/CLK _34066_/D VGND VGND VPWR VPWR _34066_/Q sky130_fd_sc_hd__dfxtp_1
X_22080_ _22433_/A VGND VGND VPWR VPWR _22080_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_133_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31278_ _31278_/A VGND VGND VPWR VPWR _35859_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21031_ _32096_/Q _32288_/Q _32352_/Q _35872_/Q _20821_/X _20962_/X VGND VGND VPWR
+ VPWR _21031_/X sky130_fd_sc_hd__mux4_1
X_33017_ _36025_/CLK _33017_/D VGND VGND VPWR VPWR _33017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30229_ _35362_/Q _29367_/X _30243_/S VGND VGND VPWR VPWR _30230_/A sky130_fd_sc_hd__mux2_1
XFILLER_236_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_330_CLK clkbuf_6_38__f_CLK/X VGND VGND VPWR VPWR _36021_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_113_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34968_ _35609_/CLK _34968_/D VGND VGND VPWR VPWR _34968_/Q sky130_fd_sc_hd__dfxtp_1
X_25770_ _25770_/A VGND VGND VPWR VPWR _33345_/D sky130_fd_sc_hd__clkbuf_1
X_22982_ _22980_/X _32052_/Q _23009_/S VGND VGND VPWR VPWR _22983_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21933_ _21933_/A _21933_/B _21933_/C _21933_/D VGND VGND VPWR VPWR _21934_/A sky130_fd_sc_hd__or4_1
X_24721_ _22974_/X _32882_/Q _24723_/S VGND VGND VPWR VPWR _24722_/A sky130_fd_sc_hd__mux2_1
X_33919_ _35711_/CLK _33919_/D VGND VGND VPWR VPWR _33919_/Q sky130_fd_sc_hd__dfxtp_1
X_34899_ _34963_/CLK _34899_/D VGND VGND VPWR VPWR _34899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24652_ _24652_/A VGND VGND VPWR VPWR _32849_/D sky130_fd_sc_hd__clkbuf_1
X_27440_ _34103_/Q _27137_/X _27452_/S VGND VGND VPWR VPWR _27441_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21864_ _34935_/Q _34871_/Q _34807_/Q _34743_/Q _21760_/X _21761_/X VGND VGND VPWR
+ VPWR _21864_/X sky130_fd_sc_hd__mux4_1
XFILLER_83_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23603_ _23603_/A VGND VGND VPWR VPWR _32293_/D sky130_fd_sc_hd__clkbuf_1
X_20815_ _20747_/X _20813_/X _20814_/X _20750_/X VGND VGND VPWR VPWR _20815_/X sky130_fd_sc_hd__a22o_1
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27371_ _34070_/Q _27033_/X _27389_/S VGND VGND VPWR VPWR _27372_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_397_CLK clkbuf_6_41__f_CLK/X VGND VGND VPWR VPWR _36151_/CLK sky130_fd_sc_hd__clkbuf_16
X_24583_ _24583_/A VGND VGND VPWR VPWR _32816_/D sky130_fd_sc_hd__clkbuf_1
X_21795_ _21758_/X _21793_/X _21794_/X _21763_/X VGND VGND VPWR VPWR _21795_/X sky130_fd_sc_hd__a22o_1
XFILLER_208_1244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29110_ _34862_/Q _27109_/X _29120_/S VGND VGND VPWR VPWR _29111_/A sky130_fd_sc_hd__mux2_1
X_26322_ _26322_/A VGND VGND VPWR VPWR _33607_/D sky130_fd_sc_hd__clkbuf_1
X_23534_ _32262_/Q _23447_/X _23536_/S VGND VGND VPWR VPWR _23535_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20746_ _20740_/X _20743_/X _20744_/X _20745_/X VGND VGND VPWR VPWR _20746_/X sky130_fd_sc_hd__a22o_1
XFILLER_195_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29041_ _29041_/A VGND VGND VPWR VPWR _34829_/D sky130_fd_sc_hd__clkbuf_1
X_26253_ _26253_/A VGND VGND VPWR VPWR _33574_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_149_CLK clkbuf_6_29__f_CLK/X VGND VGND VPWR VPWR _34773_/CLK sky130_fd_sc_hd__clkbuf_16
X_23465_ _23465_/A VGND VGND VPWR VPWR _32233_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20677_ _22365_/A VGND VGND VPWR VPWR _21753_/A sky130_fd_sc_hd__buf_8
XFILLER_183_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25204_ _25204_/A VGND VGND VPWR VPWR _33078_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22416_ _22304_/X _22414_/X _22415_/X _22307_/X VGND VGND VPWR VPWR _22416_/X sky130_fd_sc_hd__a22o_1
X_26184_ _24948_/X _33542_/Q _26186_/S VGND VGND VPWR VPWR _26185_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23396_ input26/X VGND VGND VPWR VPWR _23396_/X sky130_fd_sc_hd__clkbuf_4
X_25135_ _25267_/S VGND VGND VPWR VPWR _25154_/S sky130_fd_sc_hd__buf_6
X_22347_ _22309_/X _22345_/X _22346_/X _22312_/X VGND VGND VPWR VPWR _22347_/X sky130_fd_sc_hd__a22o_1
XFILLER_136_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29943_ _29943_/A VGND VGND VPWR VPWR _35226_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25066_ _24899_/X _33014_/Q _25080_/S VGND VGND VPWR VPWR _25067_/A sky130_fd_sc_hd__mux2_1
X_22278_ _22274_/X _22277_/X _22104_/X VGND VGND VPWR VPWR _22286_/C sky130_fd_sc_hd__o21ba_1
X_24017_ _22940_/X _32551_/Q _24021_/S VGND VGND VPWR VPWR _24018_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21229_ _33638_/Q _33574_/Q _33510_/Q _33446_/Q _21094_/X _21095_/X VGND VGND VPWR
+ VPWR _21229_/X sky130_fd_sc_hd__mux4_1
X_29874_ _35194_/Q _29441_/X _29880_/S VGND VGND VPWR VPWR _29875_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_321_CLK clkbuf_6_39__f_CLK/X VGND VGND VPWR VPWR _32882_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_137_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28825_ _34727_/Q _27087_/X _28829_/S VGND VGND VPWR VPWR _28826_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28756_ _28756_/A VGND VGND VPWR VPWR _34695_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16770_ _16770_/A VGND VGND VPWR VPWR _31977_/D sky130_fd_sc_hd__clkbuf_1
X_25968_ _25968_/A VGND VGND VPWR VPWR _33439_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_991 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27707_ _27707_/A VGND VGND VPWR VPWR _34218_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24919_ _24919_/A VGND VGND VPWR VPWR _32956_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28687_ _28687_/A VGND VGND VPWR VPWR _34662_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1024 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25899_ _25899_/A VGND VGND VPWR VPWR _33406_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_233_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18440_ _20159_/A VGND VGND VPWR VPWR _18440_/X sky130_fd_sc_hd__buf_4
XFILLER_2_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27638_ _27638_/A VGND VGND VPWR VPWR _34197_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18371_ _20077_/A VGND VGND VPWR VPWR _20169_/A sky130_fd_sc_hd__buf_12
XFILLER_15_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27569_ _34164_/Q _27127_/X _27587_/S VGND VGND VPWR VPWR _27570_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_388_CLK clkbuf_6_40__f_CLK/X VGND VGND VPWR VPWR _36090_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29308_ _34956_/Q _27202_/X _29318_/S VGND VGND VPWR VPWR _29309_/A sky130_fd_sc_hd__mux2_1
XFILLER_202_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17322_ _35449_/Q _35385_/Q _35321_/Q _35257_/Q _17254_/X _17255_/X VGND VGND VPWR
+ VPWR _17322_/X sky130_fd_sc_hd__mux4_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_1153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30580_ _30580_/A VGND VGND VPWR VPWR _35528_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17253_ _16998_/X _17251_/X _17252_/X _17001_/X VGND VGND VPWR VPWR _17253_/X sky130_fd_sc_hd__a22o_1
X_29239_ _34923_/Q _27100_/X _29255_/S VGND VGND VPWR VPWR _29240_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16204_ _34393_/Q _36121_/Q _34265_/Q _34201_/Q _16170_/X _16171_/X VGND VGND VPWR
+ VPWR _16204_/X sky130_fd_sc_hd__mux4_1
XFILLER_31_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32250_ _35835_/CLK _32250_/D VGND VGND VPWR VPWR _32250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17184_ _35637_/Q _34997_/Q _34357_/Q _33717_/Q _17144_/X _17145_/X VGND VGND VPWR
+ VPWR _17184_/X sky130_fd_sc_hd__mux4_1
XFILLER_183_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31201_ _31201_/A VGND VGND VPWR VPWR _35822_/D sky130_fd_sc_hd__clkbuf_1
X_16135_ _34903_/Q _34839_/Q _34775_/Q _34711_/Q _16096_/X _16098_/X VGND VGND VPWR
+ VPWR _16135_/X sky130_fd_sc_hd__mux4_1
X_32181_ _35547_/CLK _32181_/D VGND VGND VPWR VPWR _32181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31132_ _31132_/A VGND VGND VPWR VPWR _35790_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16066_ _17982_/A VGND VGND VPWR VPWR _17935_/A sky130_fd_sc_hd__buf_12
XFILLER_29_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_312_CLK clkbuf_6_50__f_CLK/X VGND VGND VPWR VPWR _35975_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_9_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31063_ _31063_/A VGND VGND VPWR VPWR _35757_/D sky130_fd_sc_hd__clkbuf_1
X_35940_ _36007_/CLK _35940_/D VGND VGND VPWR VPWR _35940_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19825_ _33407_/Q _33343_/Q _33279_/Q _33215_/Q _19780_/X _19781_/X VGND VGND VPWR
+ VPWR _19825_/X sky130_fd_sc_hd__mux4_1
XFILLER_123_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30014_ _30014_/A VGND VGND VPWR VPWR _35260_/D sky130_fd_sc_hd__clkbuf_1
X_35871_ _35871_/CLK _35871_/D VGND VGND VPWR VPWR _35871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34822_ _36167_/CLK _34822_/D VGND VGND VPWR VPWR _34822_/Q sky130_fd_sc_hd__dfxtp_1
X_19756_ _19712_/X _19754_/X _19755_/X _19718_/X VGND VGND VPWR VPWR _19756_/X sky130_fd_sc_hd__a22o_1
X_16968_ _16645_/X _16966_/X _16967_/X _16648_/X VGND VGND VPWR VPWR _16968_/X sky130_fd_sc_hd__a22o_1
XFILLER_49_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18707_ _18597_/X _18705_/X _18706_/X _18600_/X VGND VGND VPWR VPWR _18707_/X sky130_fd_sc_hd__a22o_1
X_34753_ _36104_/CLK _34753_/D VGND VGND VPWR VPWR _34753_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_5_16_0_CLK clkbuf_2_2_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_16_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_209_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31965_ _34148_/CLK _31965_/D VGND VGND VPWR VPWR _31965_/Q sky130_fd_sc_hd__dfxtp_1
X_19687_ _19367_/X _19685_/X _19686_/X _19371_/X VGND VGND VPWR VPWR _19687_/X sky130_fd_sc_hd__a22o_1
X_16899_ _35629_/Q _34989_/Q _34349_/Q _33709_/Q _16791_/X _16792_/X VGND VGND VPWR
+ VPWR _16899_/X sky130_fd_sc_hd__mux4_1
XFILLER_65_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33704_ _35559_/CLK _33704_/D VGND VGND VPWR VPWR _33704_/Q sky130_fd_sc_hd__dfxtp_1
X_18638_ _35165_/Q _35101_/Q _35037_/Q _32157_/Q _18604_/X _18605_/X VGND VGND VPWR
+ VPWR _18638_/X sky130_fd_sc_hd__mux4_1
X_30916_ _35688_/Q input10/X _30918_/S VGND VGND VPWR VPWR _30917_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34684_ _35644_/CLK _34684_/D VGND VGND VPWR VPWR _34684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31896_ _23402_/X _36152_/Q _31906_/S VGND VGND VPWR VPWR _31897_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_791 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33635_ _34148_/CLK _33635_/D VGND VGND VPWR VPWR _33635_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18569_ _18378_/X _18567_/X _18568_/X _18388_/X VGND VGND VPWR VPWR _18569_/X sky130_fd_sc_hd__a22o_1
XFILLER_206_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30847_ _30847_/A VGND VGND VPWR VPWR _35655_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_379_CLK clkbuf_6_42__f_CLK/X VGND VGND VPWR VPWR _34172_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_40_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20600_ _22373_/A VGND VGND VPWR VPWR _22464_/A sky130_fd_sc_hd__buf_12
XFILLER_36_1114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33566_ _36191_/CLK _33566_/D VGND VGND VPWR VPWR _33566_/Q sky130_fd_sc_hd__dfxtp_1
X_21580_ _21580_/A _21580_/B _21580_/C _21580_/D VGND VGND VPWR VPWR _21581_/A sky130_fd_sc_hd__or4_4
XFILLER_178_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30778_ _30778_/A VGND VGND VPWR VPWR _35622_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35305_ _35433_/CLK _35305_/D VGND VGND VPWR VPWR _35305_/Q sky130_fd_sc_hd__dfxtp_1
X_32517_ _35973_/CLK _32517_/D VGND VGND VPWR VPWR _32517_/Q sky130_fd_sc_hd__dfxtp_1
X_20531_ _19458_/A _20529_/X _20530_/X _19463_/A VGND VGND VPWR VPWR _20531_/X sky130_fd_sc_hd__a22o_1
XFILLER_32_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33497_ _34009_/CLK _33497_/D VGND VGND VPWR VPWR _33497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23250_ _32156_/Q _23249_/X _23259_/S VGND VGND VPWR VPWR _23251_/A sky130_fd_sc_hd__mux2_1
X_35236_ _35817_/CLK _35236_/D VGND VGND VPWR VPWR _35236_/Q sky130_fd_sc_hd__dfxtp_1
X_20462_ _33426_/Q _33362_/Q _33298_/Q _33234_/Q _18337_/X _18339_/X VGND VGND VPWR
+ VPWR _20462_/X sky130_fd_sc_hd__mux4_1
XFILLER_165_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32448_ _36075_/CLK _32448_/D VGND VGND VPWR VPWR _32448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22201_ _32897_/Q _32833_/Q _32769_/Q _32705_/Q _21946_/X _21947_/X VGND VGND VPWR
+ VPWR _22201_/X sky130_fd_sc_hd__mux4_1
XFILLER_119_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35167_ _35609_/CLK _35167_/D VGND VGND VPWR VPWR _35167_/Q sky130_fd_sc_hd__dfxtp_1
X_23181_ _23181_/A VGND VGND VPWR VPWR _32128_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20393_ _34447_/Q _36175_/Q _34319_/Q _34255_/Q _20235_/X _20236_/X VGND VGND VPWR
+ VPWR _20393_/X sky130_fd_sc_hd__mux4_1
XFILLER_173_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32379_ _32889_/CLK _32379_/D VGND VGND VPWR VPWR _32379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_1237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34118_ _34182_/CLK _34118_/D VGND VGND VPWR VPWR _34118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22132_ _32127_/Q _32319_/Q _32383_/Q _35903_/Q _21880_/X _22021_/X VGND VGND VPWR
+ VPWR _22132_/X sky130_fd_sc_hd__mux4_1
XFILLER_133_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35098_ _35162_/CLK _35098_/D VGND VGND VPWR VPWR _35098_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput230 _32426_/Q VGND VGND VPWR VPWR D3[20] sky130_fd_sc_hd__buf_2
XTAP_6607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput241 _32436_/Q VGND VGND VPWR VPWR D3[30] sky130_fd_sc_hd__buf_2
XFILLER_161_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput252 _32446_/Q VGND VGND VPWR VPWR D3[40] sky130_fd_sc_hd__buf_2
XTAP_6618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34049_ _36159_/CLK _34049_/D VGND VGND VPWR VPWR _34049_/Q sky130_fd_sc_hd__dfxtp_1
X_26940_ _26940_/A VGND VGND VPWR VPWR _33897_/D sky130_fd_sc_hd__clkbuf_1
Xoutput263 _32456_/Q VGND VGND VPWR VPWR D3[50] sky130_fd_sc_hd__buf_2
X_22063_ _21951_/X _22061_/X _22062_/X _21954_/X VGND VGND VPWR VPWR _22063_/X sky130_fd_sc_hd__a22o_1
XFILLER_245_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_303_CLK clkbuf_6_51__f_CLK/X VGND VGND VPWR VPWR _35463_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_161_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput274 _32466_/Q VGND VGND VPWR VPWR D3[60] sky130_fd_sc_hd__buf_2
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21014_ _20691_/X _21012_/X _21013_/X _20701_/X VGND VGND VPWR VPWR _21014_/X sky130_fd_sc_hd__a22o_1
XTAP_5917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26871_ _26871_/A VGND VGND VPWR VPWR _33864_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28610_ _28610_/A VGND VGND VPWR VPWR _34626_/D sky130_fd_sc_hd__clkbuf_1
X_25822_ _24812_/X _33370_/Q _25832_/S VGND VGND VPWR VPWR _25823_/A sky130_fd_sc_hd__mux2_1
XFILLER_134_1279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29590_ _29590_/A VGND VGND VPWR VPWR _35059_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28541_ _28541_/A VGND VGND VPWR VPWR _34593_/D sky130_fd_sc_hd__clkbuf_1
X_25753_ _25753_/A VGND VGND VPWR VPWR _33337_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22965_ input18/X VGND VGND VPWR VPWR _22965_/X sky130_fd_sc_hd__buf_2
XFILLER_216_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_243_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24704_ _24794_/S VGND VGND VPWR VPWR _24723_/S sky130_fd_sc_hd__buf_4
XFILLER_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28472_ _27776_/X _34561_/Q _28484_/S VGND VGND VPWR VPWR _28473_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21916_ _21912_/X _21915_/X _21740_/X _21741_/X VGND VGND VPWR VPWR _21933_/B sky130_fd_sc_hd__o211a_1
X_22896_ _22896_/A VGND VGND VPWR VPWR _32024_/D sky130_fd_sc_hd__clkbuf_1
X_25684_ _25684_/A VGND VGND VPWR VPWR _33304_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27423_ _34095_/Q _27112_/X _27431_/S VGND VGND VPWR VPWR _27424_/A sky130_fd_sc_hd__mux2_1
X_24635_ _23046_/X _32841_/Q _24651_/S VGND VGND VPWR VPWR _24636_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21847_ _32119_/Q _32311_/Q _32375_/Q _35895_/Q _21527_/X _21668_/X VGND VGND VPWR
+ VPWR _21847_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27354_ _27354_/A VGND VGND VPWR VPWR _34062_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24566_ _24566_/A VGND VGND VPWR VPWR _32808_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21778_ _21659_/X _21776_/X _21777_/X _21665_/X VGND VGND VPWR VPWR _21778_/X sky130_fd_sc_hd__a22o_1
XFILLER_168_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26305_ _24927_/X _33599_/Q _26321_/S VGND VGND VPWR VPWR _26306_/A sky130_fd_sc_hd__mux2_1
X_20729_ _20660_/X _20727_/X _20728_/X _20672_/X VGND VGND VPWR VPWR _20729_/X sky130_fd_sc_hd__a22o_1
X_23517_ _23565_/S VGND VGND VPWR VPWR _23536_/S sky130_fd_sc_hd__buf_4
X_24497_ _24524_/S VGND VGND VPWR VPWR _24516_/S sky130_fd_sc_hd__buf_4
X_27285_ _27285_/A VGND VGND VPWR VPWR _34029_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29024_ _29024_/A VGND VGND VPWR VPWR _34821_/D sky130_fd_sc_hd__clkbuf_1
X_23448_ _32228_/Q _23447_/X _23451_/S VGND VGND VPWR VPWR _23449_/A sky130_fd_sc_hd__mux2_1
X_26236_ _26236_/A VGND VGND VPWR VPWR _33566_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_221_1263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26167_ _26215_/S VGND VGND VPWR VPWR _26186_/S sky130_fd_sc_hd__buf_6
X_23379_ _32205_/Q _23364_/X _23385_/S VGND VGND VPWR VPWR _23380_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25118_ _24976_/X _33039_/Q _25122_/S VGND VGND VPWR VPWR _25119_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26098_ _24821_/X _33501_/Q _26102_/S VGND VGND VPWR VPWR _26099_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17940_ _17934_/X _17939_/X _17871_/X VGND VGND VPWR VPWR _17941_/D sky130_fd_sc_hd__o21ba_1
X_29926_ _35219_/Q _29518_/X _29930_/S VGND VGND VPWR VPWR _29927_/A sky130_fd_sc_hd__mux2_1
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25049_ _24874_/X _33006_/Q _25059_/S VGND VGND VPWR VPWR _25050_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17871_ _17871_/A VGND VGND VPWR VPWR _17871_/X sky130_fd_sc_hd__buf_2
XFILLER_120_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29857_ _35186_/Q _29416_/X _29859_/S VGND VGND VPWR VPWR _29858_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19610_ _32633_/Q _32569_/Q _32505_/Q _35961_/Q _19576_/X _19360_/X VGND VGND VPWR
+ VPWR _19610_/X sky130_fd_sc_hd__mux4_1
X_28808_ _34719_/Q _27062_/X _28808_/S VGND VGND VPWR VPWR _28809_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16822_ _16818_/X _16821_/X _16779_/X VGND VGND VPWR VPWR _16844_/A sky130_fd_sc_hd__o21ba_1
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29788_ _29788_/A VGND VGND VPWR VPWR _35153_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19541_ _33911_/Q _33847_/Q _33783_/Q _36087_/Q _19324_/X _19325_/X VGND VGND VPWR
+ VPWR _19541_/X sky130_fd_sc_hd__mux4_1
X_28739_ _34687_/Q _27162_/X _28755_/S VGND VGND VPWR VPWR _28740_/A sky130_fd_sc_hd__mux2_1
X_16753_ _16714_/X _16751_/X _16752_/X _16718_/X VGND VGND VPWR VPWR _16753_/X sky130_fd_sc_hd__a22o_1
XFILLER_235_932 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_588 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31750_ _36083_/Q input22/X _31750_/S VGND VGND VPWR VPWR _31751_/A sky130_fd_sc_hd__mux2_1
X_19472_ _33397_/Q _33333_/Q _33269_/Q _33205_/Q _19427_/X _19428_/X VGND VGND VPWR
+ VPWR _19472_/X sky130_fd_sc_hd__mux4_1
XFILLER_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16684_ _35623_/Q _34983_/Q _34343_/Q _33703_/Q _16438_/X _16439_/X VGND VGND VPWR
+ VPWR _16684_/X sky130_fd_sc_hd__mux4_1
XFILLER_34_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18423_ _18419_/X _18422_/X _18344_/X _18346_/X VGND VGND VPWR VPWR _18438_/B sky130_fd_sc_hd__o211a_1
X_30701_ _35586_/Q _29466_/X _30711_/S VGND VGND VPWR VPWR _30702_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31681_ _31681_/A VGND VGND VPWR VPWR _36050_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33420_ _33420_/CLK _33420_/D VGND VGND VPWR VPWR _33420_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18354_ _20066_/A VGND VGND VPWR VPWR _20299_/A sky130_fd_sc_hd__buf_12
X_30632_ _35553_/Q _29364_/X _30648_/S VGND VGND VPWR VPWR _30633_/A sky130_fd_sc_hd__mux2_1
XFILLER_221_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17305_ _17199_/X _17303_/X _17304_/X _17204_/X VGND VGND VPWR VPWR _17305_/X sky130_fd_sc_hd__a22o_1
XFILLER_203_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33351_ _33415_/CLK _33351_/D VGND VGND VPWR VPWR _33351_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18285_ input78/X VGND VGND VPWR VPWR _18363_/A sky130_fd_sc_hd__buf_6
X_30563_ _30563_/A VGND VGND VPWR VPWR _35520_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32302_ _32877_/CLK _32302_/D VGND VGND VPWR VPWR _32302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36070_ _36070_/CLK _36070_/D VGND VGND VPWR VPWR _36070_/Q sky130_fd_sc_hd__dfxtp_1
X_17236_ _17236_/A VGND VGND VPWR VPWR _31990_/D sky130_fd_sc_hd__clkbuf_1
X_33282_ _36099_/CLK _33282_/D VGND VGND VPWR VPWR _33282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30494_ _30605_/S VGND VGND VPWR VPWR _30513_/S sky130_fd_sc_hd__buf_4
XFILLER_200_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35021_ _35661_/CLK _35021_/D VGND VGND VPWR VPWR _35021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32233_ _35724_/CLK _32233_/D VGND VGND VPWR VPWR _32233_/Q sky130_fd_sc_hd__dfxtp_1
X_17167_ _17167_/A _17167_/B _17167_/C _17167_/D VGND VGND VPWR VPWR _17168_/A sky130_fd_sc_hd__or4_4
XFILLER_143_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_1202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16118_ _33111_/Q _35991_/Q _32983_/Q _32919_/Q _16024_/X _16025_/X VGND VGND VPWR
+ VPWR _16118_/X sky130_fd_sc_hd__mux4_1
XFILLER_127_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32164_ _35168_/CLK _32164_/D VGND VGND VPWR VPWR _32164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17098_ _33907_/Q _33843_/Q _33779_/Q _36083_/Q _17024_/X _17025_/X VGND VGND VPWR
+ VPWR _17098_/X sky130_fd_sc_hd__mux4_1
XFILLER_171_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_817 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31115_ _31115_/A VGND VGND VPWR VPWR _35782_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16049_ _17799_/A VGND VGND VPWR VPWR _16049_/X sky130_fd_sc_hd__buf_6
X_32095_ _35870_/CLK _32095_/D VGND VGND VPWR VPWR _32095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35923_ _35986_/CLK _35923_/D VGND VGND VPWR VPWR _35923_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31046_ _31046_/A VGND VGND VPWR VPWR _35749_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19808_ _35198_/Q _35134_/Q _35070_/Q _32254_/Q _19663_/X _19664_/X VGND VGND VPWR
+ VPWR _19808_/X sky130_fd_sc_hd__mux4_1
XFILLER_84_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35854_ _35855_/CLK _35854_/D VGND VGND VPWR VPWR _35854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34805_ _35829_/CLK _34805_/D VGND VGND VPWR VPWR _34805_/Q sky130_fd_sc_hd__dfxtp_1
X_19739_ _34428_/Q _36156_/Q _34300_/Q _34236_/Q _19529_/X _19530_/X VGND VGND VPWR
+ VPWR _19739_/X sky130_fd_sc_hd__mux4_1
X_35785_ _35785_/CLK _35785_/D VGND VGND VPWR VPWR _35785_/Q sky130_fd_sc_hd__dfxtp_1
X_32997_ _34593_/CLK _32997_/D VGND VGND VPWR VPWR _32997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22750_ _34705_/Q _34641_/Q _34577_/Q _34513_/Q _22598_/X _22599_/X VGND VGND VPWR
+ VPWR _22750_/X sky130_fd_sc_hd__mux4_1
X_31948_ _23484_/X _36177_/Q _31948_/S VGND VGND VPWR VPWR _31949_/A sky130_fd_sc_hd__mux2_1
X_34736_ _34927_/CLK _34736_/D VGND VGND VPWR VPWR _34736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_823 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21701_ _32627_/Q _32563_/Q _32499_/Q _35955_/Q _21523_/X _21660_/X VGND VGND VPWR
+ VPWR _21701_/X sky130_fd_sc_hd__mux4_1
XFILLER_25_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22681_ _22373_/X _22679_/X _22680_/X _22377_/X VGND VGND VPWR VPWR _22681_/X sky130_fd_sc_hd__a22o_1
XFILLER_20_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34667_ _35564_/CLK _34667_/D VGND VGND VPWR VPWR _34667_/Q sky130_fd_sc_hd__dfxtp_1
X_31879_ _23340_/X _36144_/Q _31885_/S VGND VGND VPWR VPWR _31880_/A sky130_fd_sc_hd__mux2_1
X_24420_ _22928_/X _32739_/Q _24432_/S VGND VGND VPWR VPWR _24421_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33618_ _33875_/CLK _33618_/D VGND VGND VPWR VPWR _33618_/Q sky130_fd_sc_hd__dfxtp_1
X_21632_ _32113_/Q _32305_/Q _32369_/Q _35889_/Q _21527_/X _21315_/X VGND VGND VPWR
+ VPWR _21632_/X sky130_fd_sc_hd__mux4_1
XFILLER_40_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34598_ _36135_/CLK _34598_/D VGND VGND VPWR VPWR _34598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24351_ _24351_/A VGND VGND VPWR VPWR _32706_/D sky130_fd_sc_hd__clkbuf_1
X_33549_ _34441_/CLK _33549_/D VGND VGND VPWR VPWR _33549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21563_ _21559_/X _21562_/X _21387_/X _21388_/X VGND VGND VPWR VPWR _21580_/B sky130_fd_sc_hd__o211a_1
XFILLER_240_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23302_ input16/X VGND VGND VPWR VPWR _23302_/X sky130_fd_sc_hd__clkbuf_4
X_20514_ _34963_/Q _34899_/Q _34835_/Q _34771_/Q _18383_/X _18385_/X VGND VGND VPWR
+ VPWR _20514_/X sky130_fd_sc_hd__mux4_1
X_27070_ _33953_/Q _27069_/X _27094_/S VGND VGND VPWR VPWR _27071_/A sky130_fd_sc_hd__mux2_1
X_24282_ _24282_/A VGND VGND VPWR VPWR _32673_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21494_ _32109_/Q _32301_/Q _32365_/Q _35885_/Q _21174_/X _21315_/X VGND VGND VPWR
+ VPWR _21494_/X sky130_fd_sc_hd__mux4_1
XFILLER_14_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23233_ _23233_/A VGND VGND VPWR VPWR _32150_/D sky130_fd_sc_hd__clkbuf_1
X_35219_ _36114_/CLK _35219_/D VGND VGND VPWR VPWR _35219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26021_ _26021_/A VGND VGND VPWR VPWR _33464_/D sky130_fd_sc_hd__clkbuf_1
X_20445_ _18281_/X _20443_/X _20444_/X _18291_/X VGND VGND VPWR VPWR _20445_/X sky130_fd_sc_hd__a22o_1
XFILLER_180_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_238_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36199_ _36202_/CLK _36199_/D VGND VGND VPWR VPWR _36199_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_80_CLK clkbuf_leaf_81_CLK/A VGND VGND VPWR VPWR _36054_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_134_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23164_ _23164_/A VGND VGND VPWR VPWR _32120_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20376_ _32655_/Q _32591_/Q _32527_/Q _35983_/Q _20282_/X _20066_/X VGND VGND VPWR
+ VPWR _20376_/X sky130_fd_sc_hd__mux4_1
XTAP_7116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22115_ _34942_/Q _34878_/Q _34814_/Q _34750_/Q _22113_/X _22114_/X VGND VGND VPWR
+ VPWR _22115_/X sky130_fd_sc_hd__mux4_1
XTAP_6404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27972_ _27972_/A VGND VGND VPWR VPWR _34324_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23095_ _23095_/A VGND VGND VPWR VPWR _32087_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29711_ _29711_/A VGND VGND VPWR VPWR _35116_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26923_ _33889_/Q _23265_/X _26939_/S VGND VGND VPWR VPWR _26924_/A sky130_fd_sc_hd__mux2_1
X_22046_ _22560_/A VGND VGND VPWR VPWR _22046_/X sky130_fd_sc_hd__buf_8
XTAP_6459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29642_ _35084_/Q _29497_/X _29652_/S VGND VGND VPWR VPWR _29643_/A sky130_fd_sc_hd__mux2_1
XTAP_5747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26854_ _26854_/A VGND VGND VPWR VPWR _33856_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25805_ _25805_/A VGND VGND VPWR VPWR _33362_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_229_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29573_ _35051_/Q _29395_/X _29589_/S VGND VGND VPWR VPWR _29574_/A sky130_fd_sc_hd__mux2_1
X_26785_ _26896_/S VGND VGND VPWR VPWR _26804_/S sky130_fd_sc_hd__buf_4
X_23997_ _23997_/A VGND VGND VPWR VPWR _32541_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28524_ _28524_/A VGND VGND VPWR VPWR _34585_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_217_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25736_ _25736_/A VGND VGND VPWR VPWR _33329_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22948_ _22948_/A VGND VGND VPWR VPWR _32041_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28455_ _27751_/X _34553_/Q _28463_/S VGND VGND VPWR VPWR _28456_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25667_ _24982_/X _33297_/Q _25667_/S VGND VGND VPWR VPWR _25668_/A sky130_fd_sc_hd__mux2_1
XFILLER_189_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22879_ input1/X VGND VGND VPWR VPWR _22879_/X sky130_fd_sc_hd__buf_2
X_27406_ _34087_/Q _27087_/X _27410_/S VGND VGND VPWR VPWR _27407_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24618_ _23021_/X _32833_/Q _24630_/S VGND VGND VPWR VPWR _24619_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28386_ _27649_/X _34520_/Q _28400_/S VGND VGND VPWR VPWR _28387_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25598_ _24880_/X _33264_/Q _25604_/S VGND VGND VPWR VPWR _25599_/A sky130_fd_sc_hd__mux2_1
XFILLER_231_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27337_ _27337_/A VGND VGND VPWR VPWR _34054_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_832 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24549_ _22918_/X _32800_/Q _24567_/S VGND VGND VPWR VPWR _24550_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18070_ _34191_/Q _34127_/Q _34063_/Q _33999_/Q _17799_/X _17800_/X VGND VGND VPWR
+ VPWR _18070_/X sky130_fd_sc_hd__mux4_1
XFILLER_157_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27268_ _27268_/A VGND VGND VPWR VPWR _34021_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17021_ _34161_/Q _34097_/Q _34033_/Q _33969_/Q _16740_/X _16741_/X VGND VGND VPWR
+ VPWR _17021_/X sky130_fd_sc_hd__mux4_1
X_29007_ _29007_/A VGND VGND VPWR VPWR _34813_/D sky130_fd_sc_hd__clkbuf_1
X_26219_ _24796_/X _33558_/Q _26237_/S VGND VGND VPWR VPWR _26220_/A sky130_fd_sc_hd__mux2_1
X_27199_ input49/X VGND VGND VPWR VPWR _27199_/X sky130_fd_sc_hd__buf_4
XFILLER_171_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_71_CLK clkbuf_leaf_73_CLK/A VGND VGND VPWR VPWR _35870_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_137_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_952 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18972_ _20151_/A VGND VGND VPWR VPWR _18972_/X sky130_fd_sc_hd__buf_4
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17923_ _17773_/X _17921_/X _17922_/X _17777_/X VGND VGND VPWR VPWR _17923_/X sky130_fd_sc_hd__a22o_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29909_ _29909_/A VGND VGND VPWR VPWR _35210_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32920_ _35992_/CLK _32920_/D VGND VGND VPWR VPWR _32920_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17854_ _35464_/Q _35400_/Q _35336_/Q _35272_/Q _17607_/X _17608_/X VGND VGND VPWR
+ VPWR _17854_/X sky130_fd_sc_hd__mux4_1
XTAP_6993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16805_ _17158_/A VGND VGND VPWR VPWR _16805_/X sky130_fd_sc_hd__clkbuf_4
X_32851_ _35985_/CLK _32851_/D VGND VGND VPWR VPWR _32851_/Q sky130_fd_sc_hd__dfxtp_1
X_17785_ _17936_/A VGND VGND VPWR VPWR _17785_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_130_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31802_ _31802_/A VGND VGND VPWR VPWR _36107_/D sky130_fd_sc_hd__clkbuf_1
X_19524_ _19303_/X _19522_/X _19523_/X _19306_/X VGND VGND VPWR VPWR _19524_/X sky130_fd_sc_hd__a22o_1
X_35570_ _35764_/CLK _35570_/D VGND VGND VPWR VPWR _35570_/Q sky130_fd_sc_hd__dfxtp_1
X_16736_ _16732_/X _16735_/X _16459_/X VGND VGND VPWR VPWR _16737_/D sky130_fd_sc_hd__o21ba_1
XFILLER_75_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32782_ _32913_/CLK _32782_/D VGND VGND VPWR VPWR _32782_/Q sky130_fd_sc_hd__dfxtp_1
X_34521_ _34903_/CLK _34521_/D VGND VGND VPWR VPWR _34521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31733_ _31733_/A VGND VGND VPWR VPWR _36074_/D sky130_fd_sc_hd__clkbuf_1
X_19455_ _35188_/Q _35124_/Q _35060_/Q _32231_/Q _19310_/X _19311_/X VGND VGND VPWR
+ VPWR _19455_/X sky130_fd_sc_hd__mux4_1
X_16667_ _33639_/Q _33575_/Q _33511_/Q _33447_/Q _16494_/X _16495_/X VGND VGND VPWR
+ VPWR _16667_/X sky130_fd_sc_hd__mux4_1
XFILLER_179_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18406_ _18406_/A _18406_/B _18406_/C _18406_/D VGND VGND VPWR VPWR _18407_/A sky130_fd_sc_hd__or4_2
X_34452_ _36180_/CLK _34452_/D VGND VGND VPWR VPWR _34452_/Q sky130_fd_sc_hd__dfxtp_1
X_31664_ _27804_/X _36042_/Q _31678_/S VGND VGND VPWR VPWR _31665_/A sky130_fd_sc_hd__mux2_1
X_19386_ _34418_/Q _36146_/Q _34290_/Q _34226_/Q _19176_/X _19177_/X VGND VGND VPWR
+ VPWR _19386_/X sky130_fd_sc_hd__mux4_1
X_16598_ _34149_/Q _34085_/Q _34021_/Q _33957_/Q _16387_/X _16388_/X VGND VGND VPWR
+ VPWR _16598_/X sky130_fd_sc_hd__mux4_1
XFILLER_188_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33403_ _36092_/CLK _33403_/D VGND VGND VPWR VPWR _33403_/Q sky130_fd_sc_hd__dfxtp_1
X_18337_ _20133_/A VGND VGND VPWR VPWR _18337_/X sky130_fd_sc_hd__clkbuf_8
X_30615_ _35545_/Q _29339_/X _30627_/S VGND VGND VPWR VPWR _30616_/A sky130_fd_sc_hd__mux2_1
XFILLER_188_872 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34383_ _35663_/CLK _34383_/D VGND VGND VPWR VPWR _34383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31595_ _31595_/A VGND VGND VPWR VPWR _36009_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36122_ _36125_/CLK _36122_/D VGND VGND VPWR VPWR _36122_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33334_ _36087_/CLK _33334_/D VGND VGND VPWR VPWR _33334_/Q sky130_fd_sc_hd__dfxtp_1
X_18268_ _16001_/X _18266_/X _18267_/X _16007_/X VGND VGND VPWR VPWR _18268_/X sky130_fd_sc_hd__a22o_1
XFILLER_136_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30546_ _30546_/A VGND VGND VPWR VPWR _35512_/D sky130_fd_sc_hd__clkbuf_1
X_36053_ _36053_/CLK _36053_/D VGND VGND VPWR VPWR _36053_/Q sky130_fd_sc_hd__dfxtp_1
X_17219_ _35702_/Q _32211_/Q _35574_/Q _35510_/Q _16964_/X _16965_/X VGND VGND VPWR
+ VPWR _17219_/X sky130_fd_sc_hd__mux4_1
XFILLER_159_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33265_ _33904_/CLK _33265_/D VGND VGND VPWR VPWR _33265_/Q sky130_fd_sc_hd__dfxtp_1
X_30477_ _30477_/A VGND VGND VPWR VPWR _35479_/D sky130_fd_sc_hd__clkbuf_1
X_18199_ _32147_/Q _32339_/Q _32403_/Q _35923_/Q _17986_/X _17011_/A VGND VGND VPWR
+ VPWR _18199_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_506_CLK clkbuf_leaf_2_CLK/A VGND VGND VPWR VPWR _33573_/CLK sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_62_CLK clkbuf_leaf_65_CLK/A VGND VGND VPWR VPWR _35921_/CLK sky130_fd_sc_hd__clkbuf_16
X_35004_ _35645_/CLK _35004_/D VGND VGND VPWR VPWR _35004_/Q sky130_fd_sc_hd__dfxtp_1
X_20230_ _20009_/X _20228_/X _20229_/X _20012_/X VGND VGND VPWR VPWR _20230_/X sky130_fd_sc_hd__a22o_1
X_32216_ _35709_/CLK _32216_/D VGND VGND VPWR VPWR _32216_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33196_ _36076_/CLK _33196_/D VGND VGND VPWR VPWR _33196_/Q sky130_fd_sc_hd__dfxtp_1
X_20161_ _35208_/Q _35144_/Q _35080_/Q _32264_/Q _20016_/X _20017_/X VGND VGND VPWR
+ VPWR _20161_/X sky130_fd_sc_hd__mux4_1
X_32147_ _35986_/CLK _32147_/D VGND VGND VPWR VPWR _32147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20092_ _34438_/Q _36166_/Q _34310_/Q _34246_/Q _19882_/X _19883_/X VGND VGND VPWR
+ VPWR _20092_/X sky130_fd_sc_hd__mux4_1
X_32078_ _35855_/CLK _32078_/D VGND VGND VPWR VPWR _32078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31029_ _31029_/A VGND VGND VPWR VPWR _35741_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35906_ _35970_/CLK _35906_/D VGND VGND VPWR VPWR _35906_/Q sky130_fd_sc_hd__dfxtp_1
X_23920_ _23920_/A VGND VGND VPWR VPWR _32505_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23851_ _23851_/A VGND VGND VPWR VPWR _32472_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35837_ _36029_/CLK _35837_/D VGND VGND VPWR VPWR _35837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_242_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22802_ _22798_/X _22801_/X _22446_/A _22447_/A VGND VGND VPWR VPWR _22817_/B sky130_fd_sc_hd__o211a_1
X_26570_ _24917_/X _33724_/Q _26572_/S VGND VGND VPWR VPWR _26571_/A sky130_fd_sc_hd__mux2_1
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20994_ _20990_/X _20993_/X _20615_/X VGND VGND VPWR VPWR _21016_/A sky130_fd_sc_hd__o21ba_1
X_35768_ _35768_/CLK _35768_/D VGND VGND VPWR VPWR _35768_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23782_ _22996_/X _32377_/Q _23790_/S VGND VGND VPWR VPWR _23783_/A sky130_fd_sc_hd__mux2_1
X_25521_ _25521_/A VGND VGND VPWR VPWR _33227_/D sky130_fd_sc_hd__clkbuf_1
X_34719_ _34911_/CLK _34719_/D VGND VGND VPWR VPWR _34719_/Q sky130_fd_sc_hd__dfxtp_1
X_22733_ _33937_/Q _33873_/Q _33809_/Q _36113_/Q _20662_/X _20664_/X VGND VGND VPWR
+ VPWR _22733_/X sky130_fd_sc_hd__mux4_1
XFILLER_25_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35699_ _35699_/CLK _35699_/D VGND VGND VPWR VPWR _35699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28240_ _28240_/A VGND VGND VPWR VPWR _34451_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22664_ _34958_/Q _34894_/Q _34830_/Q _34766_/Q _22466_/X _22467_/X VGND VGND VPWR
+ VPWR _22664_/X sky130_fd_sc_hd__mux4_1
XFILLER_197_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25452_ _25452_/A VGND VGND VPWR VPWR _33194_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_240_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24403_ _22903_/X _32731_/Q _24411_/S VGND VGND VPWR VPWR _24404_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21615_ _34928_/Q _34864_/Q _34800_/Q _34736_/Q _21407_/X _21408_/X VGND VGND VPWR
+ VPWR _21615_/X sky130_fd_sc_hd__mux4_1
XFILLER_55_1364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28171_ _28171_/A VGND VGND VPWR VPWR _34418_/D sky130_fd_sc_hd__clkbuf_1
X_22595_ _33100_/Q _32076_/Q _35852_/Q _35788_/Q _22384_/X _22385_/X VGND VGND VPWR
+ VPWR _22595_/X sky130_fd_sc_hd__mux4_1
X_25383_ _33163_/Q _23466_/X _25395_/S VGND VGND VPWR VPWR _25384_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27122_ _33970_/Q _27121_/X _27125_/S VGND VGND VPWR VPWR _27123_/A sky130_fd_sc_hd__mux2_1
X_21546_ _21405_/X _21544_/X _21545_/X _21410_/X VGND VGND VPWR VPWR _21546_/X sky130_fd_sc_hd__a22o_1
X_24334_ _24334_/A VGND VGND VPWR VPWR _32698_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24265_ _24265_/A VGND VGND VPWR VPWR _32665_/D sky130_fd_sc_hd__clkbuf_1
X_27053_ input61/X VGND VGND VPWR VPWR _27053_/X sky130_fd_sc_hd__buf_4
XFILLER_5_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21477_ _21477_/A VGND VGND VPWR VPWR _21477_/X sky130_fd_sc_hd__buf_4
XFILLER_14_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_53_CLK clkbuf_leaf_57_CLK/A VGND VGND VPWR VPWR _32356_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_119_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23216_ _23216_/A VGND VGND VPWR VPWR _32145_/D sky130_fd_sc_hd__clkbuf_1
X_26004_ _26004_/A VGND VGND VPWR VPWR _33456_/D sky130_fd_sc_hd__clkbuf_1
X_20428_ _20428_/A VGND VGND VPWR VPWR _32464_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_153_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24196_ _24196_/A VGND VGND VPWR VPWR _32634_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_901 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23147_ _23147_/A VGND VGND VPWR VPWR _32112_/D sky130_fd_sc_hd__clkbuf_1
X_20359_ _20355_/X _20358_/X _20157_/X VGND VGND VPWR VPWR _20367_/C sky130_fd_sc_hd__o21ba_1
XTAP_6201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27955_ _27810_/X _34316_/Q _27965_/S VGND VGND VPWR VPWR _27956_/A sky130_fd_sc_hd__mux2_1
XTAP_6245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23078_ _23078_/A VGND VGND VPWR VPWR _32083_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26906_ _33881_/Q _23240_/X _26918_/S VGND VGND VPWR VPWR _26907_/A sky130_fd_sc_hd__mux2_1
X_22029_ _21951_/X _22027_/X _22028_/X _21954_/X VGND VGND VPWR VPWR _22029_/X sky130_fd_sc_hd__a22o_1
XTAP_6289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27886_ _27708_/X _34283_/Q _27902_/S VGND VGND VPWR VPWR _27887_/A sky130_fd_sc_hd__mux2_1
XFILLER_212_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29625_ _35076_/Q _29472_/X _29631_/S VGND VGND VPWR VPWR _29626_/A sky130_fd_sc_hd__mux2_1
XTAP_4832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26837_ _26837_/A VGND VGND VPWR VPWR _33848_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17570_ _17420_/X _17568_/X _17569_/X _17424_/X VGND VGND VPWR VPWR _17570_/X sky130_fd_sc_hd__a22o_1
X_29556_ _35043_/Q _29370_/X _29568_/S VGND VGND VPWR VPWR _29557_/A sky130_fd_sc_hd__mux2_1
X_26768_ _26768_/A VGND VGND VPWR VPWR _33815_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28507_ _27828_/X _34578_/Q _28513_/S VGND VGND VPWR VPWR _28508_/A sky130_fd_sc_hd__mux2_1
XFILLER_205_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16521_ _35170_/Q _35106_/Q _35042_/Q _32162_/Q _16304_/X _16305_/X VGND VGND VPWR
+ VPWR _16521_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25719_ _25719_/A VGND VGND VPWR VPWR _33321_/D sky130_fd_sc_hd__clkbuf_1
X_29487_ _29487_/A VGND VGND VPWR VPWR _35016_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26699_ _33783_/Q _23399_/X _26711_/S VGND VGND VPWR VPWR _26700_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19240_ _20299_/A VGND VGND VPWR VPWR _19240_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_232_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28438_ _27726_/X _34545_/Q _28442_/S VGND VGND VPWR VPWR _28439_/A sky130_fd_sc_hd__mux2_1
X_16452_ _17158_/A VGND VGND VPWR VPWR _16452_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_108_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19171_ _18950_/X _19169_/X _19170_/X _18953_/X VGND VGND VPWR VPWR _19171_/X sky130_fd_sc_hd__a22o_1
X_28369_ _28369_/A VGND VGND VPWR VPWR _34512_/D sky130_fd_sc_hd__clkbuf_1
X_16383_ _16379_/X _16382_/X _16104_/X VGND VGND VPWR VPWR _16384_/D sky130_fd_sc_hd__o21ba_2
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18122_ _17859_/X _18120_/X _18121_/X _17862_/X VGND VGND VPWR VPWR _18122_/X sky130_fd_sc_hd__a22o_1
X_30400_ _30400_/A VGND VGND VPWR VPWR _35443_/D sky130_fd_sc_hd__clkbuf_1
XPHY_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31380_ _31380_/A VGND VGND VPWR VPWR _35907_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18053_ _35726_/Q _32237_/Q _35598_/Q _35534_/Q _15993_/X _15995_/X VGND VGND VPWR
+ VPWR _18053_/X sky130_fd_sc_hd__mux4_1
X_30331_ _35411_/Q _29518_/X _30335_/S VGND VGND VPWR VPWR _30332_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_44_CLK clkbuf_6_6__f_CLK/X VGND VGND VPWR VPWR _35943_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_201_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17004_ _35440_/Q _35376_/Q _35312_/Q _35248_/Q _16901_/X _16902_/X VGND VGND VPWR
+ VPWR _17004_/X sky130_fd_sc_hd__mux4_1
X_33050_ _34135_/CLK _33050_/D VGND VGND VPWR VPWR _33050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30262_ _35378_/Q _29416_/X _30264_/S VGND VGND VPWR VPWR _30263_/A sky130_fd_sc_hd__mux2_1
X_32001_ _36207_/CLK _32001_/D VGND VGND VPWR VPWR _32001_/Q sky130_fd_sc_hd__dfxtp_1
X_30193_ _30193_/A VGND VGND VPWR VPWR _35345_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_1240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18955_ _18949_/X _18954_/X _18745_/X VGND VGND VPWR VPWR _18965_/C sky130_fd_sc_hd__o21ba_1
XFILLER_80_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17906_ _17906_/A VGND VGND VPWR VPWR _17906_/X sky130_fd_sc_hd__buf_6
XFILLER_140_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18886_ _20298_/A VGND VGND VPWR VPWR _18886_/X sky130_fd_sc_hd__buf_6
X_33952_ _36202_/CLK _33952_/D VGND VGND VPWR VPWR _33952_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17837_ _17559_/X _17835_/X _17836_/X _17562_/X VGND VGND VPWR VPWR _17837_/X sky130_fd_sc_hd__a22o_1
X_32903_ _32903_/CLK _32903_/D VGND VGND VPWR VPWR _32903_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33883_ _36059_/CLK _33883_/D VGND VGND VPWR VPWR _33883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_212_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32834_ _32894_/CLK _32834_/D VGND VGND VPWR VPWR _32834_/Q sky130_fd_sc_hd__dfxtp_1
X_35622_ _35622_/CLK _35622_/D VGND VGND VPWR VPWR _35622_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17768_ _17986_/A VGND VGND VPWR VPWR _17768_/X sky130_fd_sc_hd__buf_4
XFILLER_214_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_212_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19507_ _33398_/Q _33334_/Q _33270_/Q _33206_/Q _19427_/X _19428_/X VGND VGND VPWR
+ VPWR _19507_/X sky130_fd_sc_hd__mux4_1
X_16719_ _16714_/X _16716_/X _16717_/X _16718_/X VGND VGND VPWR VPWR _16719_/X sky130_fd_sc_hd__a22o_1
X_32765_ _32891_/CLK _32765_/D VGND VGND VPWR VPWR _32765_/Q sky130_fd_sc_hd__dfxtp_1
X_35553_ _35553_/CLK _35553_/D VGND VGND VPWR VPWR _35553_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_6_56__f_CLK clkbuf_5_28_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_56__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_17699_ _17833_/A VGND VGND VPWR VPWR _17699_/X sky130_fd_sc_hd__buf_4
XFILLER_179_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_826 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34504_ _35208_/CLK _34504_/D VGND VGND VPWR VPWR _34504_/Q sky130_fd_sc_hd__dfxtp_1
X_31716_ _31716_/A VGND VGND VPWR VPWR _36066_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19438_ _32884_/Q _32820_/Q _32756_/Q _32692_/Q _19293_/X _19294_/X VGND VGND VPWR
+ VPWR _19438_/X sky130_fd_sc_hd__mux4_1
X_35484_ _36058_/CLK _35484_/D VGND VGND VPWR VPWR _35484_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32696_ _32901_/CLK _32696_/D VGND VGND VPWR VPWR _32696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_245_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34435_ _36163_/CLK _34435_/D VGND VGND VPWR VPWR _34435_/Q sky130_fd_sc_hd__dfxtp_1
X_31647_ _27779_/X _36034_/Q _31657_/S VGND VGND VPWR VPWR _31648_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19369_ _32114_/Q _32306_/Q _32370_/Q _35890_/Q _19227_/X _19368_/X VGND VGND VPWR
+ VPWR _19369_/X sky130_fd_sc_hd__mux4_1
XFILLER_188_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21400_ _21753_/A VGND VGND VPWR VPWR _21400_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_148_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22380_ _35718_/Q _32228_/Q _35590_/Q _35526_/Q _22270_/X _22271_/X VGND VGND VPWR
+ VPWR _22380_/X sky130_fd_sc_hd__mux4_1
X_34366_ _35777_/CLK _34366_/D VGND VGND VPWR VPWR _34366_/Q sky130_fd_sc_hd__dfxtp_1
X_31578_ _27677_/X _36001_/Q _31594_/S VGND VGND VPWR VPWR _31579_/A sky130_fd_sc_hd__mux2_1
XFILLER_191_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36105_ _36105_/CLK _36105_/D VGND VGND VPWR VPWR _36105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33317_ _36068_/CLK _33317_/D VGND VGND VPWR VPWR _33317_/Q sky130_fd_sc_hd__dfxtp_1
X_21331_ _35176_/Q _35112_/Q _35048_/Q _32168_/Q _21257_/X _21258_/X VGND VGND VPWR
+ VPWR _21331_/X sky130_fd_sc_hd__mux4_1
XFILLER_108_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30529_ _30529_/A VGND VGND VPWR VPWR _35504_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34297_ _36152_/CLK _34297_/D VGND VGND VPWR VPWR _34297_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_35_CLK clkbuf_6_7__f_CLK/X VGND VGND VPWR VPWR _36003_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_11_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24050_ _24050_/A VGND VGND VPWR VPWR _32566_/D sky130_fd_sc_hd__clkbuf_1
X_36036_ _36038_/CLK _36036_/D VGND VGND VPWR VPWR _36036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33248_ _36065_/CLK _33248_/D VGND VGND VPWR VPWR _33248_/Q sky130_fd_sc_hd__dfxtp_1
X_21262_ _34918_/Q _34854_/Q _34790_/Q _34726_/Q _21054_/X _21055_/X VGND VGND VPWR
+ VPWR _21262_/X sky130_fd_sc_hd__mux4_1
XFILLER_163_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23001_ _23001_/A VGND VGND VPWR VPWR _32058_/D sky130_fd_sc_hd__clkbuf_1
X_20213_ _33418_/Q _33354_/Q _33290_/Q _33226_/Q _20133_/X _20134_/X VGND VGND VPWR
+ VPWR _20213_/X sky130_fd_sc_hd__mux4_1
XFILLER_11_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33179_ _35547_/CLK _33179_/D VGND VGND VPWR VPWR _33179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21193_ _21052_/X _21191_/X _21192_/X _21057_/X VGND VGND VPWR VPWR _21193_/X sky130_fd_sc_hd__a22o_1
XFILLER_103_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20144_ _32904_/Q _32840_/Q _32776_/Q _32712_/Q _19999_/X _20000_/X VGND VGND VPWR
+ VPWR _20144_/X sky130_fd_sc_hd__mux4_1
XFILLER_58_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27740_ _27739_/X _34229_/Q _27764_/S VGND VGND VPWR VPWR _27741_/A sky130_fd_sc_hd__mux2_1
X_24952_ _24951_/X _32967_/Q _24952_/S VGND VGND VPWR VPWR _24953_/A sky130_fd_sc_hd__mux2_1
XTAP_4106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20075_ _32134_/Q _32326_/Q _32390_/Q _35910_/Q _19933_/X _20074_/X VGND VGND VPWR
+ VPWR _20075_/X sky130_fd_sc_hd__mux4_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23903_ _23903_/A VGND VGND VPWR VPWR _32497_/D sky130_fd_sc_hd__clkbuf_1
X_27671_ _27670_/X _34207_/Q _27671_/S VGND VGND VPWR VPWR _27672_/A sky130_fd_sc_hd__mux2_1
XTAP_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24883_ input20/X VGND VGND VPWR VPWR _24883_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29410_ input19/X VGND VGND VPWR VPWR _29410_/X sky130_fd_sc_hd__buf_2
XFILLER_73_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26622_ _24994_/X _33749_/Q _26622_/S VGND VGND VPWR VPWR _26623_/A sky130_fd_sc_hd__mux2_1
XTAP_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23834_ _23073_/X _32402_/Q _23840_/S VGND VGND VPWR VPWR _23835_/A sky130_fd_sc_hd__mux2_1
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29341_ _29341_/A VGND VGND VPWR VPWR _34969_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26553_ _26622_/S VGND VGND VPWR VPWR _26572_/S sky130_fd_sc_hd__buf_6
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20977_ _34654_/Q _34590_/Q _34526_/Q _34462_/Q _20833_/X _20834_/X VGND VGND VPWR
+ VPWR _20977_/X sky130_fd_sc_hd__mux4_1
XFILLER_57_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23765_ _22971_/X _32369_/Q _23769_/S VGND VGND VPWR VPWR _23766_/A sky130_fd_sc_hd__mux2_1
XFILLER_199_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25504_ _25504_/A VGND VGND VPWR VPWR _33219_/D sky130_fd_sc_hd__clkbuf_1
X_22716_ _35472_/Q _35408_/Q _35344_/Q _35280_/Q _22560_/X _22561_/X VGND VGND VPWR
+ VPWR _22716_/X sky130_fd_sc_hd__mux4_1
XFILLER_13_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29272_ _34939_/Q _27149_/X _29276_/S VGND VGND VPWR VPWR _29273_/A sky130_fd_sc_hd__mux2_1
X_26484_ _33684_/Q _23495_/X _26486_/S VGND VGND VPWR VPWR _26485_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23696_ _23073_/X _32338_/Q _23702_/S VGND VGND VPWR VPWR _23697_/A sky130_fd_sc_hd__mux2_1
X_28223_ _27807_/X _34443_/Q _28235_/S VGND VGND VPWR VPWR _28224_/A sky130_fd_sc_hd__mux2_1
XFILLER_202_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25435_ _25435_/A VGND VGND VPWR VPWR _33186_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22647_ _33166_/Q _36046_/Q _33038_/Q _32974_/Q _22368_/X _22369_/X VGND VGND VPWR
+ VPWR _22647_/X sky130_fd_sc_hd__mux4_1
XFILLER_22_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28154_ _27704_/X _34410_/Q _28172_/S VGND VGND VPWR VPWR _28155_/A sky130_fd_sc_hd__mux2_1
X_22578_ _33420_/Q _33356_/Q _33292_/Q _33228_/Q _22433_/X _22434_/X VGND VGND VPWR
+ VPWR _22578_/X sky130_fd_sc_hd__mux4_1
X_25366_ _33155_/Q _23438_/X _25374_/S VGND VGND VPWR VPWR _25367_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27105_ _27105_/A VGND VGND VPWR VPWR _33964_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24317_ _24317_/A VGND VGND VPWR VPWR _32690_/D sky130_fd_sc_hd__clkbuf_1
X_28085_ _28085_/A VGND VGND VPWR VPWR _34377_/D sky130_fd_sc_hd__clkbuf_1
X_21529_ _32878_/Q _32814_/Q _32750_/Q _32686_/Q _21240_/X _21241_/X VGND VGND VPWR
+ VPWR _21529_/X sky130_fd_sc_hd__mux4_1
X_25297_ _33122_/Q _23268_/X _25311_/S VGND VGND VPWR VPWR _25298_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_26_CLK clkbuf_6_5__f_CLK/X VGND VGND VPWR VPWR _35297_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_154_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27036_ _33942_/Q _27033_/X _27063_/S VGND VGND VPWR VPWR _27037_/A sky130_fd_sc_hd__mux2_1
X_24248_ _24248_/A VGND VGND VPWR VPWR _32659_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24179_ _24179_/A VGND VGND VPWR VPWR _32626_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28987_ _29056_/S VGND VGND VPWR VPWR _29006_/S sky130_fd_sc_hd__buf_4
XTAP_6042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput96 _31973_/Q VGND VGND VPWR VPWR D1[15] sky130_fd_sc_hd__buf_2
XTAP_6064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18740_ _35616_/Q _34976_/Q _34336_/Q _33696_/Q _18738_/X _18739_/X VGND VGND VPWR
+ VPWR _18740_/X sky130_fd_sc_hd__mux4_1
XFILLER_62_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27938_ _27785_/X _34308_/Q _27944_/S VGND VGND VPWR VPWR _27939_/A sky130_fd_sc_hd__mux2_1
XTAP_5330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18671_ _35422_/Q _35358_/Q _35294_/Q _35230_/Q _18495_/X _18496_/X VGND VGND VPWR
+ VPWR _18671_/X sky130_fd_sc_hd__mux4_1
XFILLER_76_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27869_ _27683_/X _34275_/Q _27881_/S VGND VGND VPWR VPWR _27870_/A sky130_fd_sc_hd__mux2_1
XTAP_4651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17622_ _33666_/Q _33602_/Q _33538_/Q _33474_/Q _17553_/X _17554_/X VGND VGND VPWR
+ VPWR _17622_/X sky130_fd_sc_hd__mux4_1
XTAP_4662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_726 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29608_ _35068_/Q _29447_/X _29610_/S VGND VGND VPWR VPWR _29609_/A sky130_fd_sc_hd__mux2_1
X_30880_ _30880_/A VGND VGND VPWR VPWR _35670_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17553_ _17906_/A VGND VGND VPWR VPWR _17553_/X sky130_fd_sc_hd__buf_4
X_29539_ _35035_/Q _29345_/X _29547_/S VGND VGND VPWR VPWR _29540_/A sky130_fd_sc_hd__mux2_1
XTAP_3972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16504_ _16500_/X _16501_/X _16502_/X _16503_/X VGND VGND VPWR VPWR _16504_/X sky130_fd_sc_hd__a22o_1
XFILLER_60_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32550_ _35945_/CLK _32550_/D VGND VGND VPWR VPWR _32550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17484_ _17206_/X _17482_/X _17483_/X _17209_/X VGND VGND VPWR VPWR _17484_/X sky130_fd_sc_hd__a22o_1
XFILLER_177_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19223_ _20282_/A VGND VGND VPWR VPWR _19223_/X sky130_fd_sc_hd__buf_6
X_31501_ _27763_/X _35965_/Q _31501_/S VGND VGND VPWR VPWR _31502_/A sky130_fd_sc_hd__mux2_1
X_16435_ _17847_/A VGND VGND VPWR VPWR _16435_/X sky130_fd_sc_hd__buf_2
XFILLER_108_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32481_ _33119_/CLK _32481_/D VGND VGND VPWR VPWR _32481_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34220_ _34413_/CLK _34220_/D VGND VGND VPWR VPWR _34220_/Q sky130_fd_sc_hd__dfxtp_1
X_31432_ _27661_/X _35932_/Q _31438_/S VGND VGND VPWR VPWR _31433_/A sky130_fd_sc_hd__mux2_1
X_19154_ _33388_/Q _33324_/Q _33260_/Q _33196_/Q _19074_/X _19075_/X VGND VGND VPWR
+ VPWR _19154_/X sky130_fd_sc_hd__mux4_1
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16366_ _16361_/X _16363_/X _16364_/X _16365_/X VGND VGND VPWR VPWR _16366_/X sky130_fd_sc_hd__a22o_1
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18105_ _18101_/X _18104_/X _17838_/X VGND VGND VPWR VPWR _18127_/A sky130_fd_sc_hd__o21ba_2
XFILLER_145_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34151_ _34151_/CLK _34151_/D VGND VGND VPWR VPWR _34151_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19085_ _32874_/Q _32810_/Q _32746_/Q _32682_/Q _18940_/X _18941_/X VGND VGND VPWR
+ VPWR _19085_/X sky130_fd_sc_hd__mux4_1
X_31363_ _31363_/A VGND VGND VPWR VPWR _35899_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_185_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_17_CLK clkbuf_6_6__f_CLK/X VGND VGND VPWR VPWR _35747_/CLK sky130_fd_sc_hd__clkbuf_16
X_16297_ _17864_/A VGND VGND VPWR VPWR _16297_/X sky130_fd_sc_hd__buf_4
XFILLER_199_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33102_ _35853_/CLK _33102_/D VGND VGND VPWR VPWR _33102_/Q sky130_fd_sc_hd__dfxtp_1
X_18036_ _18032_/X _18035_/X _17871_/X VGND VGND VPWR VPWR _18037_/D sky130_fd_sc_hd__o21ba_1
X_30314_ _30314_/A VGND VGND VPWR VPWR _35402_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34082_ _34085_/CLK _34082_/D VGND VGND VPWR VPWR _34082_/Q sky130_fd_sc_hd__dfxtp_1
X_31294_ _31294_/A VGND VGND VPWR VPWR _35866_/D sky130_fd_sc_hd__clkbuf_1
X_33033_ _36042_/CLK _33033_/D VGND VGND VPWR VPWR _33033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30245_ _30335_/S VGND VGND VPWR VPWR _30264_/S sky130_fd_sc_hd__buf_6
XFILLER_67_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30176_ _35337_/Q _29488_/X _30192_/S VGND VGND VPWR VPWR _30177_/A sky130_fd_sc_hd__mux2_1
XFILLER_207_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19987_ _19987_/A VGND VGND VPWR VPWR _32451_/D sky130_fd_sc_hd__buf_2
XFILLER_45_1330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18938_ _18653_/X _18936_/X _18937_/X _18659_/X VGND VGND VPWR VPWR _18938_/X sky130_fd_sc_hd__a22o_1
.ends

