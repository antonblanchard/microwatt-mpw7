magic
tech sky130A
magscale 1 2
timestamp 1662419416
<< obsli1 >>
rect 552 527 234140 19601
<< obsm1 >>
rect 14 8 234140 36848
<< metal2 >>
rect 6274 36688 6330 37088
rect 8022 36688 8078 37088
rect 9770 36688 9826 37088
rect 11518 36688 11574 37088
rect 13266 36688 13322 37088
rect 15014 36688 15070 37088
rect 16762 36688 16818 37088
rect 18510 36688 18566 37088
rect 20258 36688 20314 37088
rect 22006 36688 22062 37088
rect 23754 36688 23810 37088
rect 25502 36688 25558 37088
rect 27250 36688 27306 37088
rect 28998 36688 29054 37088
rect 30746 36688 30802 37088
rect 32494 36688 32550 37088
rect 34242 36688 34298 37088
rect 35990 36688 36046 37088
rect 37738 36688 37794 37088
rect 39486 36688 39542 37088
rect 41234 36688 41290 37088
rect 42982 36688 43038 37088
rect 44730 36688 44786 37088
rect 46478 36688 46534 37088
rect 48226 36688 48282 37088
rect 49974 36688 50030 37088
rect 51722 36688 51778 37088
rect 53470 36688 53526 37088
rect 55218 36688 55274 37088
rect 56966 36688 57022 37088
rect 58714 36688 58770 37088
rect 60462 36688 60518 37088
rect 62210 36688 62266 37088
rect 63958 36688 64014 37088
rect 65706 36688 65762 37088
rect 67454 36688 67510 37088
rect 69202 36688 69258 37088
rect 70950 36688 71006 37088
rect 72698 36688 72754 37088
rect 74446 36688 74502 37088
rect 76194 36688 76250 37088
rect 77942 36688 77998 37088
rect 79690 36688 79746 37088
rect 81438 36688 81494 37088
rect 83186 36688 83242 37088
rect 84934 36688 84990 37088
rect 86682 36688 86738 37088
rect 88430 36688 88486 37088
rect 90178 36688 90234 37088
rect 91926 36688 91982 37088
rect 93674 36688 93730 37088
rect 95422 36688 95478 37088
rect 97170 36688 97226 37088
rect 98918 36688 98974 37088
rect 100666 36688 100722 37088
rect 102414 36688 102470 37088
rect 104162 36688 104218 37088
rect 105910 36688 105966 37088
rect 107658 36688 107714 37088
rect 109406 36688 109462 37088
rect 111154 36688 111210 37088
rect 112902 36688 112958 37088
rect 114650 36688 114706 37088
rect 116398 36688 116454 37088
rect 118146 36688 118202 37088
rect 119894 36688 119950 37088
rect 121642 36688 121698 37088
rect 123390 36688 123446 37088
rect 125138 36688 125194 37088
rect 126886 36688 126942 37088
rect 128634 36688 128690 37088
rect 130382 36688 130438 37088
rect 132130 36688 132186 37088
rect 133878 36688 133934 37088
rect 135626 36688 135682 37088
rect 137374 36688 137430 37088
rect 139122 36688 139178 37088
rect 140870 36688 140926 37088
rect 142618 36688 142674 37088
rect 144366 36688 144422 37088
rect 146114 36688 146170 37088
rect 147862 36688 147918 37088
rect 149610 36688 149666 37088
rect 151358 36688 151414 37088
rect 153106 36688 153162 37088
rect 154854 36688 154910 37088
rect 156602 36688 156658 37088
rect 158350 36688 158406 37088
rect 160098 36688 160154 37088
rect 161846 36688 161902 37088
rect 163594 36688 163650 37088
rect 165342 36688 165398 37088
rect 167090 36688 167146 37088
rect 168838 36688 168894 37088
rect 170586 36688 170642 37088
rect 172334 36688 172390 37088
rect 174082 36688 174138 37088
rect 175830 36688 175886 37088
rect 177578 36688 177634 37088
rect 179326 36688 179382 37088
rect 181074 36688 181130 37088
rect 182822 36688 182878 37088
rect 184570 36688 184626 37088
rect 186318 36688 186374 37088
rect 188066 36688 188122 37088
rect 189814 36688 189870 37088
rect 191562 36688 191618 37088
rect 193310 36688 193366 37088
rect 195058 36688 195114 37088
rect 196806 36688 196862 37088
rect 198554 36688 198610 37088
rect 200302 36688 200358 37088
rect 202050 36688 202106 37088
rect 203798 36688 203854 37088
rect 205546 36688 205602 37088
rect 207294 36688 207350 37088
rect 209042 36688 209098 37088
rect 210790 36688 210846 37088
rect 212538 36688 212594 37088
rect 214286 36688 214342 37088
rect 216034 36688 216090 37088
rect 217782 36688 217838 37088
rect 219530 36688 219586 37088
rect 221278 36688 221334 37088
rect 223026 36688 223082 37088
rect 224774 36688 224830 37088
rect 226522 36688 226578 37088
rect 228270 36688 228326 37088
rect 4250 0 4306 400
rect 7838 0 7894 400
rect 11426 0 11482 400
rect 15014 0 15070 400
rect 18602 0 18658 400
rect 22190 0 22246 400
rect 25778 0 25834 400
rect 29366 0 29422 400
rect 32954 0 33010 400
rect 36542 0 36598 400
rect 40130 0 40186 400
rect 43718 0 43774 400
rect 47306 0 47362 400
rect 50894 0 50950 400
rect 54482 0 54538 400
rect 58070 0 58126 400
rect 61658 0 61714 400
rect 65246 0 65302 400
rect 68834 0 68890 400
rect 72422 0 72478 400
rect 76010 0 76066 400
rect 79598 0 79654 400
rect 83186 0 83242 400
rect 86774 0 86830 400
rect 90362 0 90418 400
rect 93950 0 94006 400
rect 97538 0 97594 400
rect 101126 0 101182 400
rect 104714 0 104770 400
rect 108302 0 108358 400
rect 111890 0 111946 400
rect 115478 0 115534 400
rect 119066 0 119122 400
rect 122654 0 122710 400
rect 126242 0 126298 400
rect 129830 0 129886 400
rect 133418 0 133474 400
rect 137006 0 137062 400
rect 140594 0 140650 400
rect 144182 0 144238 400
rect 147770 0 147826 400
rect 151358 0 151414 400
rect 154946 0 155002 400
rect 158534 0 158590 400
rect 162122 0 162178 400
rect 165710 0 165766 400
rect 169298 0 169354 400
rect 172886 0 172942 400
rect 176474 0 176530 400
rect 180062 0 180118 400
rect 183650 0 183706 400
rect 187238 0 187294 400
rect 190826 0 190882 400
rect 194414 0 194470 400
rect 198002 0 198058 400
rect 201590 0 201646 400
rect 205178 0 205234 400
rect 208766 0 208822 400
rect 212354 0 212410 400
rect 215942 0 215998 400
rect 219530 0 219586 400
rect 223118 0 223174 400
rect 226706 0 226762 400
rect 230294 0 230350 400
<< obsm2 >>
rect 20 36632 6218 36854
rect 6386 36632 7966 36854
rect 8134 36632 9714 36854
rect 9882 36632 11462 36854
rect 11630 36632 13210 36854
rect 13378 36632 14958 36854
rect 15126 36632 16706 36854
rect 16874 36632 18454 36854
rect 18622 36632 20202 36854
rect 20370 36632 21950 36854
rect 22118 36632 23698 36854
rect 23866 36632 25446 36854
rect 25614 36632 27194 36854
rect 27362 36632 28942 36854
rect 29110 36632 30690 36854
rect 30858 36632 32438 36854
rect 32606 36632 34186 36854
rect 34354 36632 35934 36854
rect 36102 36632 37682 36854
rect 37850 36632 39430 36854
rect 39598 36632 41178 36854
rect 41346 36632 42926 36854
rect 43094 36632 44674 36854
rect 44842 36632 46422 36854
rect 46590 36632 48170 36854
rect 48338 36632 49918 36854
rect 50086 36632 51666 36854
rect 51834 36632 53414 36854
rect 53582 36632 55162 36854
rect 55330 36632 56910 36854
rect 57078 36632 58658 36854
rect 58826 36632 60406 36854
rect 60574 36632 62154 36854
rect 62322 36632 63902 36854
rect 64070 36632 65650 36854
rect 65818 36632 67398 36854
rect 67566 36632 69146 36854
rect 69314 36632 70894 36854
rect 71062 36632 72642 36854
rect 72810 36632 74390 36854
rect 74558 36632 76138 36854
rect 76306 36632 77886 36854
rect 78054 36632 79634 36854
rect 79802 36632 81382 36854
rect 81550 36632 83130 36854
rect 83298 36632 84878 36854
rect 85046 36632 86626 36854
rect 86794 36632 88374 36854
rect 88542 36632 90122 36854
rect 90290 36632 91870 36854
rect 92038 36632 93618 36854
rect 93786 36632 95366 36854
rect 95534 36632 97114 36854
rect 97282 36632 98862 36854
rect 99030 36632 100610 36854
rect 100778 36632 102358 36854
rect 102526 36632 104106 36854
rect 104274 36632 105854 36854
rect 106022 36632 107602 36854
rect 107770 36632 109350 36854
rect 109518 36632 111098 36854
rect 111266 36632 112846 36854
rect 113014 36632 114594 36854
rect 114762 36632 116342 36854
rect 116510 36632 118090 36854
rect 118258 36632 119838 36854
rect 120006 36632 121586 36854
rect 121754 36632 123334 36854
rect 123502 36632 125082 36854
rect 125250 36632 126830 36854
rect 126998 36632 128578 36854
rect 128746 36632 130326 36854
rect 130494 36632 132074 36854
rect 132242 36632 133822 36854
rect 133990 36632 135570 36854
rect 135738 36632 137318 36854
rect 137486 36632 139066 36854
rect 139234 36632 140814 36854
rect 140982 36632 142562 36854
rect 142730 36632 144310 36854
rect 144478 36632 146058 36854
rect 146226 36632 147806 36854
rect 147974 36632 149554 36854
rect 149722 36632 151302 36854
rect 151470 36632 153050 36854
rect 153218 36632 154798 36854
rect 154966 36632 156546 36854
rect 156714 36632 158294 36854
rect 158462 36632 160042 36854
rect 160210 36632 161790 36854
rect 161958 36632 163538 36854
rect 163706 36632 165286 36854
rect 165454 36632 167034 36854
rect 167202 36632 168782 36854
rect 168950 36632 170530 36854
rect 170698 36632 172278 36854
rect 172446 36632 174026 36854
rect 174194 36632 175774 36854
rect 175942 36632 177522 36854
rect 177690 36632 179270 36854
rect 179438 36632 181018 36854
rect 181186 36632 182766 36854
rect 182934 36632 184514 36854
rect 184682 36632 186262 36854
rect 186430 36632 188010 36854
rect 188178 36632 189758 36854
rect 189926 36632 191506 36854
rect 191674 36632 193254 36854
rect 193422 36632 195002 36854
rect 195170 36632 196750 36854
rect 196918 36632 198498 36854
rect 198666 36632 200246 36854
rect 200414 36632 201994 36854
rect 202162 36632 203742 36854
rect 203910 36632 205490 36854
rect 205658 36632 207238 36854
rect 207406 36632 208986 36854
rect 209154 36632 210734 36854
rect 210902 36632 212482 36854
rect 212650 36632 214230 36854
rect 214398 36632 215978 36854
rect 216146 36632 217726 36854
rect 217894 36632 219474 36854
rect 219642 36632 221222 36854
rect 221390 36632 222970 36854
rect 223138 36632 224718 36854
rect 224886 36632 226466 36854
rect 226634 36632 228214 36854
rect 228382 36632 233936 36854
rect 20 456 233936 36632
rect 20 2 4194 456
rect 4362 2 7782 456
rect 7950 2 11370 456
rect 11538 2 14958 456
rect 15126 2 18546 456
rect 18714 2 22134 456
rect 22302 2 25722 456
rect 25890 2 29310 456
rect 29478 2 32898 456
rect 33066 2 36486 456
rect 36654 2 40074 456
rect 40242 2 43662 456
rect 43830 2 47250 456
rect 47418 2 50838 456
rect 51006 2 54426 456
rect 54594 2 58014 456
rect 58182 2 61602 456
rect 61770 2 65190 456
rect 65358 2 68778 456
rect 68946 2 72366 456
rect 72534 2 75954 456
rect 76122 2 79542 456
rect 79710 2 83130 456
rect 83298 2 86718 456
rect 86886 2 90306 456
rect 90474 2 93894 456
rect 94062 2 97482 456
rect 97650 2 101070 456
rect 101238 2 104658 456
rect 104826 2 108246 456
rect 108414 2 111834 456
rect 112002 2 115422 456
rect 115590 2 119010 456
rect 119178 2 122598 456
rect 122766 2 126186 456
rect 126354 2 129774 456
rect 129942 2 133362 456
rect 133530 2 136950 456
rect 137118 2 140538 456
rect 140706 2 144126 456
rect 144294 2 147714 456
rect 147882 2 151302 456
rect 151470 2 154890 456
rect 155058 2 158478 456
rect 158646 2 162066 456
rect 162234 2 165654 456
rect 165822 2 169242 456
rect 169410 2 172830 456
rect 172998 2 176418 456
rect 176586 2 180006 456
rect 180174 2 183594 456
rect 183762 2 187182 456
rect 187350 2 190770 456
rect 190938 2 194358 456
rect 194526 2 197946 456
rect 198114 2 201534 456
rect 201702 2 205122 456
rect 205290 2 208710 456
rect 208878 2 212298 456
rect 212466 2 215886 456
rect 216054 2 219474 456
rect 219642 2 223062 456
rect 223230 2 226650 456
rect 226818 2 230238 456
rect 230406 2 233936 456
<< metal3 >>
rect 234292 35232 234692 35352
rect 0 34416 400 34536
rect 234292 32648 234692 32768
rect 234292 30064 234692 30184
rect 0 29112 400 29232
rect 234292 27480 234692 27600
rect 234292 24896 234692 25016
rect 0 23808 400 23928
rect 234292 22312 234692 22432
rect 234292 19728 234692 19848
rect 0 18504 400 18624
rect 234292 17144 234692 17264
rect 234292 14560 234692 14680
rect 0 13200 400 13320
rect 234292 11976 234692 12096
rect 234292 9392 234692 9512
rect 0 7896 400 8016
rect 234292 6808 234692 6928
rect 234292 4224 234692 4344
rect 0 2592 400 2712
rect 234292 1640 234692 1760
<< obsm3 >>
rect 197 35432 234292 36481
rect 197 35152 234212 35432
rect 197 34616 234292 35152
rect 480 34336 234292 34616
rect 197 32848 234292 34336
rect 197 32568 234212 32848
rect 197 30264 234292 32568
rect 197 29984 234212 30264
rect 197 29312 234292 29984
rect 480 29032 234292 29312
rect 197 27680 234292 29032
rect 197 27400 234212 27680
rect 197 25096 234292 27400
rect 197 24816 234212 25096
rect 197 24008 234292 24816
rect 480 23728 234292 24008
rect 197 22512 234292 23728
rect 197 22232 234212 22512
rect 197 19928 234292 22232
rect 197 19648 234212 19928
rect 197 18704 234292 19648
rect 480 18424 234292 18704
rect 197 17344 234292 18424
rect 197 17064 234212 17344
rect 197 14760 234292 17064
rect 197 14480 234212 14760
rect 197 13400 234292 14480
rect 480 13120 234292 13400
rect 197 12176 234292 13120
rect 197 11896 234212 12176
rect 197 9592 234292 11896
rect 197 9312 234212 9592
rect 197 8096 234292 9312
rect 480 7816 234292 8096
rect 197 7008 234292 7816
rect 197 6728 234212 7008
rect 197 4424 234292 6728
rect 197 4144 234212 4424
rect 197 2792 234292 4144
rect 480 2512 234292 2792
rect 197 1840 234292 2512
rect 197 1560 234212 1840
rect 197 35 234292 1560
<< metal4 >>
rect 1242 496 1862 36496
rect 19242 496 19862 36496
rect 37242 496 37862 36496
rect 55242 496 55862 36496
rect 73242 496 73862 36496
rect 91242 496 91862 36496
rect 109242 496 109862 36496
rect 127242 496 127862 36496
rect 145242 496 145862 36496
rect 163242 496 163862 36496
rect 181242 496 181862 36496
rect 199242 496 199862 36496
rect 217242 496 217862 36496
<< obsm4 >>
rect 795 987 1162 35053
rect 1942 987 19162 35053
rect 19942 987 37162 35053
rect 37942 987 55162 35053
rect 55942 987 73162 35053
rect 73942 987 91162 35053
rect 91942 987 109162 35053
rect 109942 987 127162 35053
rect 127942 987 145162 35053
rect 145942 987 163162 35053
rect 163942 987 181162 35053
rect 181942 987 199162 35053
rect 199942 987 214117 35053
<< labels >>
rlabel metal3 s 234292 24896 234692 25016 6 A0[0]
port 1 nsew signal input
rlabel metal3 s 234292 27480 234692 27600 6 A0[1]
port 2 nsew signal input
rlabel metal3 s 234292 30064 234692 30184 6 A0[2]
port 3 nsew signal input
rlabel metal3 s 234292 32648 234692 32768 6 A0[3]
port 4 nsew signal input
rlabel metal3 s 234292 35232 234692 35352 6 A0[4]
port 5 nsew signal input
rlabel metal3 s 0 7896 400 8016 6 A1[0]
port 6 nsew signal input
rlabel metal3 s 0 13200 400 13320 6 A1[1]
port 7 nsew signal input
rlabel metal3 s 0 18504 400 18624 6 A1[2]
port 8 nsew signal input
rlabel metal3 s 0 23808 400 23928 6 A1[3]
port 9 nsew signal input
rlabel metal3 s 0 29112 400 29232 6 A1[4]
port 10 nsew signal input
rlabel metal3 s 0 2592 400 2712 6 CLK
port 11 nsew signal input
rlabel metal2 s 4250 0 4306 400 6 Di0[0]
port 12 nsew signal input
rlabel metal2 s 40130 0 40186 400 6 Di0[10]
port 13 nsew signal input
rlabel metal2 s 43718 0 43774 400 6 Di0[11]
port 14 nsew signal input
rlabel metal2 s 47306 0 47362 400 6 Di0[12]
port 15 nsew signal input
rlabel metal2 s 50894 0 50950 400 6 Di0[13]
port 16 nsew signal input
rlabel metal2 s 54482 0 54538 400 6 Di0[14]
port 17 nsew signal input
rlabel metal2 s 58070 0 58126 400 6 Di0[15]
port 18 nsew signal input
rlabel metal2 s 61658 0 61714 400 6 Di0[16]
port 19 nsew signal input
rlabel metal2 s 65246 0 65302 400 6 Di0[17]
port 20 nsew signal input
rlabel metal2 s 68834 0 68890 400 6 Di0[18]
port 21 nsew signal input
rlabel metal2 s 72422 0 72478 400 6 Di0[19]
port 22 nsew signal input
rlabel metal2 s 7838 0 7894 400 6 Di0[1]
port 23 nsew signal input
rlabel metal2 s 76010 0 76066 400 6 Di0[20]
port 24 nsew signal input
rlabel metal2 s 79598 0 79654 400 6 Di0[21]
port 25 nsew signal input
rlabel metal2 s 83186 0 83242 400 6 Di0[22]
port 26 nsew signal input
rlabel metal2 s 86774 0 86830 400 6 Di0[23]
port 27 nsew signal input
rlabel metal2 s 90362 0 90418 400 6 Di0[24]
port 28 nsew signal input
rlabel metal2 s 93950 0 94006 400 6 Di0[25]
port 29 nsew signal input
rlabel metal2 s 97538 0 97594 400 6 Di0[26]
port 30 nsew signal input
rlabel metal2 s 101126 0 101182 400 6 Di0[27]
port 31 nsew signal input
rlabel metal2 s 104714 0 104770 400 6 Di0[28]
port 32 nsew signal input
rlabel metal2 s 108302 0 108358 400 6 Di0[29]
port 33 nsew signal input
rlabel metal2 s 11426 0 11482 400 6 Di0[2]
port 34 nsew signal input
rlabel metal2 s 111890 0 111946 400 6 Di0[30]
port 35 nsew signal input
rlabel metal2 s 115478 0 115534 400 6 Di0[31]
port 36 nsew signal input
rlabel metal2 s 119066 0 119122 400 6 Di0[32]
port 37 nsew signal input
rlabel metal2 s 122654 0 122710 400 6 Di0[33]
port 38 nsew signal input
rlabel metal2 s 126242 0 126298 400 6 Di0[34]
port 39 nsew signal input
rlabel metal2 s 129830 0 129886 400 6 Di0[35]
port 40 nsew signal input
rlabel metal2 s 133418 0 133474 400 6 Di0[36]
port 41 nsew signal input
rlabel metal2 s 137006 0 137062 400 6 Di0[37]
port 42 nsew signal input
rlabel metal2 s 140594 0 140650 400 6 Di0[38]
port 43 nsew signal input
rlabel metal2 s 144182 0 144238 400 6 Di0[39]
port 44 nsew signal input
rlabel metal2 s 15014 0 15070 400 6 Di0[3]
port 45 nsew signal input
rlabel metal2 s 147770 0 147826 400 6 Di0[40]
port 46 nsew signal input
rlabel metal2 s 151358 0 151414 400 6 Di0[41]
port 47 nsew signal input
rlabel metal2 s 154946 0 155002 400 6 Di0[42]
port 48 nsew signal input
rlabel metal2 s 158534 0 158590 400 6 Di0[43]
port 49 nsew signal input
rlabel metal2 s 162122 0 162178 400 6 Di0[44]
port 50 nsew signal input
rlabel metal2 s 165710 0 165766 400 6 Di0[45]
port 51 nsew signal input
rlabel metal2 s 169298 0 169354 400 6 Di0[46]
port 52 nsew signal input
rlabel metal2 s 172886 0 172942 400 6 Di0[47]
port 53 nsew signal input
rlabel metal2 s 176474 0 176530 400 6 Di0[48]
port 54 nsew signal input
rlabel metal2 s 180062 0 180118 400 6 Di0[49]
port 55 nsew signal input
rlabel metal2 s 18602 0 18658 400 6 Di0[4]
port 56 nsew signal input
rlabel metal2 s 183650 0 183706 400 6 Di0[50]
port 57 nsew signal input
rlabel metal2 s 187238 0 187294 400 6 Di0[51]
port 58 nsew signal input
rlabel metal2 s 190826 0 190882 400 6 Di0[52]
port 59 nsew signal input
rlabel metal2 s 194414 0 194470 400 6 Di0[53]
port 60 nsew signal input
rlabel metal2 s 198002 0 198058 400 6 Di0[54]
port 61 nsew signal input
rlabel metal2 s 201590 0 201646 400 6 Di0[55]
port 62 nsew signal input
rlabel metal2 s 205178 0 205234 400 6 Di0[56]
port 63 nsew signal input
rlabel metal2 s 208766 0 208822 400 6 Di0[57]
port 64 nsew signal input
rlabel metal2 s 212354 0 212410 400 6 Di0[58]
port 65 nsew signal input
rlabel metal2 s 215942 0 215998 400 6 Di0[59]
port 66 nsew signal input
rlabel metal2 s 22190 0 22246 400 6 Di0[5]
port 67 nsew signal input
rlabel metal2 s 219530 0 219586 400 6 Di0[60]
port 68 nsew signal input
rlabel metal2 s 223118 0 223174 400 6 Di0[61]
port 69 nsew signal input
rlabel metal2 s 226706 0 226762 400 6 Di0[62]
port 70 nsew signal input
rlabel metal2 s 230294 0 230350 400 6 Di0[63]
port 71 nsew signal input
rlabel metal2 s 25778 0 25834 400 6 Di0[6]
port 72 nsew signal input
rlabel metal2 s 29366 0 29422 400 6 Di0[7]
port 73 nsew signal input
rlabel metal2 s 32954 0 33010 400 6 Di0[8]
port 74 nsew signal input
rlabel metal2 s 36542 0 36598 400 6 Di0[9]
port 75 nsew signal input
rlabel metal2 s 6274 36688 6330 37088 6 Do0[0]
port 76 nsew signal output
rlabel metal2 s 23754 36688 23810 37088 6 Do0[10]
port 77 nsew signal output
rlabel metal2 s 27250 36688 27306 37088 6 Do0[11]
port 78 nsew signal output
rlabel metal2 s 30746 36688 30802 37088 6 Do0[12]
port 79 nsew signal output
rlabel metal2 s 34242 36688 34298 37088 6 Do0[13]
port 80 nsew signal output
rlabel metal2 s 37738 36688 37794 37088 6 Do0[14]
port 81 nsew signal output
rlabel metal2 s 41234 36688 41290 37088 6 Do0[15]
port 82 nsew signal output
rlabel metal2 s 44730 36688 44786 37088 6 Do0[16]
port 83 nsew signal output
rlabel metal2 s 48226 36688 48282 37088 6 Do0[17]
port 84 nsew signal output
rlabel metal2 s 51722 36688 51778 37088 6 Do0[18]
port 85 nsew signal output
rlabel metal2 s 55218 36688 55274 37088 6 Do0[19]
port 86 nsew signal output
rlabel metal2 s 8022 36688 8078 37088 6 Do0[1]
port 87 nsew signal output
rlabel metal2 s 58714 36688 58770 37088 6 Do0[20]
port 88 nsew signal output
rlabel metal2 s 60462 36688 60518 37088 6 Do0[21]
port 89 nsew signal output
rlabel metal2 s 62210 36688 62266 37088 6 Do0[22]
port 90 nsew signal output
rlabel metal2 s 63958 36688 64014 37088 6 Do0[23]
port 91 nsew signal output
rlabel metal2 s 65706 36688 65762 37088 6 Do0[24]
port 92 nsew signal output
rlabel metal2 s 67454 36688 67510 37088 6 Do0[25]
port 93 nsew signal output
rlabel metal2 s 69202 36688 69258 37088 6 Do0[26]
port 94 nsew signal output
rlabel metal2 s 70950 36688 71006 37088 6 Do0[27]
port 95 nsew signal output
rlabel metal2 s 72698 36688 72754 37088 6 Do0[28]
port 96 nsew signal output
rlabel metal2 s 74446 36688 74502 37088 6 Do0[29]
port 97 nsew signal output
rlabel metal2 s 9770 36688 9826 37088 6 Do0[2]
port 98 nsew signal output
rlabel metal2 s 76194 36688 76250 37088 6 Do0[30]
port 99 nsew signal output
rlabel metal2 s 77942 36688 77998 37088 6 Do0[31]
port 100 nsew signal output
rlabel metal2 s 79690 36688 79746 37088 6 Do0[32]
port 101 nsew signal output
rlabel metal2 s 81438 36688 81494 37088 6 Do0[33]
port 102 nsew signal output
rlabel metal2 s 83186 36688 83242 37088 6 Do0[34]
port 103 nsew signal output
rlabel metal2 s 84934 36688 84990 37088 6 Do0[35]
port 104 nsew signal output
rlabel metal2 s 86682 36688 86738 37088 6 Do0[36]
port 105 nsew signal output
rlabel metal2 s 88430 36688 88486 37088 6 Do0[37]
port 106 nsew signal output
rlabel metal2 s 90178 36688 90234 37088 6 Do0[38]
port 107 nsew signal output
rlabel metal2 s 91926 36688 91982 37088 6 Do0[39]
port 108 nsew signal output
rlabel metal2 s 11518 36688 11574 37088 6 Do0[3]
port 109 nsew signal output
rlabel metal2 s 93674 36688 93730 37088 6 Do0[40]
port 110 nsew signal output
rlabel metal2 s 95422 36688 95478 37088 6 Do0[41]
port 111 nsew signal output
rlabel metal2 s 97170 36688 97226 37088 6 Do0[42]
port 112 nsew signal output
rlabel metal2 s 98918 36688 98974 37088 6 Do0[43]
port 113 nsew signal output
rlabel metal2 s 100666 36688 100722 37088 6 Do0[44]
port 114 nsew signal output
rlabel metal2 s 102414 36688 102470 37088 6 Do0[45]
port 115 nsew signal output
rlabel metal2 s 104162 36688 104218 37088 6 Do0[46]
port 116 nsew signal output
rlabel metal2 s 105910 36688 105966 37088 6 Do0[47]
port 117 nsew signal output
rlabel metal2 s 107658 36688 107714 37088 6 Do0[48]
port 118 nsew signal output
rlabel metal2 s 109406 36688 109462 37088 6 Do0[49]
port 119 nsew signal output
rlabel metal2 s 13266 36688 13322 37088 6 Do0[4]
port 120 nsew signal output
rlabel metal2 s 111154 36688 111210 37088 6 Do0[50]
port 121 nsew signal output
rlabel metal2 s 112902 36688 112958 37088 6 Do0[51]
port 122 nsew signal output
rlabel metal2 s 114650 36688 114706 37088 6 Do0[52]
port 123 nsew signal output
rlabel metal2 s 116398 36688 116454 37088 6 Do0[53]
port 124 nsew signal output
rlabel metal2 s 118146 36688 118202 37088 6 Do0[54]
port 125 nsew signal output
rlabel metal2 s 119894 36688 119950 37088 6 Do0[55]
port 126 nsew signal output
rlabel metal2 s 121642 36688 121698 37088 6 Do0[56]
port 127 nsew signal output
rlabel metal2 s 123390 36688 123446 37088 6 Do0[57]
port 128 nsew signal output
rlabel metal2 s 125138 36688 125194 37088 6 Do0[58]
port 129 nsew signal output
rlabel metal2 s 126886 36688 126942 37088 6 Do0[59]
port 130 nsew signal output
rlabel metal2 s 15014 36688 15070 37088 6 Do0[5]
port 131 nsew signal output
rlabel metal2 s 128634 36688 128690 37088 6 Do0[60]
port 132 nsew signal output
rlabel metal2 s 130382 36688 130438 37088 6 Do0[61]
port 133 nsew signal output
rlabel metal2 s 132130 36688 132186 37088 6 Do0[62]
port 134 nsew signal output
rlabel metal2 s 133878 36688 133934 37088 6 Do0[63]
port 135 nsew signal output
rlabel metal2 s 16762 36688 16818 37088 6 Do0[6]
port 136 nsew signal output
rlabel metal2 s 18510 36688 18566 37088 6 Do0[7]
port 137 nsew signal output
rlabel metal2 s 20258 36688 20314 37088 6 Do0[8]
port 138 nsew signal output
rlabel metal2 s 22006 36688 22062 37088 6 Do0[9]
port 139 nsew signal output
rlabel metal2 s 25502 36688 25558 37088 6 Do1[0]
port 140 nsew signal output
rlabel metal2 s 135626 36688 135682 37088 6 Do1[10]
port 141 nsew signal output
rlabel metal2 s 137374 36688 137430 37088 6 Do1[11]
port 142 nsew signal output
rlabel metal2 s 139122 36688 139178 37088 6 Do1[12]
port 143 nsew signal output
rlabel metal2 s 140870 36688 140926 37088 6 Do1[13]
port 144 nsew signal output
rlabel metal2 s 142618 36688 142674 37088 6 Do1[14]
port 145 nsew signal output
rlabel metal2 s 144366 36688 144422 37088 6 Do1[15]
port 146 nsew signal output
rlabel metal2 s 146114 36688 146170 37088 6 Do1[16]
port 147 nsew signal output
rlabel metal2 s 147862 36688 147918 37088 6 Do1[17]
port 148 nsew signal output
rlabel metal2 s 149610 36688 149666 37088 6 Do1[18]
port 149 nsew signal output
rlabel metal2 s 151358 36688 151414 37088 6 Do1[19]
port 150 nsew signal output
rlabel metal2 s 28998 36688 29054 37088 6 Do1[1]
port 151 nsew signal output
rlabel metal2 s 153106 36688 153162 37088 6 Do1[20]
port 152 nsew signal output
rlabel metal2 s 154854 36688 154910 37088 6 Do1[21]
port 153 nsew signal output
rlabel metal2 s 156602 36688 156658 37088 6 Do1[22]
port 154 nsew signal output
rlabel metal2 s 158350 36688 158406 37088 6 Do1[23]
port 155 nsew signal output
rlabel metal2 s 160098 36688 160154 37088 6 Do1[24]
port 156 nsew signal output
rlabel metal2 s 161846 36688 161902 37088 6 Do1[25]
port 157 nsew signal output
rlabel metal2 s 163594 36688 163650 37088 6 Do1[26]
port 158 nsew signal output
rlabel metal2 s 165342 36688 165398 37088 6 Do1[27]
port 159 nsew signal output
rlabel metal2 s 167090 36688 167146 37088 6 Do1[28]
port 160 nsew signal output
rlabel metal2 s 168838 36688 168894 37088 6 Do1[29]
port 161 nsew signal output
rlabel metal2 s 32494 36688 32550 37088 6 Do1[2]
port 162 nsew signal output
rlabel metal2 s 170586 36688 170642 37088 6 Do1[30]
port 163 nsew signal output
rlabel metal2 s 172334 36688 172390 37088 6 Do1[31]
port 164 nsew signal output
rlabel metal2 s 174082 36688 174138 37088 6 Do1[32]
port 165 nsew signal output
rlabel metal2 s 175830 36688 175886 37088 6 Do1[33]
port 166 nsew signal output
rlabel metal2 s 177578 36688 177634 37088 6 Do1[34]
port 167 nsew signal output
rlabel metal2 s 179326 36688 179382 37088 6 Do1[35]
port 168 nsew signal output
rlabel metal2 s 181074 36688 181130 37088 6 Do1[36]
port 169 nsew signal output
rlabel metal2 s 182822 36688 182878 37088 6 Do1[37]
port 170 nsew signal output
rlabel metal2 s 184570 36688 184626 37088 6 Do1[38]
port 171 nsew signal output
rlabel metal2 s 186318 36688 186374 37088 6 Do1[39]
port 172 nsew signal output
rlabel metal2 s 35990 36688 36046 37088 6 Do1[3]
port 173 nsew signal output
rlabel metal2 s 188066 36688 188122 37088 6 Do1[40]
port 174 nsew signal output
rlabel metal2 s 189814 36688 189870 37088 6 Do1[41]
port 175 nsew signal output
rlabel metal2 s 191562 36688 191618 37088 6 Do1[42]
port 176 nsew signal output
rlabel metal2 s 193310 36688 193366 37088 6 Do1[43]
port 177 nsew signal output
rlabel metal2 s 195058 36688 195114 37088 6 Do1[44]
port 178 nsew signal output
rlabel metal2 s 196806 36688 196862 37088 6 Do1[45]
port 179 nsew signal output
rlabel metal2 s 198554 36688 198610 37088 6 Do1[46]
port 180 nsew signal output
rlabel metal2 s 200302 36688 200358 37088 6 Do1[47]
port 181 nsew signal output
rlabel metal2 s 202050 36688 202106 37088 6 Do1[48]
port 182 nsew signal output
rlabel metal2 s 203798 36688 203854 37088 6 Do1[49]
port 183 nsew signal output
rlabel metal2 s 39486 36688 39542 37088 6 Do1[4]
port 184 nsew signal output
rlabel metal2 s 205546 36688 205602 37088 6 Do1[50]
port 185 nsew signal output
rlabel metal2 s 207294 36688 207350 37088 6 Do1[51]
port 186 nsew signal output
rlabel metal2 s 209042 36688 209098 37088 6 Do1[52]
port 187 nsew signal output
rlabel metal2 s 210790 36688 210846 37088 6 Do1[53]
port 188 nsew signal output
rlabel metal2 s 212538 36688 212594 37088 6 Do1[54]
port 189 nsew signal output
rlabel metal2 s 214286 36688 214342 37088 6 Do1[55]
port 190 nsew signal output
rlabel metal2 s 216034 36688 216090 37088 6 Do1[56]
port 191 nsew signal output
rlabel metal2 s 217782 36688 217838 37088 6 Do1[57]
port 192 nsew signal output
rlabel metal2 s 219530 36688 219586 37088 6 Do1[58]
port 193 nsew signal output
rlabel metal2 s 221278 36688 221334 37088 6 Do1[59]
port 194 nsew signal output
rlabel metal2 s 42982 36688 43038 37088 6 Do1[5]
port 195 nsew signal output
rlabel metal2 s 223026 36688 223082 37088 6 Do1[60]
port 196 nsew signal output
rlabel metal2 s 224774 36688 224830 37088 6 Do1[61]
port 197 nsew signal output
rlabel metal2 s 226522 36688 226578 37088 6 Do1[62]
port 198 nsew signal output
rlabel metal2 s 228270 36688 228326 37088 6 Do1[63]
port 199 nsew signal output
rlabel metal2 s 46478 36688 46534 37088 6 Do1[6]
port 200 nsew signal output
rlabel metal2 s 49974 36688 50030 37088 6 Do1[7]
port 201 nsew signal output
rlabel metal2 s 53470 36688 53526 37088 6 Do1[8]
port 202 nsew signal output
rlabel metal2 s 56966 36688 57022 37088 6 Do1[9]
port 203 nsew signal output
rlabel metal3 s 234292 1640 234692 1760 6 EN0
port 204 nsew signal input
rlabel metal3 s 0 34416 400 34536 6 EN1
port 205 nsew signal input
rlabel metal4 s 19242 496 19862 36496 6 VGND
port 206 nsew ground bidirectional
rlabel metal4 s 55242 496 55862 36496 6 VGND
port 206 nsew ground bidirectional
rlabel metal4 s 91242 496 91862 36496 6 VGND
port 206 nsew ground bidirectional
rlabel metal4 s 127242 496 127862 36496 6 VGND
port 206 nsew ground bidirectional
rlabel metal4 s 163242 496 163862 36496 6 VGND
port 206 nsew ground bidirectional
rlabel metal4 s 199242 496 199862 36496 6 VGND
port 206 nsew ground bidirectional
rlabel metal4 s 1242 496 1862 36496 6 VPWR
port 207 nsew power bidirectional
rlabel metal4 s 37242 496 37862 36496 6 VPWR
port 207 nsew power bidirectional
rlabel metal4 s 73242 496 73862 36496 6 VPWR
port 207 nsew power bidirectional
rlabel metal4 s 109242 496 109862 36496 6 VPWR
port 207 nsew power bidirectional
rlabel metal4 s 145242 496 145862 36496 6 VPWR
port 207 nsew power bidirectional
rlabel metal4 s 181242 496 181862 36496 6 VPWR
port 207 nsew power bidirectional
rlabel metal4 s 217242 496 217862 36496 6 VPWR
port 207 nsew power bidirectional
rlabel metal3 s 234292 4224 234692 4344 6 WE0[0]
port 208 nsew signal input
rlabel metal3 s 234292 6808 234692 6928 6 WE0[1]
port 209 nsew signal input
rlabel metal3 s 234292 9392 234692 9512 6 WE0[2]
port 210 nsew signal input
rlabel metal3 s 234292 11976 234692 12096 6 WE0[3]
port 211 nsew signal input
rlabel metal3 s 234292 14560 234692 14680 6 WE0[4]
port 212 nsew signal input
rlabel metal3 s 234292 17144 234692 17264 6 WE0[5]
port 213 nsew signal input
rlabel metal3 s 234292 19728 234692 19848 6 WE0[6]
port 214 nsew signal input
rlabel metal3 s 234292 22312 234692 22432 6 WE0[7]
port 215 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 234692 37088
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 17561940
string GDS_FILE /mnt/dffram/build/32x64_1RW1R/openlane/runs/RUN_2022.09.05_22.57.31/results/signoff/RAM32_1RW1R.magic.gds
string GDS_START 150134
<< end >>

