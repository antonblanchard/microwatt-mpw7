VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM512
  CLASS BLOCK ;
  FOREIGN RAM512 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1583.780 BY 987.360 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 520.240 1583.780 520.840 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 574.640 1583.780 575.240 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 629.040 1583.780 629.640 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 683.440 1583.780 684.040 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 737.840 1583.780 738.440 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 792.240 1583.780 792.840 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 846.640 1583.780 847.240 ;
    END
  END A0[6]
  PIN A0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 901.040 1583.780 901.640 ;
    END
  END A0[7]
  PIN A0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 955.440 1583.780 956.040 ;
    END
  END A0[8]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 2.000 493.640 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 2.000 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 2.000 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 2.000 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 2.000 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 0.000 340.770 2.000 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.870 0.000 365.150 2.000 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 0.000 389.530 2.000 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 0.000 413.910 2.000 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 2.000 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 0.000 462.670 2.000 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 0.000 487.050 2.000 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 2.000 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.150 0.000 511.430 2.000 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.530 0.000 535.810 2.000 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.910 0.000 560.190 2.000 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.290 0.000 584.570 2.000 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 0.000 608.950 2.000 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.050 0.000 633.330 2.000 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.430 0.000 657.710 2.000 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.810 0.000 682.090 2.000 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.190 0.000 706.470 2.000 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.570 0.000 730.850 2.000 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 2.000 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.950 0.000 755.230 2.000 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 0.000 779.610 2.000 ;
    END
  END Di0[31]
  PIN Di0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.710 0.000 803.990 2.000 ;
    END
  END Di0[32]
  PIN Di0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.090 0.000 828.370 2.000 ;
    END
  END Di0[33]
  PIN Di0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.470 0.000 852.750 2.000 ;
    END
  END Di0[34]
  PIN Di0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.850 0.000 877.130 2.000 ;
    END
  END Di0[35]
  PIN Di0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.230 0.000 901.510 2.000 ;
    END
  END Di0[36]
  PIN Di0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 925.610 0.000 925.890 2.000 ;
    END
  END Di0[37]
  PIN Di0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.990 0.000 950.270 2.000 ;
    END
  END Di0[38]
  PIN Di0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 974.370 0.000 974.650 2.000 ;
    END
  END Di0[39]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 2.000 ;
    END
  END Di0[3]
  PIN Di0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.750 0.000 999.030 2.000 ;
    END
  END Di0[40]
  PIN Di0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1023.130 0.000 1023.410 2.000 ;
    END
  END Di0[41]
  PIN Di0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.510 0.000 1047.790 2.000 ;
    END
  END Di0[42]
  PIN Di0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.890 0.000 1072.170 2.000 ;
    END
  END Di0[43]
  PIN Di0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1096.270 0.000 1096.550 2.000 ;
    END
  END Di0[44]
  PIN Di0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.650 0.000 1120.930 2.000 ;
    END
  END Di0[45]
  PIN Di0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.030 0.000 1145.310 2.000 ;
    END
  END Di0[46]
  PIN Di0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1169.410 0.000 1169.690 2.000 ;
    END
  END Di0[47]
  PIN Di0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1193.790 0.000 1194.070 2.000 ;
    END
  END Di0[48]
  PIN Di0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1218.170 0.000 1218.450 2.000 ;
    END
  END Di0[49]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 2.000 ;
    END
  END Di0[4]
  PIN Di0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1242.550 0.000 1242.830 2.000 ;
    END
  END Di0[50]
  PIN Di0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.930 0.000 1267.210 2.000 ;
    END
  END Di0[51]
  PIN Di0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.310 0.000 1291.590 2.000 ;
    END
  END Di0[52]
  PIN Di0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1315.690 0.000 1315.970 2.000 ;
    END
  END Di0[53]
  PIN Di0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.070 0.000 1340.350 2.000 ;
    END
  END Di0[54]
  PIN Di0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1364.450 0.000 1364.730 2.000 ;
    END
  END Di0[55]
  PIN Di0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1388.830 0.000 1389.110 2.000 ;
    END
  END Di0[56]
  PIN Di0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.210 0.000 1413.490 2.000 ;
    END
  END Di0[57]
  PIN Di0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1437.590 0.000 1437.870 2.000 ;
    END
  END Di0[58]
  PIN Di0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1461.970 0.000 1462.250 2.000 ;
    END
  END Di0[59]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 2.000 ;
    END
  END Di0[5]
  PIN Di0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1486.350 0.000 1486.630 2.000 ;
    END
  END Di0[60]
  PIN Di0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1510.730 0.000 1511.010 2.000 ;
    END
  END Di0[61]
  PIN Di0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1535.110 0.000 1535.390 2.000 ;
    END
  END Di0[62]
  PIN Di0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1559.490 0.000 1559.770 2.000 ;
    END
  END Di0[63]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 0.000 170.110 2.000 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 2.000 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 2.000 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 2.000 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 985.360 23.830 987.360 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 985.360 267.630 987.360 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 985.360 292.010 987.360 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 985.360 316.390 987.360 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 985.360 340.770 987.360 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.870 985.360 365.150 987.360 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 985.360 389.530 987.360 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 985.360 413.910 987.360 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 985.360 438.290 987.360 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 985.360 462.670 987.360 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 985.360 487.050 987.360 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 985.360 48.210 987.360 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.150 985.360 511.430 987.360 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.530 985.360 535.810 987.360 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.910 985.360 560.190 987.360 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.290 985.360 584.570 987.360 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 985.360 608.950 987.360 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.050 985.360 633.330 987.360 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.430 985.360 657.710 987.360 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.810 985.360 682.090 987.360 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.190 985.360 706.470 987.360 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.570 985.360 730.850 987.360 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 985.360 72.590 987.360 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.950 985.360 755.230 987.360 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 985.360 779.610 987.360 ;
    END
  END Do0[31]
  PIN Do0[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.710 985.360 803.990 987.360 ;
    END
  END Do0[32]
  PIN Do0[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.090 985.360 828.370 987.360 ;
    END
  END Do0[33]
  PIN Do0[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.470 985.360 852.750 987.360 ;
    END
  END Do0[34]
  PIN Do0[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.850 985.360 877.130 987.360 ;
    END
  END Do0[35]
  PIN Do0[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.230 985.360 901.510 987.360 ;
    END
  END Do0[36]
  PIN Do0[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 925.610 985.360 925.890 987.360 ;
    END
  END Do0[37]
  PIN Do0[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.990 985.360 950.270 987.360 ;
    END
  END Do0[38]
  PIN Do0[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 974.370 985.360 974.650 987.360 ;
    END
  END Do0[39]
  PIN Do0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 985.360 96.970 987.360 ;
    END
  END Do0[3]
  PIN Do0[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.750 985.360 999.030 987.360 ;
    END
  END Do0[40]
  PIN Do0[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1023.130 985.360 1023.410 987.360 ;
    END
  END Do0[41]
  PIN Do0[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.510 985.360 1047.790 987.360 ;
    END
  END Do0[42]
  PIN Do0[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.890 985.360 1072.170 987.360 ;
    END
  END Do0[43]
  PIN Do0[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1096.270 985.360 1096.550 987.360 ;
    END
  END Do0[44]
  PIN Do0[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.650 985.360 1120.930 987.360 ;
    END
  END Do0[45]
  PIN Do0[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.030 985.360 1145.310 987.360 ;
    END
  END Do0[46]
  PIN Do0[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1169.410 985.360 1169.690 987.360 ;
    END
  END Do0[47]
  PIN Do0[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1193.790 985.360 1194.070 987.360 ;
    END
  END Do0[48]
  PIN Do0[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1218.170 985.360 1218.450 987.360 ;
    END
  END Do0[49]
  PIN Do0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 985.360 121.350 987.360 ;
    END
  END Do0[4]
  PIN Do0[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1242.550 985.360 1242.830 987.360 ;
    END
  END Do0[50]
  PIN Do0[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.930 985.360 1267.210 987.360 ;
    END
  END Do0[51]
  PIN Do0[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.310 985.360 1291.590 987.360 ;
    END
  END Do0[52]
  PIN Do0[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1315.690 985.360 1315.970 987.360 ;
    END
  END Do0[53]
  PIN Do0[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.070 985.360 1340.350 987.360 ;
    END
  END Do0[54]
  PIN Do0[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1364.450 985.360 1364.730 987.360 ;
    END
  END Do0[55]
  PIN Do0[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1388.830 985.360 1389.110 987.360 ;
    END
  END Do0[56]
  PIN Do0[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.210 985.360 1413.490 987.360 ;
    END
  END Do0[57]
  PIN Do0[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1437.590 985.360 1437.870 987.360 ;
    END
  END Do0[58]
  PIN Do0[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1461.970 985.360 1462.250 987.360 ;
    END
  END Do0[59]
  PIN Do0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 985.360 145.730 987.360 ;
    END
  END Do0[5]
  PIN Do0[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1486.350 985.360 1486.630 987.360 ;
    END
  END Do0[60]
  PIN Do0[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1510.730 985.360 1511.010 987.360 ;
    END
  END Do0[61]
  PIN Do0[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1535.110 985.360 1535.390 987.360 ;
    END
  END Do0[62]
  PIN Do0[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1559.490 985.360 1559.770 987.360 ;
    END
  END Do0[63]
  PIN Do0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 985.360 170.110 987.360 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 985.360 194.490 987.360 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 985.360 218.870 987.360 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 985.360 243.250 987.360 ;
    END
  END Do0[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 30.640 1583.780 31.240 ;
    END
  END EN0
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 113.690 100.400 116.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 293.690 100.400 296.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 473.690 100.400 476.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 653.690 100.400 656.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 833.690 100.400 836.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1013.690 100.400 1016.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1193.690 100.400 1196.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1373.690 100.400 1376.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1553.690 100.400 1556.790 886.960 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 23.690 100.400 26.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 203.690 100.400 206.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 383.690 100.400 386.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.690 100.400 566.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 743.690 100.400 746.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 923.690 100.400 926.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1103.690 100.400 1106.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1283.690 100.400 1286.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1463.690 100.400 1466.790 886.960 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 85.040 1583.780 85.640 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 139.440 1583.780 140.040 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 193.840 1583.780 194.440 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 248.240 1583.780 248.840 ;
    END
  END WE0[3]
  PIN WE0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 302.640 1583.780 303.240 ;
    END
  END WE0[4]
  PIN WE0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 357.040 1583.780 357.640 ;
    END
  END WE0[5]
  PIN WE0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 411.440 1583.780 412.040 ;
    END
  END WE0[6]
  PIN WE0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 465.840 1583.780 466.440 ;
    END
  END WE0[7]
  OBS
      LAYER li1 ;
        RECT 20.240 100.555 1563.540 886.805 ;
      LAYER met1 ;
        RECT 3.290 0.380 1575.430 987.320 ;
      LAYER met2 ;
        RECT 3.320 985.080 23.270 987.350 ;
        RECT 24.110 985.080 47.650 987.350 ;
        RECT 48.490 985.080 72.030 987.350 ;
        RECT 72.870 985.080 96.410 987.350 ;
        RECT 97.250 985.080 120.790 987.350 ;
        RECT 121.630 985.080 145.170 987.350 ;
        RECT 146.010 985.080 169.550 987.350 ;
        RECT 170.390 985.080 193.930 987.350 ;
        RECT 194.770 985.080 218.310 987.350 ;
        RECT 219.150 985.080 242.690 987.350 ;
        RECT 243.530 985.080 267.070 987.350 ;
        RECT 267.910 985.080 291.450 987.350 ;
        RECT 292.290 985.080 315.830 987.350 ;
        RECT 316.670 985.080 340.210 987.350 ;
        RECT 341.050 985.080 364.590 987.350 ;
        RECT 365.430 985.080 388.970 987.350 ;
        RECT 389.810 985.080 413.350 987.350 ;
        RECT 414.190 985.080 437.730 987.350 ;
        RECT 438.570 985.080 462.110 987.350 ;
        RECT 462.950 985.080 486.490 987.350 ;
        RECT 487.330 985.080 510.870 987.350 ;
        RECT 511.710 985.080 535.250 987.350 ;
        RECT 536.090 985.080 559.630 987.350 ;
        RECT 560.470 985.080 584.010 987.350 ;
        RECT 584.850 985.080 608.390 987.350 ;
        RECT 609.230 985.080 632.770 987.350 ;
        RECT 633.610 985.080 657.150 987.350 ;
        RECT 657.990 985.080 681.530 987.350 ;
        RECT 682.370 985.080 705.910 987.350 ;
        RECT 706.750 985.080 730.290 987.350 ;
        RECT 731.130 985.080 754.670 987.350 ;
        RECT 755.510 985.080 779.050 987.350 ;
        RECT 779.890 985.080 803.430 987.350 ;
        RECT 804.270 985.080 827.810 987.350 ;
        RECT 828.650 985.080 852.190 987.350 ;
        RECT 853.030 985.080 876.570 987.350 ;
        RECT 877.410 985.080 900.950 987.350 ;
        RECT 901.790 985.080 925.330 987.350 ;
        RECT 926.170 985.080 949.710 987.350 ;
        RECT 950.550 985.080 974.090 987.350 ;
        RECT 974.930 985.080 998.470 987.350 ;
        RECT 999.310 985.080 1022.850 987.350 ;
        RECT 1023.690 985.080 1047.230 987.350 ;
        RECT 1048.070 985.080 1071.610 987.350 ;
        RECT 1072.450 985.080 1095.990 987.350 ;
        RECT 1096.830 985.080 1120.370 987.350 ;
        RECT 1121.210 985.080 1144.750 987.350 ;
        RECT 1145.590 985.080 1169.130 987.350 ;
        RECT 1169.970 985.080 1193.510 987.350 ;
        RECT 1194.350 985.080 1217.890 987.350 ;
        RECT 1218.730 985.080 1242.270 987.350 ;
        RECT 1243.110 985.080 1266.650 987.350 ;
        RECT 1267.490 985.080 1291.030 987.350 ;
        RECT 1291.870 985.080 1315.410 987.350 ;
        RECT 1316.250 985.080 1339.790 987.350 ;
        RECT 1340.630 985.080 1364.170 987.350 ;
        RECT 1365.010 985.080 1388.550 987.350 ;
        RECT 1389.390 985.080 1412.930 987.350 ;
        RECT 1413.770 985.080 1437.310 987.350 ;
        RECT 1438.150 985.080 1461.690 987.350 ;
        RECT 1462.530 985.080 1486.070 987.350 ;
        RECT 1486.910 985.080 1510.450 987.350 ;
        RECT 1511.290 985.080 1534.830 987.350 ;
        RECT 1535.670 985.080 1559.210 987.350 ;
        RECT 1560.050 985.080 1575.410 987.350 ;
        RECT 3.320 2.280 1575.410 985.080 ;
        RECT 3.320 0.350 23.270 2.280 ;
        RECT 24.110 0.350 47.650 2.280 ;
        RECT 48.490 0.350 72.030 2.280 ;
        RECT 72.870 0.350 96.410 2.280 ;
        RECT 97.250 0.350 120.790 2.280 ;
        RECT 121.630 0.350 145.170 2.280 ;
        RECT 146.010 0.350 169.550 2.280 ;
        RECT 170.390 0.350 193.930 2.280 ;
        RECT 194.770 0.350 218.310 2.280 ;
        RECT 219.150 0.350 242.690 2.280 ;
        RECT 243.530 0.350 267.070 2.280 ;
        RECT 267.910 0.350 291.450 2.280 ;
        RECT 292.290 0.350 315.830 2.280 ;
        RECT 316.670 0.350 340.210 2.280 ;
        RECT 341.050 0.350 364.590 2.280 ;
        RECT 365.430 0.350 388.970 2.280 ;
        RECT 389.810 0.350 413.350 2.280 ;
        RECT 414.190 0.350 437.730 2.280 ;
        RECT 438.570 0.350 462.110 2.280 ;
        RECT 462.950 0.350 486.490 2.280 ;
        RECT 487.330 0.350 510.870 2.280 ;
        RECT 511.710 0.350 535.250 2.280 ;
        RECT 536.090 0.350 559.630 2.280 ;
        RECT 560.470 0.350 584.010 2.280 ;
        RECT 584.850 0.350 608.390 2.280 ;
        RECT 609.230 0.350 632.770 2.280 ;
        RECT 633.610 0.350 657.150 2.280 ;
        RECT 657.990 0.350 681.530 2.280 ;
        RECT 682.370 0.350 705.910 2.280 ;
        RECT 706.750 0.350 730.290 2.280 ;
        RECT 731.130 0.350 754.670 2.280 ;
        RECT 755.510 0.350 779.050 2.280 ;
        RECT 779.890 0.350 803.430 2.280 ;
        RECT 804.270 0.350 827.810 2.280 ;
        RECT 828.650 0.350 852.190 2.280 ;
        RECT 853.030 0.350 876.570 2.280 ;
        RECT 877.410 0.350 900.950 2.280 ;
        RECT 901.790 0.350 925.330 2.280 ;
        RECT 926.170 0.350 949.710 2.280 ;
        RECT 950.550 0.350 974.090 2.280 ;
        RECT 974.930 0.350 998.470 2.280 ;
        RECT 999.310 0.350 1022.850 2.280 ;
        RECT 1023.690 0.350 1047.230 2.280 ;
        RECT 1048.070 0.350 1071.610 2.280 ;
        RECT 1072.450 0.350 1095.990 2.280 ;
        RECT 1096.830 0.350 1120.370 2.280 ;
        RECT 1121.210 0.350 1144.750 2.280 ;
        RECT 1145.590 0.350 1169.130 2.280 ;
        RECT 1169.970 0.350 1193.510 2.280 ;
        RECT 1194.350 0.350 1217.890 2.280 ;
        RECT 1218.730 0.350 1242.270 2.280 ;
        RECT 1243.110 0.350 1266.650 2.280 ;
        RECT 1267.490 0.350 1291.030 2.280 ;
        RECT 1291.870 0.350 1315.410 2.280 ;
        RECT 1316.250 0.350 1339.790 2.280 ;
        RECT 1340.630 0.350 1364.170 2.280 ;
        RECT 1365.010 0.350 1388.550 2.280 ;
        RECT 1389.390 0.350 1412.930 2.280 ;
        RECT 1413.770 0.350 1437.310 2.280 ;
        RECT 1438.150 0.350 1461.690 2.280 ;
        RECT 1462.530 0.350 1486.070 2.280 ;
        RECT 1486.910 0.350 1510.450 2.280 ;
        RECT 1511.290 0.350 1534.830 2.280 ;
        RECT 1535.670 0.350 1559.210 2.280 ;
        RECT 1560.050 0.350 1575.410 2.280 ;
      LAYER met3 ;
        RECT 2.000 956.440 1581.780 987.185 ;
        RECT 2.000 955.040 1581.380 956.440 ;
        RECT 2.000 902.040 1581.780 955.040 ;
        RECT 2.000 900.640 1581.380 902.040 ;
        RECT 2.000 847.640 1581.780 900.640 ;
        RECT 2.000 846.240 1581.380 847.640 ;
        RECT 2.000 793.240 1581.780 846.240 ;
        RECT 2.000 791.840 1581.380 793.240 ;
        RECT 2.000 738.840 1581.780 791.840 ;
        RECT 2.000 737.440 1581.380 738.840 ;
        RECT 2.000 684.440 1581.780 737.440 ;
        RECT 2.000 683.040 1581.380 684.440 ;
        RECT 2.000 630.040 1581.780 683.040 ;
        RECT 2.000 628.640 1581.380 630.040 ;
        RECT 2.000 575.640 1581.780 628.640 ;
        RECT 2.000 574.240 1581.380 575.640 ;
        RECT 2.000 521.240 1581.780 574.240 ;
        RECT 2.000 519.840 1581.380 521.240 ;
        RECT 2.000 494.040 1581.780 519.840 ;
        RECT 2.400 492.640 1581.780 494.040 ;
        RECT 2.000 466.840 1581.780 492.640 ;
        RECT 2.000 465.440 1581.380 466.840 ;
        RECT 2.000 412.440 1581.780 465.440 ;
        RECT 2.000 411.040 1581.380 412.440 ;
        RECT 2.000 358.040 1581.780 411.040 ;
        RECT 2.000 356.640 1581.380 358.040 ;
        RECT 2.000 303.640 1581.780 356.640 ;
        RECT 2.000 302.240 1581.380 303.640 ;
        RECT 2.000 249.240 1581.780 302.240 ;
        RECT 2.000 247.840 1581.380 249.240 ;
        RECT 2.000 194.840 1581.780 247.840 ;
        RECT 2.000 193.440 1581.380 194.840 ;
        RECT 2.000 140.440 1581.780 193.440 ;
        RECT 2.000 139.040 1581.380 140.440 ;
        RECT 2.000 86.040 1581.780 139.040 ;
        RECT 2.000 84.640 1581.380 86.040 ;
        RECT 2.000 31.640 1581.780 84.640 ;
        RECT 2.000 30.240 1581.380 31.640 ;
        RECT 2.000 0.855 1581.780 30.240 ;
      LAYER met4 ;
        RECT 41.695 887.360 1566.465 987.185 ;
        RECT 41.695 100.000 113.290 887.360 ;
        RECT 117.190 100.000 203.290 887.360 ;
        RECT 207.190 100.000 293.290 887.360 ;
        RECT 297.190 100.000 383.290 887.360 ;
        RECT 387.190 100.000 473.290 887.360 ;
        RECT 477.190 100.000 563.290 887.360 ;
        RECT 567.190 100.000 653.290 887.360 ;
        RECT 657.190 100.000 743.290 887.360 ;
        RECT 747.190 100.000 833.290 887.360 ;
        RECT 837.190 100.000 923.290 887.360 ;
        RECT 927.190 100.000 1013.290 887.360 ;
        RECT 1017.190 100.000 1103.290 887.360 ;
        RECT 1107.190 100.000 1193.290 887.360 ;
        RECT 1197.190 100.000 1283.290 887.360 ;
        RECT 1287.190 100.000 1373.290 887.360 ;
        RECT 1377.190 100.000 1463.290 887.360 ;
        RECT 1467.190 100.000 1553.290 887.360 ;
        RECT 1557.190 100.000 1566.465 887.360 ;
        RECT 41.695 4.255 1566.465 100.000 ;
  END
END RAM512
END LIBRARY

